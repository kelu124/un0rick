// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Oct 7 2018 03:23:06

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MATTY_MAIN_VHDL" view "INTERFACE"

module MATTY_MAIN_VHDL (
    RAM_DATA,
    RAM_ADD,
    spi_sclk_ft,
    button_trig,
    ADC9,
    spi_cs_ft,
    poff,
    RAM_nOE,
    ADC0,
    spi_mosi_flash,
    spi_miso_flash,
    trig_ft,
    spi_miso_rpi,
    RAM_nWE,
    DAC_cs,
    ADC6,
    spi_select,
    clk,
    ADC4,
    trig_rpi,
    top_tour2,
    spi_cs_rpi,
    DAC_sclk,
    ADC_clk,
    ADC3,
    trig_ext,
    spi_mosi_rpi,
    spi_mosi_ft,
    cs_rpi2flash,
    spi_cs_flash,
    pon,
    RAM_nCE,
    LED3,
    ADC1,
    reset_rpi,
    RAM_nLB,
    LED_MODE,
    ADC8,
    spi_sclk_rpi,
    ADC7,
    top_tour1,
    spi_miso_ft,
    button_mode,
    DAC_mosi,
    ADC5,
    reset_ft,
    LED_ACQ,
    spi_sclk_flash,
    reset_alim,
    RAM_nUB,
    ADC2);

    inout [15:0] RAM_DATA;
    output [18:0] RAM_ADD;
    input spi_sclk_ft;
    input button_trig;
    input ADC9;
    input spi_cs_ft;
    output poff;
    output RAM_nOE;
    input ADC0;
    output spi_mosi_flash;
    input spi_miso_flash;
    input trig_ft;
    output spi_miso_rpi;
    output RAM_nWE;
    output DAC_cs;
    input ADC6;
    input spi_select;
    input clk;
    input ADC4;
    input trig_rpi;
    input top_tour2;
    input spi_cs_rpi;
    output DAC_sclk;
    output ADC_clk;
    input ADC3;
    input trig_ext;
    input spi_mosi_rpi;
    input spi_mosi_ft;
    input cs_rpi2flash;
    output spi_cs_flash;
    output pon;
    output RAM_nCE;
    output LED3;
    input ADC1;
    input reset_rpi;
    output RAM_nLB;
    output LED_MODE;
    input ADC8;
    input spi_sclk_rpi;
    input ADC7;
    input top_tour1;
    output spi_miso_ft;
    input button_mode;
    output DAC_mosi;
    input ADC5;
    input reset_ft;
    output LED_ACQ;
    output spi_sclk_flash;
    input reset_alim;
    output RAM_nUB;
    input ADC2;

    wire N__53520;
    wire N__53519;
    wire N__53518;
    wire N__53511;
    wire N__53510;
    wire N__53509;
    wire N__53502;
    wire N__53501;
    wire N__53500;
    wire N__53493;
    wire N__53492;
    wire N__53491;
    wire N__53484;
    wire N__53483;
    wire N__53482;
    wire N__53475;
    wire N__53474;
    wire N__53473;
    wire N__53466;
    wire N__53465;
    wire N__53464;
    wire N__53457;
    wire N__53456;
    wire N__53455;
    wire N__53448;
    wire N__53447;
    wire N__53446;
    wire N__53439;
    wire N__53438;
    wire N__53437;
    wire N__53430;
    wire N__53429;
    wire N__53428;
    wire N__53421;
    wire N__53420;
    wire N__53419;
    wire N__53412;
    wire N__53411;
    wire N__53410;
    wire N__53403;
    wire N__53402;
    wire N__53401;
    wire N__53394;
    wire N__53393;
    wire N__53392;
    wire N__53385;
    wire N__53384;
    wire N__53383;
    wire N__53376;
    wire N__53375;
    wire N__53374;
    wire N__53367;
    wire N__53366;
    wire N__53365;
    wire N__53358;
    wire N__53357;
    wire N__53356;
    wire N__53349;
    wire N__53348;
    wire N__53347;
    wire N__53340;
    wire N__53339;
    wire N__53338;
    wire N__53331;
    wire N__53330;
    wire N__53329;
    wire N__53322;
    wire N__53321;
    wire N__53320;
    wire N__53313;
    wire N__53312;
    wire N__53311;
    wire N__53304;
    wire N__53303;
    wire N__53302;
    wire N__53295;
    wire N__53294;
    wire N__53293;
    wire N__53286;
    wire N__53285;
    wire N__53284;
    wire N__53277;
    wire N__53276;
    wire N__53275;
    wire N__53268;
    wire N__53267;
    wire N__53266;
    wire N__53259;
    wire N__53258;
    wire N__53257;
    wire N__53250;
    wire N__53249;
    wire N__53248;
    wire N__53241;
    wire N__53240;
    wire N__53239;
    wire N__53232;
    wire N__53231;
    wire N__53230;
    wire N__53223;
    wire N__53222;
    wire N__53221;
    wire N__53214;
    wire N__53213;
    wire N__53212;
    wire N__53205;
    wire N__53204;
    wire N__53203;
    wire N__53196;
    wire N__53195;
    wire N__53194;
    wire N__53187;
    wire N__53186;
    wire N__53185;
    wire N__53178;
    wire N__53177;
    wire N__53176;
    wire N__53169;
    wire N__53168;
    wire N__53167;
    wire N__53160;
    wire N__53159;
    wire N__53158;
    wire N__53151;
    wire N__53150;
    wire N__53149;
    wire N__53142;
    wire N__53141;
    wire N__53140;
    wire N__53133;
    wire N__53132;
    wire N__53131;
    wire N__53124;
    wire N__53123;
    wire N__53122;
    wire N__53115;
    wire N__53114;
    wire N__53113;
    wire N__53106;
    wire N__53105;
    wire N__53104;
    wire N__53097;
    wire N__53096;
    wire N__53095;
    wire N__53088;
    wire N__53087;
    wire N__53086;
    wire N__53079;
    wire N__53078;
    wire N__53077;
    wire N__53070;
    wire N__53069;
    wire N__53068;
    wire N__53061;
    wire N__53060;
    wire N__53059;
    wire N__53052;
    wire N__53051;
    wire N__53050;
    wire N__53043;
    wire N__53042;
    wire N__53041;
    wire N__53034;
    wire N__53033;
    wire N__53032;
    wire N__53025;
    wire N__53024;
    wire N__53023;
    wire N__53016;
    wire N__53015;
    wire N__53014;
    wire N__53007;
    wire N__53006;
    wire N__53005;
    wire N__52998;
    wire N__52997;
    wire N__52996;
    wire N__52989;
    wire N__52988;
    wire N__52987;
    wire N__52980;
    wire N__52979;
    wire N__52978;
    wire N__52971;
    wire N__52970;
    wire N__52969;
    wire N__52962;
    wire N__52961;
    wire N__52960;
    wire N__52953;
    wire N__52952;
    wire N__52951;
    wire N__52944;
    wire N__52943;
    wire N__52942;
    wire N__52935;
    wire N__52934;
    wire N__52933;
    wire N__52926;
    wire N__52925;
    wire N__52924;
    wire N__52917;
    wire N__52916;
    wire N__52915;
    wire N__52908;
    wire N__52907;
    wire N__52906;
    wire N__52899;
    wire N__52898;
    wire N__52897;
    wire N__52890;
    wire N__52889;
    wire N__52888;
    wire N__52881;
    wire N__52880;
    wire N__52879;
    wire N__52872;
    wire N__52871;
    wire N__52870;
    wire N__52863;
    wire N__52862;
    wire N__52861;
    wire N__52854;
    wire N__52853;
    wire N__52852;
    wire N__52845;
    wire N__52844;
    wire N__52843;
    wire N__52836;
    wire N__52835;
    wire N__52834;
    wire N__52827;
    wire N__52826;
    wire N__52825;
    wire N__52818;
    wire N__52817;
    wire N__52816;
    wire N__52809;
    wire N__52808;
    wire N__52807;
    wire N__52790;
    wire N__52789;
    wire N__52788;
    wire N__52787;
    wire N__52786;
    wire N__52785;
    wire N__52784;
    wire N__52783;
    wire N__52782;
    wire N__52781;
    wire N__52780;
    wire N__52779;
    wire N__52770;
    wire N__52769;
    wire N__52768;
    wire N__52767;
    wire N__52766;
    wire N__52765;
    wire N__52764;
    wire N__52763;
    wire N__52760;
    wire N__52759;
    wire N__52756;
    wire N__52755;
    wire N__52752;
    wire N__52751;
    wire N__52748;
    wire N__52747;
    wire N__52746;
    wire N__52745;
    wire N__52744;
    wire N__52743;
    wire N__52742;
    wire N__52739;
    wire N__52738;
    wire N__52731;
    wire N__52728;
    wire N__52721;
    wire N__52712;
    wire N__52711;
    wire N__52710;
    wire N__52709;
    wire N__52708;
    wire N__52707;
    wire N__52706;
    wire N__52705;
    wire N__52688;
    wire N__52685;
    wire N__52684;
    wire N__52681;
    wire N__52680;
    wire N__52677;
    wire N__52676;
    wire N__52673;
    wire N__52672;
    wire N__52671;
    wire N__52670;
    wire N__52669;
    wire N__52668;
    wire N__52661;
    wire N__52658;
    wire N__52651;
    wire N__52650;
    wire N__52649;
    wire N__52646;
    wire N__52643;
    wire N__52640;
    wire N__52639;
    wire N__52636;
    wire N__52633;
    wire N__52630;
    wire N__52627;
    wire N__52626;
    wire N__52625;
    wire N__52624;
    wire N__52623;
    wire N__52620;
    wire N__52603;
    wire N__52602;
    wire N__52599;
    wire N__52598;
    wire N__52595;
    wire N__52594;
    wire N__52591;
    wire N__52590;
    wire N__52587;
    wire N__52586;
    wire N__52579;
    wire N__52574;
    wire N__52573;
    wire N__52572;
    wire N__52571;
    wire N__52570;
    wire N__52563;
    wire N__52552;
    wire N__52549;
    wire N__52548;
    wire N__52545;
    wire N__52544;
    wire N__52541;
    wire N__52540;
    wire N__52537;
    wire N__52536;
    wire N__52531;
    wire N__52514;
    wire N__52511;
    wire N__52510;
    wire N__52507;
    wire N__52504;
    wire N__52503;
    wire N__52500;
    wire N__52499;
    wire N__52496;
    wire N__52495;
    wire N__52492;
    wire N__52491;
    wire N__52488;
    wire N__52485;
    wire N__52482;
    wire N__52465;
    wire N__52460;
    wire N__52455;
    wire N__52450;
    wire N__52433;
    wire N__52428;
    wire N__52425;
    wire N__52420;
    wire N__52417;
    wire N__52414;
    wire N__52409;
    wire N__52408;
    wire N__52405;
    wire N__52402;
    wire N__52399;
    wire N__52396;
    wire N__52393;
    wire N__52390;
    wire N__52385;
    wire N__52380;
    wire N__52377;
    wire N__52372;
    wire N__52367;
    wire N__52364;
    wire N__52361;
    wire N__52358;
    wire N__52355;
    wire N__52352;
    wire N__52349;
    wire N__52348;
    wire N__52347;
    wire N__52346;
    wire N__52345;
    wire N__52344;
    wire N__52343;
    wire N__52342;
    wire N__52341;
    wire N__52340;
    wire N__52339;
    wire N__52338;
    wire N__52337;
    wire N__52336;
    wire N__52335;
    wire N__52334;
    wire N__52333;
    wire N__52332;
    wire N__52331;
    wire N__52330;
    wire N__52329;
    wire N__52328;
    wire N__52327;
    wire N__52326;
    wire N__52325;
    wire N__52324;
    wire N__52323;
    wire N__52322;
    wire N__52321;
    wire N__52320;
    wire N__52319;
    wire N__52318;
    wire N__52317;
    wire N__52316;
    wire N__52315;
    wire N__52314;
    wire N__52313;
    wire N__52312;
    wire N__52311;
    wire N__52310;
    wire N__52309;
    wire N__52308;
    wire N__52307;
    wire N__52306;
    wire N__52305;
    wire N__52304;
    wire N__52303;
    wire N__52302;
    wire N__52301;
    wire N__52300;
    wire N__52299;
    wire N__52298;
    wire N__52297;
    wire N__52296;
    wire N__52295;
    wire N__52294;
    wire N__52293;
    wire N__52292;
    wire N__52291;
    wire N__52290;
    wire N__52289;
    wire N__52288;
    wire N__52287;
    wire N__52286;
    wire N__52285;
    wire N__52284;
    wire N__52283;
    wire N__52282;
    wire N__52281;
    wire N__52280;
    wire N__52279;
    wire N__52278;
    wire N__52277;
    wire N__52276;
    wire N__52275;
    wire N__52274;
    wire N__52273;
    wire N__52272;
    wire N__52271;
    wire N__52270;
    wire N__52269;
    wire N__52268;
    wire N__52267;
    wire N__52266;
    wire N__52265;
    wire N__52264;
    wire N__52263;
    wire N__52262;
    wire N__52261;
    wire N__52260;
    wire N__52259;
    wire N__52258;
    wire N__52257;
    wire N__52256;
    wire N__52255;
    wire N__52254;
    wire N__52253;
    wire N__52252;
    wire N__52251;
    wire N__52250;
    wire N__52249;
    wire N__52248;
    wire N__52247;
    wire N__52246;
    wire N__52245;
    wire N__52244;
    wire N__52243;
    wire N__52242;
    wire N__52241;
    wire N__52240;
    wire N__52239;
    wire N__52238;
    wire N__52237;
    wire N__52236;
    wire N__52235;
    wire N__52234;
    wire N__52233;
    wire N__52232;
    wire N__52231;
    wire N__52230;
    wire N__52229;
    wire N__52228;
    wire N__52227;
    wire N__52226;
    wire N__52225;
    wire N__52224;
    wire N__52223;
    wire N__52222;
    wire N__52221;
    wire N__52220;
    wire N__52219;
    wire N__52218;
    wire N__52217;
    wire N__52216;
    wire N__52215;
    wire N__52214;
    wire N__52213;
    wire N__52212;
    wire N__52211;
    wire N__52210;
    wire N__52209;
    wire N__52208;
    wire N__52207;
    wire N__52206;
    wire N__52205;
    wire N__52204;
    wire N__52203;
    wire N__52202;
    wire N__52201;
    wire N__51902;
    wire N__51899;
    wire N__51896;
    wire N__51895;
    wire N__51894;
    wire N__51891;
    wire N__51890;
    wire N__51889;
    wire N__51886;
    wire N__51883;
    wire N__51882;
    wire N__51879;
    wire N__51876;
    wire N__51873;
    wire N__51872;
    wire N__51869;
    wire N__51866;
    wire N__51863;
    wire N__51858;
    wire N__51855;
    wire N__51852;
    wire N__51849;
    wire N__51844;
    wire N__51841;
    wire N__51836;
    wire N__51827;
    wire N__51826;
    wire N__51825;
    wire N__51824;
    wire N__51823;
    wire N__51822;
    wire N__51821;
    wire N__51820;
    wire N__51819;
    wire N__51818;
    wire N__51817;
    wire N__51816;
    wire N__51815;
    wire N__51814;
    wire N__51813;
    wire N__51812;
    wire N__51811;
    wire N__51810;
    wire N__51809;
    wire N__51808;
    wire N__51807;
    wire N__51806;
    wire N__51805;
    wire N__51804;
    wire N__51803;
    wire N__51802;
    wire N__51801;
    wire N__51800;
    wire N__51799;
    wire N__51798;
    wire N__51797;
    wire N__51796;
    wire N__51795;
    wire N__51794;
    wire N__51793;
    wire N__51792;
    wire N__51791;
    wire N__51790;
    wire N__51789;
    wire N__51788;
    wire N__51787;
    wire N__51786;
    wire N__51785;
    wire N__51784;
    wire N__51783;
    wire N__51782;
    wire N__51781;
    wire N__51780;
    wire N__51779;
    wire N__51778;
    wire N__51777;
    wire N__51776;
    wire N__51775;
    wire N__51774;
    wire N__51773;
    wire N__51772;
    wire N__51771;
    wire N__51770;
    wire N__51769;
    wire N__51768;
    wire N__51767;
    wire N__51766;
    wire N__51765;
    wire N__51764;
    wire N__51763;
    wire N__51762;
    wire N__51761;
    wire N__51760;
    wire N__51759;
    wire N__51758;
    wire N__51757;
    wire N__51756;
    wire N__51755;
    wire N__51754;
    wire N__51753;
    wire N__51752;
    wire N__51751;
    wire N__51750;
    wire N__51749;
    wire N__51748;
    wire N__51747;
    wire N__51746;
    wire N__51745;
    wire N__51744;
    wire N__51743;
    wire N__51742;
    wire N__51741;
    wire N__51740;
    wire N__51739;
    wire N__51738;
    wire N__51737;
    wire N__51736;
    wire N__51735;
    wire N__51734;
    wire N__51733;
    wire N__51732;
    wire N__51731;
    wire N__51730;
    wire N__51729;
    wire N__51728;
    wire N__51727;
    wire N__51726;
    wire N__51725;
    wire N__51724;
    wire N__51723;
    wire N__51722;
    wire N__51721;
    wire N__51720;
    wire N__51719;
    wire N__51718;
    wire N__51717;
    wire N__51716;
    wire N__51715;
    wire N__51714;
    wire N__51713;
    wire N__51712;
    wire N__51711;
    wire N__51710;
    wire N__51709;
    wire N__51708;
    wire N__51707;
    wire N__51706;
    wire N__51705;
    wire N__51704;
    wire N__51703;
    wire N__51702;
    wire N__51701;
    wire N__51700;
    wire N__51699;
    wire N__51698;
    wire N__51697;
    wire N__51696;
    wire N__51695;
    wire N__51694;
    wire N__51693;
    wire N__51692;
    wire N__51691;
    wire N__51690;
    wire N__51689;
    wire N__51688;
    wire N__51687;
    wire N__51686;
    wire N__51685;
    wire N__51684;
    wire N__51683;
    wire N__51682;
    wire N__51681;
    wire N__51680;
    wire N__51679;
    wire N__51678;
    wire N__51677;
    wire N__51676;
    wire N__51675;
    wire N__51674;
    wire N__51673;
    wire N__51672;
    wire N__51671;
    wire N__51670;
    wire N__51669;
    wire N__51668;
    wire N__51667;
    wire N__51666;
    wire N__51665;
    wire N__51664;
    wire N__51663;
    wire N__51662;
    wire N__51661;
    wire N__51660;
    wire N__51659;
    wire N__51658;
    wire N__51657;
    wire N__51656;
    wire N__51655;
    wire N__51654;
    wire N__51653;
    wire N__51652;
    wire N__51651;
    wire N__51650;
    wire N__51649;
    wire N__51648;
    wire N__51647;
    wire N__51646;
    wire N__51645;
    wire N__51644;
    wire N__51643;
    wire N__51642;
    wire N__51269;
    wire N__51266;
    wire N__51263;
    wire N__51262;
    wire N__51259;
    wire N__51256;
    wire N__51253;
    wire N__51248;
    wire N__51245;
    wire N__51242;
    wire N__51241;
    wire N__51238;
    wire N__51235;
    wire N__51232;
    wire N__51227;
    wire N__51224;
    wire N__51223;
    wire N__51220;
    wire N__51217;
    wire N__51216;
    wire N__51215;
    wire N__51214;
    wire N__51213;
    wire N__51208;
    wire N__51205;
    wire N__51198;
    wire N__51197;
    wire N__51192;
    wire N__51191;
    wire N__51188;
    wire N__51185;
    wire N__51182;
    wire N__51179;
    wire N__51178;
    wire N__51175;
    wire N__51172;
    wire N__51169;
    wire N__51166;
    wire N__51163;
    wire N__51158;
    wire N__51151;
    wire N__51146;
    wire N__51145;
    wire N__51144;
    wire N__51143;
    wire N__51138;
    wire N__51133;
    wire N__51128;
    wire N__51125;
    wire N__51124;
    wire N__51121;
    wire N__51118;
    wire N__51113;
    wire N__51110;
    wire N__51107;
    wire N__51104;
    wire N__51101;
    wire N__51100;
    wire N__51097;
    wire N__51094;
    wire N__51089;
    wire N__51086;
    wire N__51083;
    wire N__51080;
    wire N__51077;
    wire N__51076;
    wire N__51075;
    wire N__51074;
    wire N__51071;
    wire N__51070;
    wire N__51069;
    wire N__51068;
    wire N__51065;
    wire N__51064;
    wire N__51063;
    wire N__51062;
    wire N__51059;
    wire N__51056;
    wire N__51055;
    wire N__51054;
    wire N__51053;
    wire N__51052;
    wire N__51051;
    wire N__51050;
    wire N__51047;
    wire N__51044;
    wire N__51043;
    wire N__51042;
    wire N__51041;
    wire N__51040;
    wire N__51039;
    wire N__51038;
    wire N__51037;
    wire N__51034;
    wire N__51031;
    wire N__51030;
    wire N__51029;
    wire N__51026;
    wire N__51023;
    wire N__51020;
    wire N__51019;
    wire N__51018;
    wire N__51017;
    wire N__51014;
    wire N__51009;
    wire N__51006;
    wire N__51003;
    wire N__51000;
    wire N__50997;
    wire N__50994;
    wire N__50991;
    wire N__50986;
    wire N__50985;
    wire N__50984;
    wire N__50983;
    wire N__50982;
    wire N__50979;
    wire N__50976;
    wire N__50973;
    wire N__50970;
    wire N__50967;
    wire N__50964;
    wire N__50961;
    wire N__50956;
    wire N__50953;
    wire N__50950;
    wire N__50943;
    wire N__50940;
    wire N__50939;
    wire N__50938;
    wire N__50935;
    wire N__50932;
    wire N__50931;
    wire N__50930;
    wire N__50929;
    wire N__50928;
    wire N__50925;
    wire N__50914;
    wire N__50907;
    wire N__50904;
    wire N__50903;
    wire N__50900;
    wire N__50899;
    wire N__50898;
    wire N__50897;
    wire N__50896;
    wire N__50893;
    wire N__50892;
    wire N__50889;
    wire N__50884;
    wire N__50883;
    wire N__50882;
    wire N__50881;
    wire N__50880;
    wire N__50879;
    wire N__50878;
    wire N__50877;
    wire N__50872;
    wire N__50861;
    wire N__50858;
    wire N__50855;
    wire N__50852;
    wire N__50851;
    wire N__50848;
    wire N__50845;
    wire N__50840;
    wire N__50837;
    wire N__50834;
    wire N__50831;
    wire N__50828;
    wire N__50825;
    wire N__50820;
    wire N__50817;
    wire N__50816;
    wire N__50815;
    wire N__50814;
    wire N__50811;
    wire N__50808;
    wire N__50805;
    wire N__50802;
    wire N__50799;
    wire N__50796;
    wire N__50793;
    wire N__50790;
    wire N__50787;
    wire N__50784;
    wire N__50781;
    wire N__50778;
    wire N__50775;
    wire N__50772;
    wire N__50769;
    wire N__50766;
    wire N__50763;
    wire N__50758;
    wire N__50755;
    wire N__50750;
    wire N__50747;
    wire N__50742;
    wire N__50739;
    wire N__50724;
    wire N__50719;
    wire N__50718;
    wire N__50717;
    wire N__50716;
    wire N__50715;
    wire N__50712;
    wire N__50707;
    wire N__50696;
    wire N__50689;
    wire N__50682;
    wire N__50667;
    wire N__50664;
    wire N__50655;
    wire N__50652;
    wire N__50649;
    wire N__50646;
    wire N__50643;
    wire N__50634;
    wire N__50629;
    wire N__50624;
    wire N__50609;
    wire N__50606;
    wire N__50603;
    wire N__50600;
    wire N__50597;
    wire N__50594;
    wire N__50593;
    wire N__50590;
    wire N__50587;
    wire N__50584;
    wire N__50581;
    wire N__50578;
    wire N__50575;
    wire N__50570;
    wire N__50567;
    wire N__50564;
    wire N__50561;
    wire N__50558;
    wire N__50555;
    wire N__50552;
    wire N__50549;
    wire N__50546;
    wire N__50545;
    wire N__50544;
    wire N__50543;
    wire N__50542;
    wire N__50541;
    wire N__50538;
    wire N__50535;
    wire N__50532;
    wire N__50531;
    wire N__50530;
    wire N__50529;
    wire N__50528;
    wire N__50527;
    wire N__50526;
    wire N__50523;
    wire N__50520;
    wire N__50517;
    wire N__50516;
    wire N__50513;
    wire N__50508;
    wire N__50505;
    wire N__50502;
    wire N__50499;
    wire N__50496;
    wire N__50495;
    wire N__50492;
    wire N__50489;
    wire N__50488;
    wire N__50487;
    wire N__50486;
    wire N__50485;
    wire N__50484;
    wire N__50483;
    wire N__50482;
    wire N__50481;
    wire N__50480;
    wire N__50473;
    wire N__50470;
    wire N__50469;
    wire N__50468;
    wire N__50467;
    wire N__50466;
    wire N__50465;
    wire N__50464;
    wire N__50463;
    wire N__50452;
    wire N__50449;
    wire N__50446;
    wire N__50443;
    wire N__50440;
    wire N__50437;
    wire N__50434;
    wire N__50431;
    wire N__50430;
    wire N__50427;
    wire N__50424;
    wire N__50421;
    wire N__50420;
    wire N__50417;
    wire N__50414;
    wire N__50413;
    wire N__50410;
    wire N__50409;
    wire N__50408;
    wire N__50407;
    wire N__50402;
    wire N__50399;
    wire N__50396;
    wire N__50393;
    wire N__50392;
    wire N__50391;
    wire N__50388;
    wire N__50385;
    wire N__50382;
    wire N__50381;
    wire N__50380;
    wire N__50379;
    wire N__50378;
    wire N__50375;
    wire N__50374;
    wire N__50367;
    wire N__50356;
    wire N__50353;
    wire N__50346;
    wire N__50343;
    wire N__50338;
    wire N__50335;
    wire N__50334;
    wire N__50331;
    wire N__50330;
    wire N__50329;
    wire N__50328;
    wire N__50327;
    wire N__50324;
    wire N__50321;
    wire N__50318;
    wire N__50317;
    wire N__50310;
    wire N__50309;
    wire N__50308;
    wire N__50307;
    wire N__50306;
    wire N__50305;
    wire N__50302;
    wire N__50299;
    wire N__50296;
    wire N__50289;
    wire N__50286;
    wire N__50283;
    wire N__50280;
    wire N__50277;
    wire N__50274;
    wire N__50271;
    wire N__50268;
    wire N__50261;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50242;
    wire N__50239;
    wire N__50236;
    wire N__50229;
    wire N__50226;
    wire N__50225;
    wire N__50224;
    wire N__50221;
    wire N__50218;
    wire N__50215;
    wire N__50212;
    wire N__50209;
    wire N__50206;
    wire N__50199;
    wire N__50196;
    wire N__50189;
    wire N__50186;
    wire N__50183;
    wire N__50180;
    wire N__50171;
    wire N__50170;
    wire N__50169;
    wire N__50168;
    wire N__50161;
    wire N__50156;
    wire N__50153;
    wire N__50150;
    wire N__50147;
    wire N__50144;
    wire N__50131;
    wire N__50128;
    wire N__50117;
    wire N__50114;
    wire N__50111;
    wire N__50108;
    wire N__50105;
    wire N__50100;
    wire N__50089;
    wire N__50072;
    wire N__50069;
    wire N__50066;
    wire N__50063;
    wire N__50062;
    wire N__50061;
    wire N__50060;
    wire N__50059;
    wire N__50058;
    wire N__50057;
    wire N__50056;
    wire N__50055;
    wire N__50054;
    wire N__50053;
    wire N__50052;
    wire N__50051;
    wire N__50050;
    wire N__50049;
    wire N__50048;
    wire N__50047;
    wire N__50044;
    wire N__50041;
    wire N__50038;
    wire N__50037;
    wire N__50036;
    wire N__50035;
    wire N__50034;
    wire N__50033;
    wire N__50032;
    wire N__50031;
    wire N__50030;
    wire N__50029;
    wire N__50028;
    wire N__50027;
    wire N__50024;
    wire N__50023;
    wire N__50020;
    wire N__50017;
    wire N__50016;
    wire N__50013;
    wire N__50010;
    wire N__50009;
    wire N__50006;
    wire N__50003;
    wire N__50000;
    wire N__49997;
    wire N__49996;
    wire N__49995;
    wire N__49994;
    wire N__49991;
    wire N__49990;
    wire N__49987;
    wire N__49984;
    wire N__49981;
    wire N__49978;
    wire N__49973;
    wire N__49970;
    wire N__49967;
    wire N__49964;
    wire N__49961;
    wire N__49958;
    wire N__49955;
    wire N__49952;
    wire N__49949;
    wire N__49946;
    wire N__49943;
    wire N__49940;
    wire N__49939;
    wire N__49936;
    wire N__49933;
    wire N__49930;
    wire N__49929;
    wire N__49926;
    wire N__49923;
    wire N__49920;
    wire N__49915;
    wire N__49912;
    wire N__49911;
    wire N__49910;
    wire N__49905;
    wire N__49900;
    wire N__49897;
    wire N__49894;
    wire N__49893;
    wire N__49892;
    wire N__49889;
    wire N__49886;
    wire N__49883;
    wire N__49880;
    wire N__49877;
    wire N__49876;
    wire N__49875;
    wire N__49874;
    wire N__49871;
    wire N__49868;
    wire N__49867;
    wire N__49866;
    wire N__49865;
    wire N__49848;
    wire N__49847;
    wire N__49838;
    wire N__49835;
    wire N__49834;
    wire N__49833;
    wire N__49832;
    wire N__49831;
    wire N__49828;
    wire N__49823;
    wire N__49820;
    wire N__49813;
    wire N__49808;
    wire N__49805;
    wire N__49802;
    wire N__49793;
    wire N__49790;
    wire N__49789;
    wire N__49784;
    wire N__49779;
    wire N__49774;
    wire N__49771;
    wire N__49768;
    wire N__49765;
    wire N__49760;
    wire N__49757;
    wire N__49754;
    wire N__49751;
    wire N__49748;
    wire N__49745;
    wire N__49740;
    wire N__49737;
    wire N__49734;
    wire N__49731;
    wire N__49728;
    wire N__49727;
    wire N__49726;
    wire N__49719;
    wire N__49710;
    wire N__49705;
    wire N__49702;
    wire N__49699;
    wire N__49690;
    wire N__49681;
    wire N__49678;
    wire N__49673;
    wire N__49672;
    wire N__49671;
    wire N__49662;
    wire N__49659;
    wire N__49656;
    wire N__49655;
    wire N__49654;
    wire N__49651;
    wire N__49648;
    wire N__49639;
    wire N__49636;
    wire N__49629;
    wire N__49626;
    wire N__49623;
    wire N__49616;
    wire N__49613;
    wire N__49610;
    wire N__49603;
    wire N__49586;
    wire N__49583;
    wire N__49580;
    wire N__49577;
    wire N__49576;
    wire N__49573;
    wire N__49570;
    wire N__49565;
    wire N__49562;
    wire N__49561;
    wire N__49558;
    wire N__49555;
    wire N__49550;
    wire N__49547;
    wire N__49544;
    wire N__49541;
    wire N__49538;
    wire N__49537;
    wire N__49536;
    wire N__49535;
    wire N__49534;
    wire N__49533;
    wire N__49532;
    wire N__49531;
    wire N__49530;
    wire N__49529;
    wire N__49528;
    wire N__49527;
    wire N__49526;
    wire N__49519;
    wire N__49510;
    wire N__49505;
    wire N__49496;
    wire N__49495;
    wire N__49494;
    wire N__49485;
    wire N__49484;
    wire N__49483;
    wire N__49480;
    wire N__49479;
    wire N__49476;
    wire N__49473;
    wire N__49470;
    wire N__49463;
    wire N__49462;
    wire N__49453;
    wire N__49450;
    wire N__49445;
    wire N__49442;
    wire N__49441;
    wire N__49440;
    wire N__49439;
    wire N__49438;
    wire N__49437;
    wire N__49436;
    wire N__49435;
    wire N__49434;
    wire N__49433;
    wire N__49432;
    wire N__49431;
    wire N__49430;
    wire N__49429;
    wire N__49428;
    wire N__49427;
    wire N__49426;
    wire N__49423;
    wire N__49420;
    wire N__49419;
    wire N__49418;
    wire N__49417;
    wire N__49414;
    wire N__49413;
    wire N__49410;
    wire N__49407;
    wire N__49406;
    wire N__49405;
    wire N__49404;
    wire N__49401;
    wire N__49400;
    wire N__49397;
    wire N__49394;
    wire N__49391;
    wire N__49390;
    wire N__49387;
    wire N__49386;
    wire N__49383;
    wire N__49382;
    wire N__49381;
    wire N__49372;
    wire N__49369;
    wire N__49366;
    wire N__49365;
    wire N__49364;
    wire N__49363;
    wire N__49362;
    wire N__49359;
    wire N__49356;
    wire N__49355;
    wire N__49354;
    wire N__49353;
    wire N__49352;
    wire N__49349;
    wire N__49338;
    wire N__49321;
    wire N__49318;
    wire N__49315;
    wire N__49308;
    wire N__49307;
    wire N__49306;
    wire N__49305;
    wire N__49304;
    wire N__49303;
    wire N__49302;
    wire N__49299;
    wire N__49296;
    wire N__49295;
    wire N__49294;
    wire N__49293;
    wire N__49292;
    wire N__49291;
    wire N__49290;
    wire N__49289;
    wire N__49288;
    wire N__49283;
    wire N__49280;
    wire N__49275;
    wire N__49272;
    wire N__49269;
    wire N__49264;
    wire N__49261;
    wire N__49260;
    wire N__49257;
    wire N__49254;
    wire N__49253;
    wire N__49250;
    wire N__49247;
    wire N__49246;
    wire N__49241;
    wire N__49240;
    wire N__49237;
    wire N__49234;
    wire N__49231;
    wire N__49224;
    wire N__49217;
    wire N__49212;
    wire N__49203;
    wire N__49194;
    wire N__49193;
    wire N__49192;
    wire N__49191;
    wire N__49188;
    wire N__49185;
    wire N__49182;
    wire N__49179;
    wire N__49176;
    wire N__49173;
    wire N__49170;
    wire N__49167;
    wire N__49164;
    wire N__49161;
    wire N__49158;
    wire N__49155;
    wire N__49152;
    wire N__49149;
    wire N__49146;
    wire N__49145;
    wire N__49142;
    wire N__49137;
    wire N__49124;
    wire N__49117;
    wire N__49116;
    wire N__49105;
    wire N__49102;
    wire N__49099;
    wire N__49096;
    wire N__49095;
    wire N__49088;
    wire N__49085;
    wire N__49082;
    wire N__49079;
    wire N__49076;
    wire N__49073;
    wire N__49064;
    wire N__49061;
    wire N__49058;
    wire N__49053;
    wire N__49050;
    wire N__49049;
    wire N__49046;
    wire N__49043;
    wire N__49040;
    wire N__49037;
    wire N__49034;
    wire N__49027;
    wire N__49024;
    wire N__49021;
    wire N__49018;
    wire N__49015;
    wire N__49012;
    wire N__49007;
    wire N__49004;
    wire N__49001;
    wire N__48994;
    wire N__48987;
    wire N__48984;
    wire N__48979;
    wire N__48972;
    wire N__48969;
    wire N__48962;
    wire N__48961;
    wire N__48960;
    wire N__48957;
    wire N__48956;
    wire N__48953;
    wire N__48952;
    wire N__48951;
    wire N__48950;
    wire N__48949;
    wire N__48948;
    wire N__48947;
    wire N__48946;
    wire N__48943;
    wire N__48940;
    wire N__48937;
    wire N__48936;
    wire N__48935;
    wire N__48934;
    wire N__48933;
    wire N__48932;
    wire N__48931;
    wire N__48930;
    wire N__48929;
    wire N__48926;
    wire N__48923;
    wire N__48912;
    wire N__48911;
    wire N__48910;
    wire N__48909;
    wire N__48908;
    wire N__48907;
    wire N__48904;
    wire N__48903;
    wire N__48902;
    wire N__48901;
    wire N__48900;
    wire N__48899;
    wire N__48898;
    wire N__48897;
    wire N__48894;
    wire N__48889;
    wire N__48872;
    wire N__48867;
    wire N__48864;
    wire N__48853;
    wire N__48850;
    wire N__48845;
    wire N__48834;
    wire N__48815;
    wire N__48812;
    wire N__48809;
    wire N__48806;
    wire N__48803;
    wire N__48802;
    wire N__48799;
    wire N__48796;
    wire N__48791;
    wire N__48790;
    wire N__48787;
    wire N__48784;
    wire N__48781;
    wire N__48776;
    wire N__48773;
    wire N__48772;
    wire N__48771;
    wire N__48766;
    wire N__48763;
    wire N__48760;
    wire N__48755;
    wire N__48754;
    wire N__48753;
    wire N__48752;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48734;
    wire N__48731;
    wire N__48730;
    wire N__48729;
    wire N__48722;
    wire N__48719;
    wire N__48718;
    wire N__48717;
    wire N__48714;
    wire N__48713;
    wire N__48708;
    wire N__48705;
    wire N__48702;
    wire N__48699;
    wire N__48692;
    wire N__48689;
    wire N__48686;
    wire N__48685;
    wire N__48682;
    wire N__48679;
    wire N__48676;
    wire N__48671;
    wire N__48668;
    wire N__48667;
    wire N__48666;
    wire N__48665;
    wire N__48662;
    wire N__48659;
    wire N__48656;
    wire N__48653;
    wire N__48650;
    wire N__48641;
    wire N__48638;
    wire N__48637;
    wire N__48636;
    wire N__48633;
    wire N__48628;
    wire N__48623;
    wire N__48620;
    wire N__48619;
    wire N__48618;
    wire N__48615;
    wire N__48612;
    wire N__48611;
    wire N__48608;
    wire N__48601;
    wire N__48596;
    wire N__48593;
    wire N__48592;
    wire N__48591;
    wire N__48588;
    wire N__48583;
    wire N__48578;
    wire N__48575;
    wire N__48572;
    wire N__48569;
    wire N__48568;
    wire N__48565;
    wire N__48562;
    wire N__48557;
    wire N__48554;
    wire N__48553;
    wire N__48550;
    wire N__48547;
    wire N__48544;
    wire N__48539;
    wire N__48536;
    wire N__48535;
    wire N__48534;
    wire N__48533;
    wire N__48530;
    wire N__48527;
    wire N__48522;
    wire N__48515;
    wire N__48512;
    wire N__48509;
    wire N__48506;
    wire N__48505;
    wire N__48502;
    wire N__48499;
    wire N__48496;
    wire N__48491;
    wire N__48490;
    wire N__48489;
    wire N__48488;
    wire N__48487;
    wire N__48486;
    wire N__48485;
    wire N__48484;
    wire N__48483;
    wire N__48482;
    wire N__48481;
    wire N__48480;
    wire N__48479;
    wire N__48478;
    wire N__48477;
    wire N__48476;
    wire N__48475;
    wire N__48474;
    wire N__48473;
    wire N__48472;
    wire N__48471;
    wire N__48470;
    wire N__48469;
    wire N__48468;
    wire N__48467;
    wire N__48466;
    wire N__48465;
    wire N__48464;
    wire N__48463;
    wire N__48462;
    wire N__48461;
    wire N__48460;
    wire N__48459;
    wire N__48458;
    wire N__48457;
    wire N__48456;
    wire N__48455;
    wire N__48454;
    wire N__48453;
    wire N__48452;
    wire N__48451;
    wire N__48450;
    wire N__48449;
    wire N__48448;
    wire N__48447;
    wire N__48446;
    wire N__48445;
    wire N__48444;
    wire N__48347;
    wire N__48344;
    wire N__48341;
    wire N__48338;
    wire N__48335;
    wire N__48332;
    wire N__48329;
    wire N__48328;
    wire N__48325;
    wire N__48324;
    wire N__48321;
    wire N__48318;
    wire N__48315;
    wire N__48310;
    wire N__48305;
    wire N__48304;
    wire N__48303;
    wire N__48300;
    wire N__48297;
    wire N__48294;
    wire N__48289;
    wire N__48284;
    wire N__48281;
    wire N__48278;
    wire N__48275;
    wire N__48272;
    wire N__48269;
    wire N__48266;
    wire N__48265;
    wire N__48264;
    wire N__48263;
    wire N__48262;
    wire N__48261;
    wire N__48260;
    wire N__48259;
    wire N__48242;
    wire N__48239;
    wire N__48236;
    wire N__48233;
    wire N__48232;
    wire N__48231;
    wire N__48228;
    wire N__48225;
    wire N__48222;
    wire N__48219;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48207;
    wire N__48204;
    wire N__48201;
    wire N__48198;
    wire N__48191;
    wire N__48188;
    wire N__48185;
    wire N__48182;
    wire N__48179;
    wire N__48176;
    wire N__48173;
    wire N__48170;
    wire N__48167;
    wire N__48164;
    wire N__48161;
    wire N__48158;
    wire N__48155;
    wire N__48152;
    wire N__48149;
    wire N__48146;
    wire N__48143;
    wire N__48140;
    wire N__48137;
    wire N__48134;
    wire N__48131;
    wire N__48130;
    wire N__48129;
    wire N__48128;
    wire N__48127;
    wire N__48126;
    wire N__48119;
    wire N__48116;
    wire N__48113;
    wire N__48110;
    wire N__48103;
    wire N__48098;
    wire N__48097;
    wire N__48094;
    wire N__48091;
    wire N__48090;
    wire N__48089;
    wire N__48086;
    wire N__48079;
    wire N__48074;
    wire N__48073;
    wire N__48070;
    wire N__48067;
    wire N__48062;
    wire N__48059;
    wire N__48056;
    wire N__48053;
    wire N__48052;
    wire N__48051;
    wire N__48048;
    wire N__48045;
    wire N__48042;
    wire N__48041;
    wire N__48038;
    wire N__48033;
    wire N__48032;
    wire N__48029;
    wire N__48024;
    wire N__48021;
    wire N__48018;
    wire N__48015;
    wire N__48012;
    wire N__48011;
    wire N__48008;
    wire N__48007;
    wire N__48006;
    wire N__48001;
    wire N__47998;
    wire N__47995;
    wire N__47992;
    wire N__47989;
    wire N__47984;
    wire N__47977;
    wire N__47974;
    wire N__47971;
    wire N__47968;
    wire N__47965;
    wire N__47962;
    wire N__47957;
    wire N__47956;
    wire N__47951;
    wire N__47948;
    wire N__47947;
    wire N__47944;
    wire N__47941;
    wire N__47936;
    wire N__47933;
    wire N__47930;
    wire N__47929;
    wire N__47928;
    wire N__47925;
    wire N__47922;
    wire N__47919;
    wire N__47912;
    wire N__47909;
    wire N__47906;
    wire N__47903;
    wire N__47900;
    wire N__47897;
    wire N__47894;
    wire N__47893;
    wire N__47892;
    wire N__47889;
    wire N__47888;
    wire N__47887;
    wire N__47882;
    wire N__47879;
    wire N__47876;
    wire N__47873;
    wire N__47870;
    wire N__47867;
    wire N__47864;
    wire N__47861;
    wire N__47858;
    wire N__47855;
    wire N__47852;
    wire N__47849;
    wire N__47846;
    wire N__47839;
    wire N__47834;
    wire N__47831;
    wire N__47828;
    wire N__47825;
    wire N__47822;
    wire N__47819;
    wire N__47816;
    wire N__47813;
    wire N__47810;
    wire N__47807;
    wire N__47804;
    wire N__47801;
    wire N__47798;
    wire N__47795;
    wire N__47792;
    wire N__47789;
    wire N__47786;
    wire N__47783;
    wire N__47782;
    wire N__47779;
    wire N__47776;
    wire N__47773;
    wire N__47770;
    wire N__47765;
    wire N__47762;
    wire N__47759;
    wire N__47756;
    wire N__47753;
    wire N__47750;
    wire N__47747;
    wire N__47744;
    wire N__47741;
    wire N__47738;
    wire N__47735;
    wire N__47732;
    wire N__47729;
    wire N__47726;
    wire N__47723;
    wire N__47720;
    wire N__47717;
    wire N__47714;
    wire N__47711;
    wire N__47708;
    wire N__47705;
    wire N__47702;
    wire N__47699;
    wire N__47696;
    wire N__47693;
    wire N__47690;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47675;
    wire N__47672;
    wire N__47669;
    wire N__47666;
    wire N__47663;
    wire N__47660;
    wire N__47657;
    wire N__47654;
    wire N__47651;
    wire N__47648;
    wire N__47645;
    wire N__47642;
    wire N__47639;
    wire N__47636;
    wire N__47633;
    wire N__47630;
    wire N__47627;
    wire N__47624;
    wire N__47621;
    wire N__47618;
    wire N__47615;
    wire N__47612;
    wire N__47609;
    wire N__47606;
    wire N__47603;
    wire N__47600;
    wire N__47597;
    wire N__47594;
    wire N__47591;
    wire N__47588;
    wire N__47585;
    wire N__47582;
    wire N__47579;
    wire N__47576;
    wire N__47573;
    wire N__47570;
    wire N__47567;
    wire N__47564;
    wire N__47561;
    wire N__47558;
    wire N__47555;
    wire N__47554;
    wire N__47549;
    wire N__47546;
    wire N__47545;
    wire N__47542;
    wire N__47539;
    wire N__47536;
    wire N__47533;
    wire N__47530;
    wire N__47525;
    wire N__47522;
    wire N__47519;
    wire N__47516;
    wire N__47513;
    wire N__47512;
    wire N__47511;
    wire N__47508;
    wire N__47507;
    wire N__47506;
    wire N__47503;
    wire N__47502;
    wire N__47501;
    wire N__47500;
    wire N__47499;
    wire N__47498;
    wire N__47497;
    wire N__47496;
    wire N__47493;
    wire N__47492;
    wire N__47489;
    wire N__47486;
    wire N__47485;
    wire N__47484;
    wire N__47483;
    wire N__47482;
    wire N__47481;
    wire N__47480;
    wire N__47477;
    wire N__47474;
    wire N__47471;
    wire N__47468;
    wire N__47465;
    wire N__47462;
    wire N__47461;
    wire N__47460;
    wire N__47459;
    wire N__47458;
    wire N__47457;
    wire N__47454;
    wire N__47451;
    wire N__47448;
    wire N__47447;
    wire N__47446;
    wire N__47443;
    wire N__47440;
    wire N__47439;
    wire N__47438;
    wire N__47437;
    wire N__47432;
    wire N__47429;
    wire N__47426;
    wire N__47423;
    wire N__47420;
    wire N__47417;
    wire N__47414;
    wire N__47413;
    wire N__47410;
    wire N__47399;
    wire N__47396;
    wire N__47395;
    wire N__47394;
    wire N__47393;
    wire N__47390;
    wire N__47387;
    wire N__47384;
    wire N__47381;
    wire N__47380;
    wire N__47379;
    wire N__47374;
    wire N__47371;
    wire N__47368;
    wire N__47365;
    wire N__47364;
    wire N__47363;
    wire N__47358;
    wire N__47355;
    wire N__47352;
    wire N__47349;
    wire N__47348;
    wire N__47347;
    wire N__47346;
    wire N__47345;
    wire N__47344;
    wire N__47343;
    wire N__47330;
    wire N__47329;
    wire N__47328;
    wire N__47325;
    wire N__47322;
    wire N__47315;
    wire N__47312;
    wire N__47309;
    wire N__47306;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47282;
    wire N__47279;
    wire N__47276;
    wire N__47275;
    wire N__47272;
    wire N__47267;
    wire N__47264;
    wire N__47261;
    wire N__47258;
    wire N__47255;
    wire N__47252;
    wire N__47251;
    wire N__47248;
    wire N__47247;
    wire N__47246;
    wire N__47245;
    wire N__47244;
    wire N__47241;
    wire N__47238;
    wire N__47235;
    wire N__47232;
    wire N__47229;
    wire N__47224;
    wire N__47215;
    wire N__47210;
    wire N__47203;
    wire N__47202;
    wire N__47195;
    wire N__47192;
    wire N__47189;
    wire N__47178;
    wire N__47175;
    wire N__47174;
    wire N__47171;
    wire N__47170;
    wire N__47169;
    wire N__47166;
    wire N__47163;
    wire N__47160;
    wire N__47157;
    wire N__47154;
    wire N__47149;
    wire N__47144;
    wire N__47141;
    wire N__47138;
    wire N__47135;
    wire N__47130;
    wire N__47127;
    wire N__47122;
    wire N__47121;
    wire N__47120;
    wire N__47119;
    wire N__47118;
    wire N__47115;
    wire N__47110;
    wire N__47107;
    wire N__47104;
    wire N__47101;
    wire N__47098;
    wire N__47087;
    wire N__47080;
    wire N__47075;
    wire N__47070;
    wire N__47067;
    wire N__47064;
    wire N__47061;
    wire N__47058;
    wire N__47055;
    wire N__47048;
    wire N__47039;
    wire N__47018;
    wire N__47017;
    wire N__47014;
    wire N__47011;
    wire N__47006;
    wire N__47003;
    wire N__47000;
    wire N__46999;
    wire N__46996;
    wire N__46993;
    wire N__46988;
    wire N__46985;
    wire N__46982;
    wire N__46979;
    wire N__46976;
    wire N__46973;
    wire N__46970;
    wire N__46967;
    wire N__46964;
    wire N__46963;
    wire N__46962;
    wire N__46961;
    wire N__46960;
    wire N__46959;
    wire N__46958;
    wire N__46957;
    wire N__46956;
    wire N__46953;
    wire N__46944;
    wire N__46935;
    wire N__46932;
    wire N__46925;
    wire N__46924;
    wire N__46923;
    wire N__46922;
    wire N__46921;
    wire N__46920;
    wire N__46919;
    wire N__46916;
    wire N__46915;
    wire N__46914;
    wire N__46913;
    wire N__46910;
    wire N__46909;
    wire N__46908;
    wire N__46907;
    wire N__46906;
    wire N__46905;
    wire N__46902;
    wire N__46901;
    wire N__46898;
    wire N__46895;
    wire N__46892;
    wire N__46891;
    wire N__46888;
    wire N__46885;
    wire N__46882;
    wire N__46879;
    wire N__46876;
    wire N__46873;
    wire N__46870;
    wire N__46867;
    wire N__46866;
    wire N__46863;
    wire N__46860;
    wire N__46859;
    wire N__46858;
    wire N__46857;
    wire N__46856;
    wire N__46855;
    wire N__46854;
    wire N__46853;
    wire N__46852;
    wire N__46851;
    wire N__46848;
    wire N__46847;
    wire N__46844;
    wire N__46841;
    wire N__46840;
    wire N__46833;
    wire N__46830;
    wire N__46829;
    wire N__46826;
    wire N__46817;
    wire N__46810;
    wire N__46807;
    wire N__46804;
    wire N__46801;
    wire N__46798;
    wire N__46795;
    wire N__46794;
    wire N__46793;
    wire N__46790;
    wire N__46789;
    wire N__46786;
    wire N__46783;
    wire N__46780;
    wire N__46779;
    wire N__46776;
    wire N__46775;
    wire N__46774;
    wire N__46771;
    wire N__46770;
    wire N__46769;
    wire N__46766;
    wire N__46765;
    wire N__46764;
    wire N__46763;
    wire N__46762;
    wire N__46759;
    wire N__46756;
    wire N__46753;
    wire N__46752;
    wire N__46751;
    wire N__46750;
    wire N__46747;
    wire N__46746;
    wire N__46743;
    wire N__46738;
    wire N__46735;
    wire N__46726;
    wire N__46719;
    wire N__46716;
    wire N__46713;
    wire N__46710;
    wire N__46709;
    wire N__46708;
    wire N__46707;
    wire N__46704;
    wire N__46701;
    wire N__46696;
    wire N__46693;
    wire N__46690;
    wire N__46689;
    wire N__46686;
    wire N__46683;
    wire N__46680;
    wire N__46677;
    wire N__46674;
    wire N__46671;
    wire N__46668;
    wire N__46665;
    wire N__46662;
    wire N__46659;
    wire N__46656;
    wire N__46651;
    wire N__46650;
    wire N__46647;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46635;
    wire N__46632;
    wire N__46629;
    wire N__46624;
    wire N__46621;
    wire N__46614;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46604;
    wire N__46603;
    wire N__46600;
    wire N__46599;
    wire N__46598;
    wire N__46593;
    wire N__46586;
    wire N__46583;
    wire N__46572;
    wire N__46569;
    wire N__46566;
    wire N__46557;
    wire N__46554;
    wire N__46551;
    wire N__46538;
    wire N__46533;
    wire N__46522;
    wire N__46521;
    wire N__46520;
    wire N__46519;
    wire N__46518;
    wire N__46515;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46494;
    wire N__46491;
    wire N__46478;
    wire N__46475;
    wire N__46472;
    wire N__46469;
    wire N__46466;
    wire N__46463;
    wire N__46458;
    wire N__46449;
    wire N__46430;
    wire N__46427;
    wire N__46424;
    wire N__46421;
    wire N__46420;
    wire N__46417;
    wire N__46414;
    wire N__46409;
    wire N__46408;
    wire N__46405;
    wire N__46402;
    wire N__46397;
    wire N__46394;
    wire N__46391;
    wire N__46390;
    wire N__46389;
    wire N__46388;
    wire N__46387;
    wire N__46386;
    wire N__46385;
    wire N__46384;
    wire N__46383;
    wire N__46382;
    wire N__46381;
    wire N__46380;
    wire N__46379;
    wire N__46376;
    wire N__46375;
    wire N__46374;
    wire N__46371;
    wire N__46368;
    wire N__46365;
    wire N__46362;
    wire N__46359;
    wire N__46356;
    wire N__46353;
    wire N__46352;
    wire N__46349;
    wire N__46346;
    wire N__46345;
    wire N__46344;
    wire N__46343;
    wire N__46342;
    wire N__46339;
    wire N__46338;
    wire N__46335;
    wire N__46332;
    wire N__46331;
    wire N__46328;
    wire N__46325;
    wire N__46324;
    wire N__46323;
    wire N__46322;
    wire N__46321;
    wire N__46318;
    wire N__46317;
    wire N__46316;
    wire N__46315;
    wire N__46314;
    wire N__46309;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46293;
    wire N__46288;
    wire N__46285;
    wire N__46282;
    wire N__46281;
    wire N__46280;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46270;
    wire N__46267;
    wire N__46262;
    wire N__46259;
    wire N__46254;
    wire N__46251;
    wire N__46248;
    wire N__46245;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46235;
    wire N__46234;
    wire N__46233;
    wire N__46230;
    wire N__46227;
    wire N__46224;
    wire N__46215;
    wire N__46212;
    wire N__46211;
    wire N__46210;
    wire N__46209;
    wire N__46202;
    wire N__46199;
    wire N__46196;
    wire N__46193;
    wire N__46184;
    wire N__46179;
    wire N__46174;
    wire N__46167;
    wire N__46162;
    wire N__46159;
    wire N__46156;
    wire N__46153;
    wire N__46150;
    wire N__46149;
    wire N__46148;
    wire N__46147;
    wire N__46146;
    wire N__46145;
    wire N__46144;
    wire N__46143;
    wire N__46142;
    wire N__46141;
    wire N__46136;
    wire N__46131;
    wire N__46130;
    wire N__46127;
    wire N__46124;
    wire N__46121;
    wire N__46118;
    wire N__46115;
    wire N__46106;
    wire N__46101;
    wire N__46098;
    wire N__46093;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46081;
    wire N__46078;
    wire N__46075;
    wire N__46072;
    wire N__46069;
    wire N__46066;
    wire N__46063;
    wire N__46060;
    wire N__46055;
    wire N__46054;
    wire N__46053;
    wire N__46052;
    wire N__46051;
    wire N__46050;
    wire N__46047;
    wire N__46044;
    wire N__46043;
    wire N__46042;
    wire N__46039;
    wire N__46034;
    wire N__46029;
    wire N__46022;
    wire N__46019;
    wire N__46016;
    wire N__46015;
    wire N__46010;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45990;
    wire N__45987;
    wire N__45980;
    wire N__45979;
    wire N__45978;
    wire N__45977;
    wire N__45974;
    wire N__45969;
    wire N__45966;
    wire N__45963;
    wire N__45956;
    wire N__45953;
    wire N__45948;
    wire N__45945;
    wire N__45942;
    wire N__45935;
    wire N__45932;
    wire N__45927;
    wire N__45924;
    wire N__45921;
    wire N__45918;
    wire N__45911;
    wire N__45908;
    wire N__45905;
    wire N__45900;
    wire N__45889;
    wire N__45872;
    wire N__45869;
    wire N__45866;
    wire N__45863;
    wire N__45860;
    wire N__45857;
    wire N__45856;
    wire N__45853;
    wire N__45850;
    wire N__45845;
    wire N__45844;
    wire N__45841;
    wire N__45838;
    wire N__45835;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45818;
    wire N__45815;
    wire N__45812;
    wire N__45809;
    wire N__45806;
    wire N__45803;
    wire N__45800;
    wire N__45797;
    wire N__45794;
    wire N__45791;
    wire N__45788;
    wire N__45785;
    wire N__45782;
    wire N__45779;
    wire N__45776;
    wire N__45773;
    wire N__45772;
    wire N__45771;
    wire N__45768;
    wire N__45765;
    wire N__45762;
    wire N__45757;
    wire N__45752;
    wire N__45751;
    wire N__45748;
    wire N__45745;
    wire N__45744;
    wire N__45743;
    wire N__45740;
    wire N__45737;
    wire N__45732;
    wire N__45727;
    wire N__45722;
    wire N__45719;
    wire N__45718;
    wire N__45717;
    wire N__45716;
    wire N__45715;
    wire N__45714;
    wire N__45711;
    wire N__45698;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45686;
    wire N__45683;
    wire N__45680;
    wire N__45677;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45656;
    wire N__45653;
    wire N__45650;
    wire N__45647;
    wire N__45644;
    wire N__45641;
    wire N__45638;
    wire N__45635;
    wire N__45632;
    wire N__45629;
    wire N__45626;
    wire N__45623;
    wire N__45620;
    wire N__45617;
    wire N__45614;
    wire N__45611;
    wire N__45608;
    wire N__45607;
    wire N__45606;
    wire N__45605;
    wire N__45604;
    wire N__45603;
    wire N__45602;
    wire N__45601;
    wire N__45600;
    wire N__45597;
    wire N__45594;
    wire N__45593;
    wire N__45592;
    wire N__45589;
    wire N__45586;
    wire N__45585;
    wire N__45582;
    wire N__45581;
    wire N__45580;
    wire N__45579;
    wire N__45578;
    wire N__45577;
    wire N__45576;
    wire N__45575;
    wire N__45574;
    wire N__45571;
    wire N__45570;
    wire N__45569;
    wire N__45568;
    wire N__45567;
    wire N__45564;
    wire N__45563;
    wire N__45562;
    wire N__45561;
    wire N__45560;
    wire N__45559;
    wire N__45558;
    wire N__45555;
    wire N__45554;
    wire N__45551;
    wire N__45546;
    wire N__45543;
    wire N__45540;
    wire N__45535;
    wire N__45532;
    wire N__45531;
    wire N__45530;
    wire N__45529;
    wire N__45528;
    wire N__45525;
    wire N__45522;
    wire N__45519;
    wire N__45516;
    wire N__45513;
    wire N__45510;
    wire N__45509;
    wire N__45508;
    wire N__45507;
    wire N__45506;
    wire N__45503;
    wire N__45500;
    wire N__45497;
    wire N__45494;
    wire N__45491;
    wire N__45488;
    wire N__45485;
    wire N__45482;
    wire N__45481;
    wire N__45478;
    wire N__45475;
    wire N__45472;
    wire N__45469;
    wire N__45466;
    wire N__45463;
    wire N__45460;
    wire N__45457;
    wire N__45454;
    wire N__45451;
    wire N__45444;
    wire N__45439;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45414;
    wire N__45413;
    wire N__45412;
    wire N__45411;
    wire N__45410;
    wire N__45407;
    wire N__45404;
    wire N__45401;
    wire N__45398;
    wire N__45397;
    wire N__45394;
    wire N__45389;
    wire N__45388;
    wire N__45387;
    wire N__45384;
    wire N__45375;
    wire N__45374;
    wire N__45373;
    wire N__45372;
    wire N__45369;
    wire N__45360;
    wire N__45359;
    wire N__45354;
    wire N__45351;
    wire N__45350;
    wire N__45349;
    wire N__45348;
    wire N__45343;
    wire N__45338;
    wire N__45333;
    wire N__45326;
    wire N__45323;
    wire N__45320;
    wire N__45317;
    wire N__45314;
    wire N__45311;
    wire N__45308;
    wire N__45301;
    wire N__45298;
    wire N__45297;
    wire N__45296;
    wire N__45291;
    wire N__45288;
    wire N__45285;
    wire N__45280;
    wire N__45277;
    wire N__45274;
    wire N__45271;
    wire N__45268;
    wire N__45265;
    wire N__45262;
    wire N__45257;
    wire N__45254;
    wire N__45251;
    wire N__45248;
    wire N__45245;
    wire N__45238;
    wire N__45227;
    wire N__45226;
    wire N__45225;
    wire N__45224;
    wire N__45221;
    wire N__45218;
    wire N__45215;
    wire N__45212;
    wire N__45209;
    wire N__45202;
    wire N__45191;
    wire N__45178;
    wire N__45171;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45147;
    wire N__45134;
    wire N__45131;
    wire N__45128;
    wire N__45125;
    wire N__45122;
    wire N__45119;
    wire N__45118;
    wire N__45117;
    wire N__45116;
    wire N__45115;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45107;
    wire N__45106;
    wire N__45105;
    wire N__45104;
    wire N__45103;
    wire N__45102;
    wire N__45101;
    wire N__45100;
    wire N__45097;
    wire N__45096;
    wire N__45095;
    wire N__45094;
    wire N__45091;
    wire N__45090;
    wire N__45089;
    wire N__45086;
    wire N__45085;
    wire N__45082;
    wire N__45081;
    wire N__45080;
    wire N__45079;
    wire N__45078;
    wire N__45077;
    wire N__45072;
    wire N__45069;
    wire N__45068;
    wire N__45067;
    wire N__45066;
    wire N__45065;
    wire N__45064;
    wire N__45061;
    wire N__45058;
    wire N__45057;
    wire N__45056;
    wire N__45055;
    wire N__45054;
    wire N__45053;
    wire N__45050;
    wire N__45047;
    wire N__45044;
    wire N__45041;
    wire N__45038;
    wire N__45037;
    wire N__45034;
    wire N__45031;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45013;
    wire N__45010;
    wire N__45009;
    wire N__45006;
    wire N__45005;
    wire N__45002;
    wire N__45001;
    wire N__45000;
    wire N__44997;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44983;
    wire N__44982;
    wire N__44981;
    wire N__44980;
    wire N__44977;
    wire N__44974;
    wire N__44971;
    wire N__44968;
    wire N__44965;
    wire N__44962;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44952;
    wire N__44951;
    wire N__44948;
    wire N__44945;
    wire N__44942;
    wire N__44939;
    wire N__44930;
    wire N__44929;
    wire N__44928;
    wire N__44925;
    wire N__44924;
    wire N__44923;
    wire N__44920;
    wire N__44915;
    wire N__44908;
    wire N__44905;
    wire N__44902;
    wire N__44899;
    wire N__44896;
    wire N__44893;
    wire N__44890;
    wire N__44887;
    wire N__44884;
    wire N__44881;
    wire N__44876;
    wire N__44871;
    wire N__44868;
    wire N__44867;
    wire N__44864;
    wire N__44861;
    wire N__44858;
    wire N__44853;
    wire N__44842;
    wire N__44841;
    wire N__44840;
    wire N__44835;
    wire N__44834;
    wire N__44833;
    wire N__44830;
    wire N__44827;
    wire N__44820;
    wire N__44815;
    wire N__44812;
    wire N__44809;
    wire N__44806;
    wire N__44803;
    wire N__44800;
    wire N__44793;
    wire N__44788;
    wire N__44781;
    wire N__44774;
    wire N__44771;
    wire N__44764;
    wire N__44763;
    wire N__44760;
    wire N__44753;
    wire N__44748;
    wire N__44745;
    wire N__44742;
    wire N__44739;
    wire N__44734;
    wire N__44733;
    wire N__44732;
    wire N__44731;
    wire N__44730;
    wire N__44727;
    wire N__44720;
    wire N__44707;
    wire N__44702;
    wire N__44699;
    wire N__44694;
    wire N__44691;
    wire N__44684;
    wire N__44675;
    wire N__44672;
    wire N__44669;
    wire N__44666;
    wire N__44663;
    wire N__44656;
    wire N__44653;
    wire N__44648;
    wire N__44641;
    wire N__44624;
    wire N__44621;
    wire N__44618;
    wire N__44615;
    wire N__44612;
    wire N__44609;
    wire N__44606;
    wire N__44603;
    wire N__44600;
    wire N__44597;
    wire N__44594;
    wire N__44591;
    wire N__44588;
    wire N__44585;
    wire N__44582;
    wire N__44579;
    wire N__44576;
    wire N__44573;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44561;
    wire N__44558;
    wire N__44557;
    wire N__44554;
    wire N__44551;
    wire N__44548;
    wire N__44543;
    wire N__44540;
    wire N__44537;
    wire N__44534;
    wire N__44531;
    wire N__44528;
    wire N__44525;
    wire N__44522;
    wire N__44519;
    wire N__44516;
    wire N__44513;
    wire N__44510;
    wire N__44507;
    wire N__44504;
    wire N__44501;
    wire N__44498;
    wire N__44495;
    wire N__44492;
    wire N__44489;
    wire N__44486;
    wire N__44483;
    wire N__44480;
    wire N__44477;
    wire N__44474;
    wire N__44471;
    wire N__44468;
    wire N__44465;
    wire N__44462;
    wire N__44459;
    wire N__44456;
    wire N__44453;
    wire N__44450;
    wire N__44447;
    wire N__44444;
    wire N__44441;
    wire N__44438;
    wire N__44435;
    wire N__44432;
    wire N__44429;
    wire N__44426;
    wire N__44423;
    wire N__44420;
    wire N__44417;
    wire N__44414;
    wire N__44411;
    wire N__44408;
    wire N__44405;
    wire N__44402;
    wire N__44399;
    wire N__44396;
    wire N__44393;
    wire N__44390;
    wire N__44387;
    wire N__44384;
    wire N__44381;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44366;
    wire N__44363;
    wire N__44360;
    wire N__44357;
    wire N__44354;
    wire N__44351;
    wire N__44348;
    wire N__44345;
    wire N__44342;
    wire N__44339;
    wire N__44336;
    wire N__44333;
    wire N__44330;
    wire N__44327;
    wire N__44324;
    wire N__44321;
    wire N__44318;
    wire N__44315;
    wire N__44312;
    wire N__44309;
    wire N__44306;
    wire N__44303;
    wire N__44300;
    wire N__44297;
    wire N__44294;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44279;
    wire N__44278;
    wire N__44275;
    wire N__44272;
    wire N__44267;
    wire N__44264;
    wire N__44261;
    wire N__44258;
    wire N__44255;
    wire N__44252;
    wire N__44249;
    wire N__44246;
    wire N__44245;
    wire N__44244;
    wire N__44243;
    wire N__44240;
    wire N__44239;
    wire N__44238;
    wire N__44237;
    wire N__44234;
    wire N__44231;
    wire N__44228;
    wire N__44225;
    wire N__44224;
    wire N__44221;
    wire N__44218;
    wire N__44215;
    wire N__44212;
    wire N__44209;
    wire N__44206;
    wire N__44203;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44191;
    wire N__44184;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44170;
    wire N__44167;
    wire N__44164;
    wire N__44161;
    wire N__44158;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44144;
    wire N__44135;
    wire N__44132;
    wire N__44129;
    wire N__44126;
    wire N__44123;
    wire N__44120;
    wire N__44117;
    wire N__44114;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44099;
    wire N__44096;
    wire N__44093;
    wire N__44090;
    wire N__44087;
    wire N__44084;
    wire N__44081;
    wire N__44078;
    wire N__44075;
    wire N__44072;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44060;
    wire N__44057;
    wire N__44056;
    wire N__44053;
    wire N__44050;
    wire N__44045;
    wire N__44042;
    wire N__44039;
    wire N__44036;
    wire N__44033;
    wire N__44032;
    wire N__44029;
    wire N__44026;
    wire N__44023;
    wire N__44020;
    wire N__44015;
    wire N__44012;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__44000;
    wire N__43999;
    wire N__43996;
    wire N__43993;
    wire N__43988;
    wire N__43985;
    wire N__43982;
    wire N__43979;
    wire N__43976;
    wire N__43975;
    wire N__43972;
    wire N__43969;
    wire N__43966;
    wire N__43963;
    wire N__43958;
    wire N__43957;
    wire N__43956;
    wire N__43955;
    wire N__43954;
    wire N__43953;
    wire N__43952;
    wire N__43951;
    wire N__43950;
    wire N__43949;
    wire N__43948;
    wire N__43947;
    wire N__43922;
    wire N__43919;
    wire N__43916;
    wire N__43913;
    wire N__43910;
    wire N__43907;
    wire N__43904;
    wire N__43903;
    wire N__43902;
    wire N__43901;
    wire N__43898;
    wire N__43895;
    wire N__43892;
    wire N__43889;
    wire N__43888;
    wire N__43883;
    wire N__43880;
    wire N__43877;
    wire N__43874;
    wire N__43871;
    wire N__43868;
    wire N__43865;
    wire N__43862;
    wire N__43853;
    wire N__43850;
    wire N__43847;
    wire N__43844;
    wire N__43841;
    wire N__43838;
    wire N__43835;
    wire N__43832;
    wire N__43829;
    wire N__43826;
    wire N__43823;
    wire N__43820;
    wire N__43817;
    wire N__43814;
    wire N__43811;
    wire N__43808;
    wire N__43805;
    wire N__43802;
    wire N__43799;
    wire N__43796;
    wire N__43793;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43781;
    wire N__43778;
    wire N__43775;
    wire N__43772;
    wire N__43771;
    wire N__43770;
    wire N__43769;
    wire N__43768;
    wire N__43767;
    wire N__43766;
    wire N__43765;
    wire N__43762;
    wire N__43759;
    wire N__43756;
    wire N__43751;
    wire N__43748;
    wire N__43737;
    wire N__43736;
    wire N__43735;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43714;
    wire N__43709;
    wire N__43700;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43688;
    wire N__43687;
    wire N__43686;
    wire N__43683;
    wire N__43680;
    wire N__43677;
    wire N__43674;
    wire N__43671;
    wire N__43668;
    wire N__43661;
    wire N__43658;
    wire N__43655;
    wire N__43652;
    wire N__43649;
    wire N__43646;
    wire N__43645;
    wire N__43642;
    wire N__43639;
    wire N__43634;
    wire N__43631;
    wire N__43628;
    wire N__43625;
    wire N__43622;
    wire N__43621;
    wire N__43618;
    wire N__43615;
    wire N__43610;
    wire N__43607;
    wire N__43604;
    wire N__43601;
    wire N__43598;
    wire N__43595;
    wire N__43592;
    wire N__43589;
    wire N__43586;
    wire N__43583;
    wire N__43580;
    wire N__43577;
    wire N__43574;
    wire N__43573;
    wire N__43570;
    wire N__43567;
    wire N__43562;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43538;
    wire N__43535;
    wire N__43532;
    wire N__43529;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43517;
    wire N__43514;
    wire N__43511;
    wire N__43510;
    wire N__43507;
    wire N__43504;
    wire N__43499;
    wire N__43498;
    wire N__43497;
    wire N__43496;
    wire N__43495;
    wire N__43494;
    wire N__43493;
    wire N__43492;
    wire N__43491;
    wire N__43490;
    wire N__43489;
    wire N__43488;
    wire N__43487;
    wire N__43478;
    wire N__43469;
    wire N__43468;
    wire N__43467;
    wire N__43466;
    wire N__43463;
    wire N__43462;
    wire N__43459;
    wire N__43458;
    wire N__43455;
    wire N__43454;
    wire N__43451;
    wire N__43450;
    wire N__43447;
    wire N__43446;
    wire N__43445;
    wire N__43440;
    wire N__43439;
    wire N__43438;
    wire N__43433;
    wire N__43430;
    wire N__43413;
    wire N__43408;
    wire N__43405;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43385;
    wire N__43376;
    wire N__43373;
    wire N__43370;
    wire N__43367;
    wire N__43366;
    wire N__43363;
    wire N__43360;
    wire N__43355;
    wire N__43354;
    wire N__43353;
    wire N__43352;
    wire N__43351;
    wire N__43350;
    wire N__43349;
    wire N__43348;
    wire N__43347;
    wire N__43346;
    wire N__43345;
    wire N__43344;
    wire N__43343;
    wire N__43342;
    wire N__43341;
    wire N__43340;
    wire N__43339;
    wire N__43338;
    wire N__43337;
    wire N__43336;
    wire N__43335;
    wire N__43334;
    wire N__43317;
    wire N__43316;
    wire N__43315;
    wire N__43308;
    wire N__43291;
    wire N__43286;
    wire N__43283;
    wire N__43280;
    wire N__43277;
    wire N__43274;
    wire N__43265;
    wire N__43262;
    wire N__43255;
    wire N__43252;
    wire N__43249;
    wire N__43244;
    wire N__43241;
    wire N__43238;
    wire N__43235;
    wire N__43232;
    wire N__43229;
    wire N__43226;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43218;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43193;
    wire N__43190;
    wire N__43187;
    wire N__43184;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43172;
    wire N__43169;
    wire N__43166;
    wire N__43163;
    wire N__43160;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43150;
    wire N__43147;
    wire N__43142;
    wire N__43139;
    wire N__43136;
    wire N__43133;
    wire N__43130;
    wire N__43127;
    wire N__43126;
    wire N__43123;
    wire N__43120;
    wire N__43115;
    wire N__43112;
    wire N__43109;
    wire N__43106;
    wire N__43103;
    wire N__43100;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43087;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43073;
    wire N__43070;
    wire N__43069;
    wire N__43066;
    wire N__43063;
    wire N__43060;
    wire N__43055;
    wire N__43052;
    wire N__43049;
    wire N__43046;
    wire N__43043;
    wire N__43042;
    wire N__43039;
    wire N__43036;
    wire N__43033;
    wire N__43028;
    wire N__43025;
    wire N__43022;
    wire N__43019;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43007;
    wire N__43004;
    wire N__43001;
    wire N__42998;
    wire N__42995;
    wire N__42992;
    wire N__42989;
    wire N__42986;
    wire N__42983;
    wire N__42980;
    wire N__42977;
    wire N__42974;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42941;
    wire N__42938;
    wire N__42935;
    wire N__42932;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42914;
    wire N__42911;
    wire N__42908;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42896;
    wire N__42893;
    wire N__42890;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42857;
    wire N__42854;
    wire N__42851;
    wire N__42848;
    wire N__42845;
    wire N__42842;
    wire N__42839;
    wire N__42836;
    wire N__42833;
    wire N__42830;
    wire N__42827;
    wire N__42824;
    wire N__42821;
    wire N__42818;
    wire N__42815;
    wire N__42812;
    wire N__42809;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42794;
    wire N__42791;
    wire N__42788;
    wire N__42787;
    wire N__42784;
    wire N__42781;
    wire N__42776;
    wire N__42773;
    wire N__42772;
    wire N__42769;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42759;
    wire N__42756;
    wire N__42753;
    wire N__42746;
    wire N__42743;
    wire N__42740;
    wire N__42737;
    wire N__42736;
    wire N__42733;
    wire N__42730;
    wire N__42729;
    wire N__42726;
    wire N__42723;
    wire N__42720;
    wire N__42717;
    wire N__42710;
    wire N__42707;
    wire N__42706;
    wire N__42705;
    wire N__42702;
    wire N__42697;
    wire N__42692;
    wire N__42689;
    wire N__42686;
    wire N__42683;
    wire N__42680;
    wire N__42679;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42659;
    wire N__42656;
    wire N__42653;
    wire N__42650;
    wire N__42647;
    wire N__42644;
    wire N__42641;
    wire N__42640;
    wire N__42637;
    wire N__42636;
    wire N__42633;
    wire N__42630;
    wire N__42627;
    wire N__42626;
    wire N__42619;
    wire N__42616;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42604;
    wire N__42601;
    wire N__42596;
    wire N__42595;
    wire N__42592;
    wire N__42589;
    wire N__42588;
    wire N__42581;
    wire N__42580;
    wire N__42577;
    wire N__42576;
    wire N__42575;
    wire N__42574;
    wire N__42571;
    wire N__42570;
    wire N__42569;
    wire N__42568;
    wire N__42567;
    wire N__42566;
    wire N__42563;
    wire N__42560;
    wire N__42559;
    wire N__42558;
    wire N__42557;
    wire N__42556;
    wire N__42553;
    wire N__42552;
    wire N__42551;
    wire N__42550;
    wire N__42549;
    wire N__42546;
    wire N__42545;
    wire N__42538;
    wire N__42533;
    wire N__42530;
    wire N__42529;
    wire N__42528;
    wire N__42527;
    wire N__42526;
    wire N__42525;
    wire N__42524;
    wire N__42523;
    wire N__42522;
    wire N__42521;
    wire N__42516;
    wire N__42515;
    wire N__42514;
    wire N__42513;
    wire N__42512;
    wire N__42511;
    wire N__42510;
    wire N__42507;
    wire N__42500;
    wire N__42493;
    wire N__42490;
    wire N__42483;
    wire N__42478;
    wire N__42475;
    wire N__42470;
    wire N__42465;
    wire N__42462;
    wire N__42455;
    wire N__42452;
    wire N__42449;
    wire N__42446;
    wire N__42441;
    wire N__42434;
    wire N__42433;
    wire N__42432;
    wire N__42431;
    wire N__42430;
    wire N__42429;
    wire N__42428;
    wire N__42427;
    wire N__42426;
    wire N__42425;
    wire N__42424;
    wire N__42423;
    wire N__42422;
    wire N__42421;
    wire N__42418;
    wire N__42415;
    wire N__42412;
    wire N__42411;
    wire N__42408;
    wire N__42403;
    wire N__42400;
    wire N__42395;
    wire N__42388;
    wire N__42379;
    wire N__42376;
    wire N__42373;
    wire N__42370;
    wire N__42367;
    wire N__42360;
    wire N__42357;
    wire N__42352;
    wire N__42347;
    wire N__42344;
    wire N__42337;
    wire N__42334;
    wire N__42325;
    wire N__42320;
    wire N__42293;
    wire N__42290;
    wire N__42287;
    wire N__42284;
    wire N__42281;
    wire N__42278;
    wire N__42275;
    wire N__42272;
    wire N__42269;
    wire N__42266;
    wire N__42265;
    wire N__42264;
    wire N__42263;
    wire N__42260;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42249;
    wire N__42248;
    wire N__42247;
    wire N__42246;
    wire N__42245;
    wire N__42244;
    wire N__42243;
    wire N__42242;
    wire N__42241;
    wire N__42240;
    wire N__42239;
    wire N__42238;
    wire N__42235;
    wire N__42234;
    wire N__42233;
    wire N__42232;
    wire N__42231;
    wire N__42230;
    wire N__42229;
    wire N__42222;
    wire N__42219;
    wire N__42218;
    wire N__42215;
    wire N__42214;
    wire N__42213;
    wire N__42212;
    wire N__42211;
    wire N__42210;
    wire N__42209;
    wire N__42206;
    wire N__42205;
    wire N__42204;
    wire N__42203;
    wire N__42202;
    wire N__42199;
    wire N__42198;
    wire N__42197;
    wire N__42194;
    wire N__42193;
    wire N__42192;
    wire N__42191;
    wire N__42190;
    wire N__42189;
    wire N__42188;
    wire N__42185;
    wire N__42182;
    wire N__42181;
    wire N__42176;
    wire N__42175;
    wire N__42174;
    wire N__42173;
    wire N__42172;
    wire N__42171;
    wire N__42170;
    wire N__42169;
    wire N__42168;
    wire N__42167;
    wire N__42166;
    wire N__42165;
    wire N__42162;
    wire N__42161;
    wire N__42158;
    wire N__42157;
    wire N__42154;
    wire N__42153;
    wire N__42150;
    wire N__42149;
    wire N__42148;
    wire N__42147;
    wire N__42146;
    wire N__42145;
    wire N__42144;
    wire N__42143;
    wire N__42142;
    wire N__42139;
    wire N__42132;
    wire N__42125;
    wire N__42120;
    wire N__42115;
    wire N__42114;
    wire N__42113;
    wire N__42112;
    wire N__42111;
    wire N__42110;
    wire N__42109;
    wire N__42106;
    wire N__42105;
    wire N__42104;
    wire N__42101;
    wire N__42098;
    wire N__42097;
    wire N__42096;
    wire N__42095;
    wire N__42094;
    wire N__42093;
    wire N__42090;
    wire N__42083;
    wire N__42082;
    wire N__42081;
    wire N__42080;
    wire N__42077;
    wire N__42076;
    wire N__42075;
    wire N__42074;
    wire N__42073;
    wire N__42072;
    wire N__42069;
    wire N__42068;
    wire N__42067;
    wire N__42064;
    wire N__42053;
    wire N__42052;
    wire N__42049;
    wire N__42046;
    wire N__42039;
    wire N__42038;
    wire N__42037;
    wire N__42036;
    wire N__42035;
    wire N__42034;
    wire N__42033;
    wire N__42032;
    wire N__42029;
    wire N__42022;
    wire N__42019;
    wire N__42018;
    wire N__42017;
    wire N__42016;
    wire N__42015;
    wire N__42014;
    wire N__42013;
    wire N__42012;
    wire N__42011;
    wire N__42010;
    wire N__42007;
    wire N__42006;
    wire N__42003;
    wire N__42002;
    wire N__42001;
    wire N__42000;
    wire N__41997;
    wire N__41994;
    wire N__41991;
    wire N__41990;
    wire N__41989;
    wire N__41988;
    wire N__41987;
    wire N__41986;
    wire N__41985;
    wire N__41984;
    wire N__41983;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41975;
    wire N__41972;
    wire N__41965;
    wire N__41958;
    wire N__41953;
    wire N__41944;
    wire N__41937;
    wire N__41932;
    wire N__41929;
    wire N__41918;
    wire N__41911;
    wire N__41898;
    wire N__41893;
    wire N__41892;
    wire N__41891;
    wire N__41888;
    wire N__41887;
    wire N__41886;
    wire N__41885;
    wire N__41884;
    wire N__41879;
    wire N__41876;
    wire N__41875;
    wire N__41874;
    wire N__41873;
    wire N__41872;
    wire N__41869;
    wire N__41868;
    wire N__41867;
    wire N__41866;
    wire N__41865;
    wire N__41864;
    wire N__41863;
    wire N__41862;
    wire N__41861;
    wire N__41856;
    wire N__41851;
    wire N__41842;
    wire N__41841;
    wire N__41838;
    wire N__41831;
    wire N__41824;
    wire N__41821;
    wire N__41814;
    wire N__41813;
    wire N__41812;
    wire N__41811;
    wire N__41810;
    wire N__41809;
    wire N__41808;
    wire N__41807;
    wire N__41806;
    wire N__41805;
    wire N__41804;
    wire N__41801;
    wire N__41792;
    wire N__41785;
    wire N__41780;
    wire N__41777;
    wire N__41768;
    wire N__41763;
    wire N__41756;
    wire N__41749;
    wire N__41744;
    wire N__41735;
    wire N__41730;
    wire N__41723;
    wire N__41722;
    wire N__41721;
    wire N__41720;
    wire N__41717;
    wire N__41712;
    wire N__41709;
    wire N__41702;
    wire N__41689;
    wire N__41684;
    wire N__41675;
    wire N__41666;
    wire N__41659;
    wire N__41658;
    wire N__41657;
    wire N__41652;
    wire N__41643;
    wire N__41640;
    wire N__41631;
    wire N__41622;
    wire N__41615;
    wire N__41610;
    wire N__41609;
    wire N__41608;
    wire N__41607;
    wire N__41606;
    wire N__41605;
    wire N__41596;
    wire N__41587;
    wire N__41582;
    wire N__41579;
    wire N__41572;
    wire N__41567;
    wire N__41566;
    wire N__41565;
    wire N__41564;
    wire N__41563;
    wire N__41560;
    wire N__41557;
    wire N__41548;
    wire N__41541;
    wire N__41538;
    wire N__41537;
    wire N__41536;
    wire N__41533;
    wire N__41526;
    wire N__41523;
    wire N__41506;
    wire N__41501;
    wire N__41494;
    wire N__41489;
    wire N__41484;
    wire N__41479;
    wire N__41476;
    wire N__41471;
    wire N__41464;
    wire N__41457;
    wire N__41448;
    wire N__41441;
    wire N__41436;
    wire N__41431;
    wire N__41424;
    wire N__41419;
    wire N__41412;
    wire N__41387;
    wire N__41384;
    wire N__41381;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41369;
    wire N__41366;
    wire N__41363;
    wire N__41360;
    wire N__41357;
    wire N__41354;
    wire N__41351;
    wire N__41348;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41303;
    wire N__41300;
    wire N__41297;
    wire N__41294;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41276;
    wire N__41275;
    wire N__41272;
    wire N__41269;
    wire N__41266;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41249;
    wire N__41246;
    wire N__41243;
    wire N__41240;
    wire N__41237;
    wire N__41234;
    wire N__41231;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41213;
    wire N__41210;
    wire N__41207;
    wire N__41204;
    wire N__41201;
    wire N__41198;
    wire N__41195;
    wire N__41192;
    wire N__41189;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41165;
    wire N__41162;
    wire N__41159;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41147;
    wire N__41144;
    wire N__41141;
    wire N__41138;
    wire N__41135;
    wire N__41132;
    wire N__41129;
    wire N__41126;
    wire N__41123;
    wire N__41120;
    wire N__41117;
    wire N__41114;
    wire N__41111;
    wire N__41108;
    wire N__41105;
    wire N__41102;
    wire N__41099;
    wire N__41096;
    wire N__41093;
    wire N__41090;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41078;
    wire N__41075;
    wire N__41072;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41060;
    wire N__41057;
    wire N__41054;
    wire N__41051;
    wire N__41048;
    wire N__41045;
    wire N__41042;
    wire N__41039;
    wire N__41036;
    wire N__41033;
    wire N__41030;
    wire N__41027;
    wire N__41026;
    wire N__41023;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41011;
    wire N__41010;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__41000;
    wire N__40999;
    wire N__40998;
    wire N__40997;
    wire N__40996;
    wire N__40995;
    wire N__40994;
    wire N__40991;
    wire N__40986;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40978;
    wire N__40977;
    wire N__40976;
    wire N__40973;
    wire N__40970;
    wire N__40969;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40961;
    wire N__40960;
    wire N__40957;
    wire N__40956;
    wire N__40951;
    wire N__40950;
    wire N__40949;
    wire N__40940;
    wire N__40937;
    wire N__40934;
    wire N__40931;
    wire N__40922;
    wire N__40915;
    wire N__40910;
    wire N__40907;
    wire N__40904;
    wire N__40901;
    wire N__40900;
    wire N__40897;
    wire N__40896;
    wire N__40895;
    wire N__40894;
    wire N__40889;
    wire N__40882;
    wire N__40877;
    wire N__40872;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40864;
    wire N__40863;
    wire N__40862;
    wire N__40861;
    wire N__40854;
    wire N__40851;
    wire N__40844;
    wire N__40839;
    wire N__40836;
    wire N__40829;
    wire N__40826;
    wire N__40811;
    wire N__40810;
    wire N__40809;
    wire N__40806;
    wire N__40801;
    wire N__40800;
    wire N__40799;
    wire N__40798;
    wire N__40797;
    wire N__40796;
    wire N__40795;
    wire N__40794;
    wire N__40793;
    wire N__40790;
    wire N__40787;
    wire N__40786;
    wire N__40785;
    wire N__40784;
    wire N__40775;
    wire N__40766;
    wire N__40761;
    wire N__40754;
    wire N__40753;
    wire N__40752;
    wire N__40751;
    wire N__40748;
    wire N__40747;
    wire N__40746;
    wire N__40745;
    wire N__40744;
    wire N__40743;
    wire N__40742;
    wire N__40741;
    wire N__40740;
    wire N__40733;
    wire N__40726;
    wire N__40723;
    wire N__40720;
    wire N__40715;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40676;
    wire N__40675;
    wire N__40674;
    wire N__40673;
    wire N__40670;
    wire N__40669;
    wire N__40660;
    wire N__40659;
    wire N__40658;
    wire N__40655;
    wire N__40654;
    wire N__40653;
    wire N__40652;
    wire N__40651;
    wire N__40648;
    wire N__40647;
    wire N__40646;
    wire N__40645;
    wire N__40642;
    wire N__40633;
    wire N__40632;
    wire N__40627;
    wire N__40624;
    wire N__40621;
    wire N__40620;
    wire N__40619;
    wire N__40618;
    wire N__40617;
    wire N__40616;
    wire N__40615;
    wire N__40610;
    wire N__40605;
    wire N__40604;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40592;
    wire N__40589;
    wire N__40580;
    wire N__40577;
    wire N__40572;
    wire N__40567;
    wire N__40562;
    wire N__40547;
    wire N__40546;
    wire N__40545;
    wire N__40540;
    wire N__40537;
    wire N__40534;
    wire N__40533;
    wire N__40532;
    wire N__40531;
    wire N__40528;
    wire N__40525;
    wire N__40522;
    wire N__40521;
    wire N__40520;
    wire N__40517;
    wire N__40516;
    wire N__40513;
    wire N__40510;
    wire N__40509;
    wire N__40508;
    wire N__40507;
    wire N__40504;
    wire N__40501;
    wire N__40500;
    wire N__40497;
    wire N__40496;
    wire N__40493;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40479;
    wire N__40474;
    wire N__40469;
    wire N__40466;
    wire N__40461;
    wire N__40456;
    wire N__40439;
    wire N__40438;
    wire N__40437;
    wire N__40434;
    wire N__40433;
    wire N__40430;
    wire N__40429;
    wire N__40428;
    wire N__40419;
    wire N__40418;
    wire N__40417;
    wire N__40416;
    wire N__40413;
    wire N__40412;
    wire N__40411;
    wire N__40410;
    wire N__40409;
    wire N__40408;
    wire N__40407;
    wire N__40406;
    wire N__40405;
    wire N__40404;
    wire N__40403;
    wire N__40402;
    wire N__40399;
    wire N__40396;
    wire N__40391;
    wire N__40386;
    wire N__40385;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40377;
    wire N__40374;
    wire N__40367;
    wire N__40364;
    wire N__40357;
    wire N__40354;
    wire N__40351;
    wire N__40348;
    wire N__40343;
    wire N__40340;
    wire N__40337;
    wire N__40336;
    wire N__40335;
    wire N__40334;
    wire N__40329;
    wire N__40326;
    wire N__40315;
    wire N__40308;
    wire N__40307;
    wire N__40306;
    wire N__40305;
    wire N__40304;
    wire N__40303;
    wire N__40302;
    wire N__40301;
    wire N__40300;
    wire N__40299;
    wire N__40298;
    wire N__40297;
    wire N__40296;
    wire N__40295;
    wire N__40294;
    wire N__40289;
    wire N__40286;
    wire N__40281;
    wire N__40278;
    wire N__40275;
    wire N__40270;
    wire N__40269;
    wire N__40264;
    wire N__40255;
    wire N__40252;
    wire N__40241;
    wire N__40236;
    wire N__40233;
    wire N__40224;
    wire N__40221;
    wire N__40218;
    wire N__40199;
    wire N__40198;
    wire N__40197;
    wire N__40196;
    wire N__40195;
    wire N__40192;
    wire N__40191;
    wire N__40190;
    wire N__40189;
    wire N__40186;
    wire N__40181;
    wire N__40180;
    wire N__40177;
    wire N__40176;
    wire N__40175;
    wire N__40164;
    wire N__40163;
    wire N__40162;
    wire N__40161;
    wire N__40160;
    wire N__40159;
    wire N__40158;
    wire N__40157;
    wire N__40154;
    wire N__40151;
    wire N__40148;
    wire N__40143;
    wire N__40140;
    wire N__40139;
    wire N__40134;
    wire N__40129;
    wire N__40124;
    wire N__40121;
    wire N__40120;
    wire N__40117;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40097;
    wire N__40092;
    wire N__40089;
    wire N__40084;
    wire N__40073;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40054;
    wire N__40053;
    wire N__40052;
    wire N__40049;
    wire N__40046;
    wire N__40041;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40027;
    wire N__40026;
    wire N__40025;
    wire N__40024;
    wire N__40021;
    wire N__40016;
    wire N__40011;
    wire N__40010;
    wire N__40009;
    wire N__40006;
    wire N__40003;
    wire N__40002;
    wire N__39999;
    wire N__39998;
    wire N__39997;
    wire N__39992;
    wire N__39991;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39979;
    wire N__39974;
    wire N__39973;
    wire N__39972;
    wire N__39971;
    wire N__39970;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39958;
    wire N__39951;
    wire N__39948;
    wire N__39945;
    wire N__39940;
    wire N__39937;
    wire N__39920;
    wire N__39917;
    wire N__39914;
    wire N__39911;
    wire N__39908;
    wire N__39905;
    wire N__39902;
    wire N__39899;
    wire N__39896;
    wire N__39893;
    wire N__39890;
    wire N__39887;
    wire N__39884;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39866;
    wire N__39863;
    wire N__39860;
    wire N__39857;
    wire N__39854;
    wire N__39851;
    wire N__39848;
    wire N__39845;
    wire N__39842;
    wire N__39839;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39821;
    wire N__39818;
    wire N__39815;
    wire N__39812;
    wire N__39809;
    wire N__39806;
    wire N__39803;
    wire N__39802;
    wire N__39799;
    wire N__39796;
    wire N__39791;
    wire N__39788;
    wire N__39785;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39772;
    wire N__39769;
    wire N__39766;
    wire N__39763;
    wire N__39760;
    wire N__39755;
    wire N__39752;
    wire N__39749;
    wire N__39746;
    wire N__39743;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39725;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39713;
    wire N__39712;
    wire N__39709;
    wire N__39706;
    wire N__39701;
    wire N__39698;
    wire N__39695;
    wire N__39692;
    wire N__39689;
    wire N__39686;
    wire N__39683;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39671;
    wire N__39668;
    wire N__39665;
    wire N__39662;
    wire N__39659;
    wire N__39656;
    wire N__39653;
    wire N__39650;
    wire N__39647;
    wire N__39644;
    wire N__39641;
    wire N__39638;
    wire N__39635;
    wire N__39632;
    wire N__39629;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39608;
    wire N__39605;
    wire N__39602;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39592;
    wire N__39587;
    wire N__39584;
    wire N__39583;
    wire N__39580;
    wire N__39577;
    wire N__39574;
    wire N__39569;
    wire N__39566;
    wire N__39565;
    wire N__39562;
    wire N__39559;
    wire N__39556;
    wire N__39551;
    wire N__39548;
    wire N__39547;
    wire N__39544;
    wire N__39541;
    wire N__39538;
    wire N__39533;
    wire N__39530;
    wire N__39529;
    wire N__39526;
    wire N__39523;
    wire N__39520;
    wire N__39515;
    wire N__39512;
    wire N__39511;
    wire N__39510;
    wire N__39509;
    wire N__39508;
    wire N__39507;
    wire N__39506;
    wire N__39505;
    wire N__39496;
    wire N__39487;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39475;
    wire N__39472;
    wire N__39469;
    wire N__39466;
    wire N__39461;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39445;
    wire N__39442;
    wire N__39439;
    wire N__39436;
    wire N__39433;
    wire N__39428;
    wire N__39425;
    wire N__39422;
    wire N__39421;
    wire N__39418;
    wire N__39415;
    wire N__39410;
    wire N__39409;
    wire N__39408;
    wire N__39407;
    wire N__39406;
    wire N__39405;
    wire N__39404;
    wire N__39403;
    wire N__39402;
    wire N__39401;
    wire N__39400;
    wire N__39399;
    wire N__39398;
    wire N__39397;
    wire N__39396;
    wire N__39395;
    wire N__39394;
    wire N__39393;
    wire N__39392;
    wire N__39391;
    wire N__39390;
    wire N__39389;
    wire N__39388;
    wire N__39387;
    wire N__39378;
    wire N__39369;
    wire N__39360;
    wire N__39359;
    wire N__39358;
    wire N__39357;
    wire N__39356;
    wire N__39351;
    wire N__39348;
    wire N__39347;
    wire N__39346;
    wire N__39345;
    wire N__39344;
    wire N__39343;
    wire N__39342;
    wire N__39341;
    wire N__39340;
    wire N__39331;
    wire N__39322;
    wire N__39319;
    wire N__39312;
    wire N__39303;
    wire N__39298;
    wire N__39297;
    wire N__39296;
    wire N__39295;
    wire N__39286;
    wire N__39277;
    wire N__39272;
    wire N__39269;
    wire N__39262;
    wire N__39257;
    wire N__39254;
    wire N__39249;
    wire N__39248;
    wire N__39243;
    wire N__39240;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39226;
    wire N__39225;
    wire N__39220;
    wire N__39215;
    wire N__39212;
    wire N__39209;
    wire N__39204;
    wire N__39201;
    wire N__39194;
    wire N__39191;
    wire N__39188;
    wire N__39185;
    wire N__39182;
    wire N__39179;
    wire N__39176;
    wire N__39173;
    wire N__39172;
    wire N__39169;
    wire N__39166;
    wire N__39165;
    wire N__39164;
    wire N__39163;
    wire N__39160;
    wire N__39155;
    wire N__39150;
    wire N__39145;
    wire N__39140;
    wire N__39139;
    wire N__39134;
    wire N__39131;
    wire N__39130;
    wire N__39129;
    wire N__39128;
    wire N__39127;
    wire N__39124;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39104;
    wire N__39101;
    wire N__39098;
    wire N__39095;
    wire N__39092;
    wire N__39089;
    wire N__39086;
    wire N__39083;
    wire N__39082;
    wire N__39079;
    wire N__39076;
    wire N__39071;
    wire N__39068;
    wire N__39065;
    wire N__39062;
    wire N__39059;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39047;
    wire N__39046;
    wire N__39043;
    wire N__39040;
    wire N__39037;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39025;
    wire N__39022;
    wire N__39019;
    wire N__39016;
    wire N__39011;
    wire N__39008;
    wire N__39005;
    wire N__39002;
    wire N__38999;
    wire N__38996;
    wire N__38993;
    wire N__38990;
    wire N__38987;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38975;
    wire N__38972;
    wire N__38969;
    wire N__38966;
    wire N__38963;
    wire N__38960;
    wire N__38957;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38942;
    wire N__38939;
    wire N__38936;
    wire N__38933;
    wire N__38930;
    wire N__38927;
    wire N__38924;
    wire N__38921;
    wire N__38918;
    wire N__38915;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38905;
    wire N__38902;
    wire N__38899;
    wire N__38896;
    wire N__38891;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38881;
    wire N__38876;
    wire N__38873;
    wire N__38872;
    wire N__38869;
    wire N__38866;
    wire N__38863;
    wire N__38858;
    wire N__38857;
    wire N__38854;
    wire N__38851;
    wire N__38848;
    wire N__38843;
    wire N__38840;
    wire N__38837;
    wire N__38834;
    wire N__38831;
    wire N__38830;
    wire N__38827;
    wire N__38824;
    wire N__38821;
    wire N__38816;
    wire N__38815;
    wire N__38812;
    wire N__38809;
    wire N__38806;
    wire N__38801;
    wire N__38798;
    wire N__38795;
    wire N__38794;
    wire N__38791;
    wire N__38788;
    wire N__38785;
    wire N__38780;
    wire N__38779;
    wire N__38776;
    wire N__38773;
    wire N__38770;
    wire N__38765;
    wire N__38762;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38735;
    wire N__38732;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38717;
    wire N__38714;
    wire N__38711;
    wire N__38708;
    wire N__38705;
    wire N__38702;
    wire N__38699;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38672;
    wire N__38669;
    wire N__38666;
    wire N__38663;
    wire N__38660;
    wire N__38657;
    wire N__38654;
    wire N__38653;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38639;
    wire N__38636;
    wire N__38633;
    wire N__38630;
    wire N__38627;
    wire N__38624;
    wire N__38621;
    wire N__38618;
    wire N__38615;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38591;
    wire N__38588;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38576;
    wire N__38573;
    wire N__38570;
    wire N__38567;
    wire N__38564;
    wire N__38561;
    wire N__38558;
    wire N__38557;
    wire N__38556;
    wire N__38555;
    wire N__38554;
    wire N__38553;
    wire N__38552;
    wire N__38551;
    wire N__38550;
    wire N__38547;
    wire N__38542;
    wire N__38539;
    wire N__38534;
    wire N__38533;
    wire N__38532;
    wire N__38531;
    wire N__38530;
    wire N__38527;
    wire N__38526;
    wire N__38521;
    wire N__38512;
    wire N__38511;
    wire N__38510;
    wire N__38509;
    wire N__38508;
    wire N__38507;
    wire N__38506;
    wire N__38501;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38491;
    wire N__38490;
    wire N__38489;
    wire N__38486;
    wire N__38481;
    wire N__38478;
    wire N__38477;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38461;
    wire N__38460;
    wire N__38459;
    wire N__38456;
    wire N__38453;
    wire N__38452;
    wire N__38449;
    wire N__38448;
    wire N__38445;
    wire N__38442;
    wire N__38437;
    wire N__38430;
    wire N__38427;
    wire N__38426;
    wire N__38425;
    wire N__38420;
    wire N__38415;
    wire N__38414;
    wire N__38409;
    wire N__38404;
    wire N__38403;
    wire N__38402;
    wire N__38397;
    wire N__38394;
    wire N__38391;
    wire N__38388;
    wire N__38387;
    wire N__38384;
    wire N__38375;
    wire N__38372;
    wire N__38369;
    wire N__38364;
    wire N__38361;
    wire N__38356;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38340;
    wire N__38337;
    wire N__38332;
    wire N__38321;
    wire N__38306;
    wire N__38303;
    wire N__38302;
    wire N__38301;
    wire N__38300;
    wire N__38297;
    wire N__38292;
    wire N__38291;
    wire N__38290;
    wire N__38289;
    wire N__38288;
    wire N__38287;
    wire N__38286;
    wire N__38285;
    wire N__38282;
    wire N__38277;
    wire N__38272;
    wire N__38263;
    wire N__38262;
    wire N__38259;
    wire N__38258;
    wire N__38257;
    wire N__38256;
    wire N__38255;
    wire N__38254;
    wire N__38253;
    wire N__38252;
    wire N__38251;
    wire N__38250;
    wire N__38249;
    wire N__38246;
    wire N__38239;
    wire N__38234;
    wire N__38233;
    wire N__38232;
    wire N__38231;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38218;
    wire N__38217;
    wire N__38216;
    wire N__38213;
    wire N__38212;
    wire N__38211;
    wire N__38210;
    wire N__38209;
    wire N__38208;
    wire N__38207;
    wire N__38204;
    wire N__38203;
    wire N__38202;
    wire N__38201;
    wire N__38200;
    wire N__38197;
    wire N__38196;
    wire N__38195;
    wire N__38194;
    wire N__38191;
    wire N__38190;
    wire N__38185;
    wire N__38178;
    wire N__38177;
    wire N__38174;
    wire N__38171;
    wire N__38170;
    wire N__38169;
    wire N__38168;
    wire N__38167;
    wire N__38166;
    wire N__38163;
    wire N__38156;
    wire N__38151;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38135;
    wire N__38132;
    wire N__38131;
    wire N__38130;
    wire N__38129;
    wire N__38126;
    wire N__38123;
    wire N__38122;
    wire N__38121;
    wire N__38118;
    wire N__38117;
    wire N__38116;
    wire N__38115;
    wire N__38112;
    wire N__38111;
    wire N__38108;
    wire N__38105;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38097;
    wire N__38096;
    wire N__38095;
    wire N__38092;
    wire N__38091;
    wire N__38088;
    wire N__38083;
    wire N__38080;
    wire N__38075;
    wire N__38066;
    wire N__38061;
    wire N__38056;
    wire N__38053;
    wire N__38048;
    wire N__38045;
    wire N__38042;
    wire N__38035;
    wire N__38032;
    wire N__38031;
    wire N__38030;
    wire N__38025;
    wire N__38020;
    wire N__38015;
    wire N__38012;
    wire N__38009;
    wire N__38002;
    wire N__38001;
    wire N__37998;
    wire N__37997;
    wire N__37994;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37975;
    wire N__37968;
    wire N__37959;
    wire N__37948;
    wire N__37943;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37929;
    wire N__37926;
    wire N__37919;
    wire N__37916;
    wire N__37913;
    wire N__37910;
    wire N__37907;
    wire N__37902;
    wire N__37891;
    wire N__37886;
    wire N__37873;
    wire N__37856;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37838;
    wire N__37835;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37808;
    wire N__37807;
    wire N__37806;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37796;
    wire N__37793;
    wire N__37790;
    wire N__37789;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37765;
    wire N__37760;
    wire N__37755;
    wire N__37752;
    wire N__37749;
    wire N__37746;
    wire N__37739;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37727;
    wire N__37724;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37706;
    wire N__37703;
    wire N__37700;
    wire N__37697;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37676;
    wire N__37673;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37655;
    wire N__37652;
    wire N__37649;
    wire N__37646;
    wire N__37643;
    wire N__37640;
    wire N__37637;
    wire N__37636;
    wire N__37635;
    wire N__37634;
    wire N__37633;
    wire N__37632;
    wire N__37631;
    wire N__37630;
    wire N__37629;
    wire N__37628;
    wire N__37627;
    wire N__37624;
    wire N__37621;
    wire N__37618;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37593;
    wire N__37590;
    wire N__37585;
    wire N__37584;
    wire N__37583;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37564;
    wire N__37561;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37539;
    wire N__37526;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37505;
    wire N__37502;
    wire N__37499;
    wire N__37496;
    wire N__37493;
    wire N__37490;
    wire N__37487;
    wire N__37486;
    wire N__37485;
    wire N__37482;
    wire N__37481;
    wire N__37478;
    wire N__37473;
    wire N__37472;
    wire N__37471;
    wire N__37468;
    wire N__37463;
    wire N__37462;
    wire N__37461;
    wire N__37458;
    wire N__37457;
    wire N__37456;
    wire N__37455;
    wire N__37454;
    wire N__37449;
    wire N__37446;
    wire N__37443;
    wire N__37442;
    wire N__37441;
    wire N__37440;
    wire N__37439;
    wire N__37436;
    wire N__37433;
    wire N__37428;
    wire N__37423;
    wire N__37420;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37408;
    wire N__37403;
    wire N__37396;
    wire N__37391;
    wire N__37390;
    wire N__37387;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37371;
    wire N__37368;
    wire N__37355;
    wire N__37352;
    wire N__37351;
    wire N__37348;
    wire N__37345;
    wire N__37344;
    wire N__37343;
    wire N__37342;
    wire N__37341;
    wire N__37336;
    wire N__37335;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37327;
    wire N__37324;
    wire N__37321;
    wire N__37318;
    wire N__37315;
    wire N__37312;
    wire N__37309;
    wire N__37306;
    wire N__37305;
    wire N__37302;
    wire N__37297;
    wire N__37290;
    wire N__37285;
    wire N__37282;
    wire N__37271;
    wire N__37268;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37232;
    wire N__37229;
    wire N__37226;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36964;
    wire N__36961;
    wire N__36960;
    wire N__36959;
    wire N__36956;
    wire N__36953;
    wire N__36952;
    wire N__36949;
    wire N__36946;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36924;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36910;
    wire N__36907;
    wire N__36902;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36875;
    wire N__36872;
    wire N__36869;
    wire N__36866;
    wire N__36863;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36851;
    wire N__36848;
    wire N__36845;
    wire N__36842;
    wire N__36839;
    wire N__36836;
    wire N__36833;
    wire N__36830;
    wire N__36827;
    wire N__36824;
    wire N__36821;
    wire N__36818;
    wire N__36815;
    wire N__36812;
    wire N__36809;
    wire N__36806;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36662;
    wire N__36659;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36637;
    wire N__36634;
    wire N__36631;
    wire N__36628;
    wire N__36625;
    wire N__36622;
    wire N__36619;
    wire N__36616;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36587;
    wire N__36584;
    wire N__36581;
    wire N__36578;
    wire N__36575;
    wire N__36572;
    wire N__36569;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36553;
    wire N__36550;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36540;
    wire N__36537;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36523;
    wire N__36520;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36488;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36449;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36428;
    wire N__36425;
    wire N__36422;
    wire N__36419;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36395;
    wire N__36392;
    wire N__36389;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36367;
    wire N__36364;
    wire N__36361;
    wire N__36356;
    wire N__36353;
    wire N__36350;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36323;
    wire N__36322;
    wire N__36319;
    wire N__36316;
    wire N__36311;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36290;
    wire N__36287;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36275;
    wire N__36272;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36260;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36239;
    wire N__36236;
    wire N__36233;
    wire N__36230;
    wire N__36229;
    wire N__36226;
    wire N__36223;
    wire N__36218;
    wire N__36215;
    wire N__36212;
    wire N__36209;
    wire N__36206;
    wire N__36203;
    wire N__36200;
    wire N__36197;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36182;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36163;
    wire N__36160;
    wire N__36157;
    wire N__36152;
    wire N__36149;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36131;
    wire N__36130;
    wire N__36127;
    wire N__36124;
    wire N__36119;
    wire N__36116;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36101;
    wire N__36100;
    wire N__36097;
    wire N__36094;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36058;
    wire N__36055;
    wire N__36052;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36040;
    wire N__36037;
    wire N__36034;
    wire N__36029;
    wire N__36026;
    wire N__36023;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36008;
    wire N__36005;
    wire N__36002;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35990;
    wire N__35987;
    wire N__35984;
    wire N__35983;
    wire N__35980;
    wire N__35977;
    wire N__35972;
    wire N__35969;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35945;
    wire N__35942;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35918;
    wire N__35915;
    wire N__35912;
    wire N__35909;
    wire N__35906;
    wire N__35903;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35891;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35879;
    wire N__35876;
    wire N__35873;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35839;
    wire N__35836;
    wire N__35833;
    wire N__35828;
    wire N__35825;
    wire N__35822;
    wire N__35819;
    wire N__35816;
    wire N__35813;
    wire N__35810;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35798;
    wire N__35795;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35777;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35767;
    wire N__35764;
    wire N__35761;
    wire N__35756;
    wire N__35753;
    wire N__35750;
    wire N__35747;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35737;
    wire N__35734;
    wire N__35731;
    wire N__35726;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35693;
    wire N__35690;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35671;
    wire N__35668;
    wire N__35665;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35645;
    wire N__35642;
    wire N__35639;
    wire N__35636;
    wire N__35633;
    wire N__35632;
    wire N__35629;
    wire N__35626;
    wire N__35621;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35606;
    wire N__35605;
    wire N__35602;
    wire N__35599;
    wire N__35594;
    wire N__35591;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35560;
    wire N__35557;
    wire N__35554;
    wire N__35549;
    wire N__35546;
    wire N__35543;
    wire N__35540;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35528;
    wire N__35525;
    wire N__35522;
    wire N__35519;
    wire N__35516;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35498;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35453;
    wire N__35450;
    wire N__35447;
    wire N__35444;
    wire N__35441;
    wire N__35438;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35425;
    wire N__35422;
    wire N__35419;
    wire N__35414;
    wire N__35411;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35399;
    wire N__35396;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35381;
    wire N__35378;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35359;
    wire N__35356;
    wire N__35353;
    wire N__35348;
    wire N__35345;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35333;
    wire N__35330;
    wire N__35329;
    wire N__35326;
    wire N__35323;
    wire N__35320;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35305;
    wire N__35302;
    wire N__35299;
    wire N__35296;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35284;
    wire N__35281;
    wire N__35278;
    wire N__35275;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35249;
    wire N__35248;
    wire N__35245;
    wire N__35242;
    wire N__35237;
    wire N__35234;
    wire N__35231;
    wire N__35228;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35216;
    wire N__35213;
    wire N__35210;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35180;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35165;
    wire N__35162;
    wire N__35159;
    wire N__35158;
    wire N__35155;
    wire N__35152;
    wire N__35149;
    wire N__35144;
    wire N__35141;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35126;
    wire N__35123;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35111;
    wire N__35108;
    wire N__35105;
    wire N__35102;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35090;
    wire N__35087;
    wire N__35086;
    wire N__35083;
    wire N__35080;
    wire N__35075;
    wire N__35072;
    wire N__35071;
    wire N__35068;
    wire N__35065;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35024;
    wire N__35021;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35006;
    wire N__35003;
    wire N__35000;
    wire N__34997;
    wire N__34994;
    wire N__34991;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34979;
    wire N__34976;
    wire N__34973;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34961;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34946;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34934;
    wire N__34931;
    wire N__34928;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34913;
    wire N__34910;
    wire N__34907;
    wire N__34904;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34880;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34867;
    wire N__34866;
    wire N__34863;
    wire N__34860;
    wire N__34859;
    wire N__34858;
    wire N__34857;
    wire N__34854;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34836;
    wire N__34829;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34805;
    wire N__34802;
    wire N__34799;
    wire N__34796;
    wire N__34793;
    wire N__34790;
    wire N__34787;
    wire N__34784;
    wire N__34781;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34763;
    wire N__34760;
    wire N__34757;
    wire N__34754;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34694;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34631;
    wire N__34628;
    wire N__34625;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34613;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34598;
    wire N__34595;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34580;
    wire N__34577;
    wire N__34574;
    wire N__34571;
    wire N__34568;
    wire N__34565;
    wire N__34562;
    wire N__34559;
    wire N__34556;
    wire N__34553;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34532;
    wire N__34529;
    wire N__34526;
    wire N__34523;
    wire N__34520;
    wire N__34517;
    wire N__34514;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34481;
    wire N__34478;
    wire N__34475;
    wire N__34472;
    wire N__34469;
    wire N__34466;
    wire N__34463;
    wire N__34460;
    wire N__34457;
    wire N__34454;
    wire N__34451;
    wire N__34448;
    wire N__34445;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34427;
    wire N__34424;
    wire N__34421;
    wire N__34418;
    wire N__34415;
    wire N__34412;
    wire N__34409;
    wire N__34406;
    wire N__34403;
    wire N__34400;
    wire N__34397;
    wire N__34394;
    wire N__34391;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34367;
    wire N__34364;
    wire N__34361;
    wire N__34358;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34331;
    wire N__34328;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34316;
    wire N__34313;
    wire N__34310;
    wire N__34307;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34292;
    wire N__34289;
    wire N__34286;
    wire N__34283;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34271;
    wire N__34268;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34250;
    wire N__34247;
    wire N__34244;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34217;
    wire N__34214;
    wire N__34211;
    wire N__34208;
    wire N__34205;
    wire N__34202;
    wire N__34199;
    wire N__34196;
    wire N__34193;
    wire N__34190;
    wire N__34187;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34175;
    wire N__34172;
    wire N__34169;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34145;
    wire N__34142;
    wire N__34139;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34127;
    wire N__34124;
    wire N__34121;
    wire N__34118;
    wire N__34115;
    wire N__34112;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34100;
    wire N__34097;
    wire N__34094;
    wire N__34091;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34058;
    wire N__34055;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34028;
    wire N__34025;
    wire N__34022;
    wire N__34019;
    wire N__34016;
    wire N__34015;
    wire N__34014;
    wire N__34013;
    wire N__34010;
    wire N__34007;
    wire N__34006;
    wire N__34001;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33983;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33887;
    wire N__33884;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33839;
    wire N__33836;
    wire N__33833;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33769;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33755;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33747;
    wire N__33746;
    wire N__33745;
    wire N__33744;
    wire N__33743;
    wire N__33740;
    wire N__33739;
    wire N__33734;
    wire N__33733;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33723;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33698;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33560;
    wire N__33557;
    wire N__33554;
    wire N__33551;
    wire N__33548;
    wire N__33545;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33512;
    wire N__33509;
    wire N__33508;
    wire N__33505;
    wire N__33504;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33487;
    wire N__33484;
    wire N__33481;
    wire N__33478;
    wire N__33475;
    wire N__33470;
    wire N__33467;
    wire N__33464;
    wire N__33461;
    wire N__33458;
    wire N__33455;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33434;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33392;
    wire N__33389;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33381;
    wire N__33380;
    wire N__33377;
    wire N__33376;
    wire N__33375;
    wire N__33374;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33366;
    wire N__33363;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33339;
    wire N__33336;
    wire N__33333;
    wire N__33332;
    wire N__33331;
    wire N__33326;
    wire N__33321;
    wire N__33318;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33294;
    wire N__33287;
    wire N__33278;
    wire N__33277;
    wire N__33276;
    wire N__33275;
    wire N__33274;
    wire N__33273;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33257;
    wire N__33254;
    wire N__33253;
    wire N__33250;
    wire N__33249;
    wire N__33246;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33225;
    wire N__33224;
    wire N__33223;
    wire N__33220;
    wire N__33215;
    wire N__33210;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33181;
    wire N__33170;
    wire N__33169;
    wire N__33168;
    wire N__33167;
    wire N__33166;
    wire N__33165;
    wire N__33162;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33154;
    wire N__33151;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33129;
    wire N__33126;
    wire N__33123;
    wire N__33120;
    wire N__33117;
    wire N__33116;
    wire N__33115;
    wire N__33110;
    wire N__33105;
    wire N__33102;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33078;
    wire N__33071;
    wire N__33062;
    wire N__33059;
    wire N__33058;
    wire N__33057;
    wire N__33054;
    wire N__33053;
    wire N__33052;
    wire N__33049;
    wire N__33048;
    wire N__33047;
    wire N__33046;
    wire N__33043;
    wire N__33040;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32990;
    wire N__32987;
    wire N__32976;
    wire N__32973;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32942;
    wire N__32939;
    wire N__32936;
    wire N__32933;
    wire N__32930;
    wire N__32927;
    wire N__32924;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32903;
    wire N__32900;
    wire N__32897;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32864;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32851;
    wire N__32848;
    wire N__32845;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32828;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32816;
    wire N__32813;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32792;
    wire N__32789;
    wire N__32786;
    wire N__32783;
    wire N__32780;
    wire N__32777;
    wire N__32774;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32660;
    wire N__32657;
    wire N__32654;
    wire N__32651;
    wire N__32648;
    wire N__32645;
    wire N__32642;
    wire N__32639;
    wire N__32636;
    wire N__32633;
    wire N__32630;
    wire N__32627;
    wire N__32624;
    wire N__32621;
    wire N__32618;
    wire N__32615;
    wire N__32612;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32597;
    wire N__32594;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32570;
    wire N__32567;
    wire N__32564;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32543;
    wire N__32540;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32522;
    wire N__32519;
    wire N__32516;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32498;
    wire N__32495;
    wire N__32492;
    wire N__32489;
    wire N__32486;
    wire N__32483;
    wire N__32480;
    wire N__32477;
    wire N__32474;
    wire N__32471;
    wire N__32468;
    wire N__32465;
    wire N__32462;
    wire N__32459;
    wire N__32456;
    wire N__32453;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32420;
    wire N__32417;
    wire N__32414;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32399;
    wire N__32396;
    wire N__32393;
    wire N__32390;
    wire N__32387;
    wire N__32384;
    wire N__32381;
    wire N__32378;
    wire N__32375;
    wire N__32372;
    wire N__32369;
    wire N__32366;
    wire N__32363;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32351;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32333;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32321;
    wire N__32318;
    wire N__32315;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32288;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32216;
    wire N__32213;
    wire N__32210;
    wire N__32207;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32090;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32060;
    wire N__32057;
    wire N__32054;
    wire N__32051;
    wire N__32048;
    wire N__32047;
    wire N__32046;
    wire N__32045;
    wire N__32042;
    wire N__32041;
    wire N__32038;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32027;
    wire N__32024;
    wire N__32021;
    wire N__32020;
    wire N__32019;
    wire N__32018;
    wire N__32015;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31991;
    wire N__31990;
    wire N__31987;
    wire N__31984;
    wire N__31981;
    wire N__31976;
    wire N__31973;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31951;
    wire N__31946;
    wire N__31937;
    wire N__31936;
    wire N__31935;
    wire N__31934;
    wire N__31931;
    wire N__31930;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31913;
    wire N__31910;
    wire N__31909;
    wire N__31906;
    wire N__31905;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31883;
    wire N__31882;
    wire N__31879;
    wire N__31876;
    wire N__31873;
    wire N__31866;
    wire N__31863;
    wire N__31858;
    wire N__31855;
    wire N__31852;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31838;
    wire N__31835;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31805;
    wire N__31802;
    wire N__31799;
    wire N__31796;
    wire N__31793;
    wire N__31790;
    wire N__31787;
    wire N__31784;
    wire N__31781;
    wire N__31778;
    wire N__31775;
    wire N__31772;
    wire N__31769;
    wire N__31766;
    wire N__31763;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31748;
    wire N__31747;
    wire N__31744;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31733;
    wire N__31732;
    wire N__31729;
    wire N__31726;
    wire N__31723;
    wire N__31722;
    wire N__31719;
    wire N__31718;
    wire N__31717;
    wire N__31714;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31700;
    wire N__31697;
    wire N__31694;
    wire N__31691;
    wire N__31688;
    wire N__31685;
    wire N__31682;
    wire N__31679;
    wire N__31664;
    wire N__31661;
    wire N__31660;
    wire N__31659;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31645;
    wire N__31644;
    wire N__31643;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31621;
    wire N__31614;
    wire N__31611;
    wire N__31610;
    wire N__31607;
    wire N__31602;
    wire N__31599;
    wire N__31594;
    wire N__31591;
    wire N__31580;
    wire N__31579;
    wire N__31578;
    wire N__31575;
    wire N__31574;
    wire N__31573;
    wire N__31570;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31537;
    wire N__31534;
    wire N__31531;
    wire N__31528;
    wire N__31521;
    wire N__31518;
    wire N__31517;
    wire N__31514;
    wire N__31511;
    wire N__31508;
    wire N__31505;
    wire N__31500;
    wire N__31497;
    wire N__31484;
    wire N__31481;
    wire N__31480;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31472;
    wire N__31469;
    wire N__31468;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31454;
    wire N__31451;
    wire N__31450;
    wire N__31447;
    wire N__31440;
    wire N__31437;
    wire N__31434;
    wire N__31431;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31418;
    wire N__31413;
    wire N__31410;
    wire N__31397;
    wire N__31394;
    wire N__31393;
    wire N__31390;
    wire N__31389;
    wire N__31388;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31377;
    wire N__31376;
    wire N__31373;
    wire N__31370;
    wire N__31367;
    wire N__31366;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31354;
    wire N__31351;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31338;
    wire N__31337;
    wire N__31336;
    wire N__31327;
    wire N__31324;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31302;
    wire N__31297;
    wire N__31286;
    wire N__31285;
    wire N__31284;
    wire N__31283;
    wire N__31280;
    wire N__31277;
    wire N__31276;
    wire N__31273;
    wire N__31270;
    wire N__31269;
    wire N__31268;
    wire N__31267;
    wire N__31266;
    wire N__31263;
    wire N__31262;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31222;
    wire N__31219;
    wire N__31214;
    wire N__31211;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31189;
    wire N__31178;
    wire N__31177;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31163;
    wire N__31162;
    wire N__31161;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31150;
    wire N__31149;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31124;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31076;
    wire N__31067;
    wire N__31064;
    wire N__31061;
    wire N__31060;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31052;
    wire N__31049;
    wire N__31048;
    wire N__31045;
    wire N__31042;
    wire N__31039;
    wire N__31038;
    wire N__31035;
    wire N__31034;
    wire N__31033;
    wire N__31030;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31016;
    wire N__31013;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__31001;
    wire N__31000;
    wire N__30999;
    wire N__30996;
    wire N__30991;
    wire N__30988;
    wire N__30985;
    wire N__30984;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30959;
    wire N__30956;
    wire N__30955;
    wire N__30952;
    wire N__30949;
    wire N__30946;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30920;
    wire N__30917;
    wire N__30914;
    wire N__30911;
    wire N__30908;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30900;
    wire N__30899;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30889;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30881;
    wire N__30880;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30852;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30824;
    wire N__30819;
    wire N__30816;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30790;
    wire N__30787;
    wire N__30786;
    wire N__30785;
    wire N__30782;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30774;
    wire N__30773;
    wire N__30770;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30752;
    wire N__30747;
    wire N__30744;
    wire N__30739;
    wire N__30736;
    wire N__30731;
    wire N__30728;
    wire N__30727;
    wire N__30724;
    wire N__30719;
    wire N__30714;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30683;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30675;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30667;
    wire N__30664;
    wire N__30661;
    wire N__30656;
    wire N__30653;
    wire N__30652;
    wire N__30651;
    wire N__30650;
    wire N__30649;
    wire N__30644;
    wire N__30641;
    wire N__30638;
    wire N__30635;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30605;
    wire N__30602;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30572;
    wire N__30571;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30563;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30555;
    wire N__30552;
    wire N__30551;
    wire N__30548;
    wire N__30545;
    wire N__30542;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30534;
    wire N__30533;
    wire N__30530;
    wire N__30527;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30517;
    wire N__30514;
    wire N__30509;
    wire N__30504;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30490;
    wire N__30487;
    wire N__30470;
    wire N__30467;
    wire N__30466;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30458;
    wire N__30457;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30446;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30427;
    wire N__30426;
    wire N__30423;
    wire N__30422;
    wire N__30419;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30407;
    wire N__30402;
    wire N__30399;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30362;
    wire N__30361;
    wire N__30360;
    wire N__30357;
    wire N__30354;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30346;
    wire N__30345;
    wire N__30342;
    wire N__30341;
    wire N__30338;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30315;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30281;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30241;
    wire N__30238;
    wire N__30237;
    wire N__30234;
    wire N__30233;
    wire N__30230;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30206;
    wire N__30205;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30189;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30177;
    wire N__30174;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30117;
    wire N__30112;
    wire N__30111;
    wire N__30110;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30096;
    wire N__30093;
    wire N__30090;
    wire N__30089;
    wire N__30082;
    wire N__30081;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30059;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30032;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30006;
    wire N__30005;
    wire N__30002;
    wire N__29999;
    wire N__29998;
    wire N__29997;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29983;
    wire N__29980;
    wire N__29977;
    wire N__29974;
    wire N__29971;
    wire N__29970;
    wire N__29969;
    wire N__29966;
    wire N__29961;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29931;
    wire N__29928;
    wire N__29925;
    wire N__29922;
    wire N__29919;
    wire N__29916;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29877;
    wire N__29874;
    wire N__29873;
    wire N__29872;
    wire N__29871;
    wire N__29868;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29851;
    wire N__29848;
    wire N__29845;
    wire N__29842;
    wire N__29841;
    wire N__29840;
    wire N__29833;
    wire N__29830;
    wire N__29827;
    wire N__29822;
    wire N__29819;
    wire N__29818;
    wire N__29815;
    wire N__29812;
    wire N__29807;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29759;
    wire N__29756;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29690;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29564;
    wire N__29561;
    wire N__29558;
    wire N__29557;
    wire N__29556;
    wire N__29555;
    wire N__29554;
    wire N__29551;
    wire N__29548;
    wire N__29545;
    wire N__29540;
    wire N__29535;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29507;
    wire N__29504;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29486;
    wire N__29483;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29444;
    wire N__29441;
    wire N__29438;
    wire N__29435;
    wire N__29432;
    wire N__29429;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29407;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29395;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29357;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29308;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29296;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29269;
    wire N__29266;
    wire N__29261;
    wire N__29258;
    wire N__29255;
    wire N__29252;
    wire N__29249;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29225;
    wire N__29222;
    wire N__29219;
    wire N__29216;
    wire N__29213;
    wire N__29212;
    wire N__29209;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29165;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29155;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29119;
    wire N__29116;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29063;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29051;
    wire N__29050;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29024;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29006;
    wire N__29003;
    wire N__29000;
    wire N__28997;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28973;
    wire N__28970;
    wire N__28967;
    wire N__28964;
    wire N__28961;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28943;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28904;
    wire N__28901;
    wire N__28898;
    wire N__28895;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28883;
    wire N__28880;
    wire N__28877;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28823;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28793;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28757;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28745;
    wire N__28742;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28700;
    wire N__28697;
    wire N__28694;
    wire N__28691;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28619;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28565;
    wire N__28562;
    wire N__28559;
    wire N__28556;
    wire N__28553;
    wire N__28550;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28531;
    wire N__28528;
    wire N__28523;
    wire N__28520;
    wire N__28517;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28496;
    wire N__28493;
    wire N__28490;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28445;
    wire N__28444;
    wire N__28443;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28424;
    wire N__28421;
    wire N__28418;
    wire N__28415;
    wire N__28412;
    wire N__28409;
    wire N__28406;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28391;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28372;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28357;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28337;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28322;
    wire N__28319;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28298;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28277;
    wire N__28274;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28264;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28214;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28193;
    wire N__28190;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28175;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28154;
    wire N__28151;
    wire N__28150;
    wire N__28147;
    wire N__28144;
    wire N__28141;
    wire N__28136;
    wire N__28135;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28115;
    wire N__28112;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28097;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28084;
    wire N__28081;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28064;
    wire N__28061;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28034;
    wire N__28031;
    wire N__28028;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27993;
    wire N__27990;
    wire N__27989;
    wire N__27986;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27958;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27929;
    wire N__27928;
    wire N__27927;
    wire N__27926;
    wire N__27925;
    wire N__27924;
    wire N__27923;
    wire N__27922;
    wire N__27911;
    wire N__27904;
    wire N__27899;
    wire N__27896;
    wire N__27893;
    wire N__27892;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27878;
    wire N__27877;
    wire N__27874;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27857;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27836;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27745;
    wire N__27742;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27715;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27680;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27653;
    wire N__27650;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27527;
    wire N__27524;
    wire N__27521;
    wire N__27518;
    wire N__27515;
    wire N__27512;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27479;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27464;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27443;
    wire N__27440;
    wire N__27437;
    wire N__27434;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27344;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27164;
    wire N__27161;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27095;
    wire N__27094;
    wire N__27093;
    wire N__27092;
    wire N__27091;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27073;
    wire N__27062;
    wire N__27061;
    wire N__27058;
    wire N__27057;
    wire N__27054;
    wire N__27051;
    wire N__27046;
    wire N__27043;
    wire N__27040;
    wire N__27037;
    wire N__27034;
    wire N__27031;
    wire N__27028;
    wire N__27023;
    wire N__27022;
    wire N__27021;
    wire N__27020;
    wire N__27019;
    wire N__27016;
    wire N__27015;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26992;
    wire N__26989;
    wire N__26984;
    wire N__26981;
    wire N__26978;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26950;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26933;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26900;
    wire N__26897;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26855;
    wire N__26852;
    wire N__26849;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26810;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26798;
    wire N__26795;
    wire N__26792;
    wire N__26789;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26744;
    wire N__26741;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26723;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26687;
    wire N__26684;
    wire N__26681;
    wire N__26678;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26666;
    wire N__26663;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26639;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26615;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26582;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26563;
    wire N__26562;
    wire N__26559;
    wire N__26556;
    wire N__26553;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26516;
    wire N__26513;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26389;
    wire N__26386;
    wire N__26383;
    wire N__26380;
    wire N__26377;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26197;
    wire N__26196;
    wire N__26195;
    wire N__26194;
    wire N__26193;
    wire N__26188;
    wire N__26185;
    wire N__26184;
    wire N__26179;
    wire N__26178;
    wire N__26175;
    wire N__26174;
    wire N__26171;
    wire N__26168;
    wire N__26167;
    wire N__26166;
    wire N__26165;
    wire N__26164;
    wire N__26163;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26137;
    wire N__26134;
    wire N__26131;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26099;
    wire N__26098;
    wire N__26095;
    wire N__26092;
    wire N__26091;
    wire N__26090;
    wire N__26089;
    wire N__26088;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26078;
    wire N__26073;
    wire N__26068;
    wire N__26065;
    wire N__26062;
    wire N__26059;
    wire N__26048;
    wire N__26045;
    wire N__26044;
    wire N__26043;
    wire N__26042;
    wire N__26041;
    wire N__26038;
    wire N__26031;
    wire N__26028;
    wire N__26027;
    wire N__26024;
    wire N__26019;
    wire N__26016;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25945;
    wire N__25942;
    wire N__25939;
    wire N__25936;
    wire N__25933;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25823;
    wire N__25820;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25664;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25522;
    wire N__25521;
    wire N__25520;
    wire N__25517;
    wire N__25510;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25478;
    wire N__25475;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25453;
    wire N__25450;
    wire N__25447;
    wire N__25444;
    wire N__25439;
    wire N__25436;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25421;
    wire N__25418;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25369;
    wire N__25368;
    wire N__25367;
    wire N__25366;
    wire N__25365;
    wire N__25364;
    wire N__25363;
    wire N__25362;
    wire N__25361;
    wire N__25360;
    wire N__25359;
    wire N__25358;
    wire N__25357;
    wire N__25356;
    wire N__25355;
    wire N__25354;
    wire N__25353;
    wire N__25352;
    wire N__25351;
    wire N__25350;
    wire N__25349;
    wire N__25348;
    wire N__25347;
    wire N__25340;
    wire N__25331;
    wire N__25322;
    wire N__25311;
    wire N__25302;
    wire N__25293;
    wire N__25288;
    wire N__25281;
    wire N__25274;
    wire N__25271;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25259;
    wire N__25256;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25206;
    wire N__25203;
    wire N__25200;
    wire N__25197;
    wire N__25194;
    wire N__25187;
    wire N__25184;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25160;
    wire N__25159;
    wire N__25158;
    wire N__25153;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25138;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25022;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24950;
    wire N__24947;
    wire N__24944;
    wire N__24941;
    wire N__24938;
    wire N__24935;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24920;
    wire N__24917;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24693;
    wire N__24692;
    wire N__24691;
    wire N__24686;
    wire N__24683;
    wire N__24682;
    wire N__24677;
    wire N__24672;
    wire N__24669;
    wire N__24668;
    wire N__24667;
    wire N__24664;
    wire N__24659;
    wire N__24656;
    wire N__24653;
    wire N__24652;
    wire N__24651;
    wire N__24650;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24638;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24550;
    wire N__24547;
    wire N__24544;
    wire N__24543;
    wire N__24538;
    wire N__24535;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24513;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24499;
    wire N__24496;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24461;
    wire N__24460;
    wire N__24459;
    wire N__24456;
    wire N__24455;
    wire N__24454;
    wire N__24451;
    wire N__24448;
    wire N__24445;
    wire N__24442;
    wire N__24439;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24399;
    wire N__24392;
    wire N__24389;
    wire N__24388;
    wire N__24387;
    wire N__24386;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24363;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24349;
    wire N__24346;
    wire N__24339;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24304;
    wire N__24301;
    wire N__24298;
    wire N__24295;
    wire N__24290;
    wire N__24287;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24256;
    wire N__24255;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24243;
    wire N__24240;
    wire N__24235;
    wire N__24232;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24158;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24119;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24083;
    wire N__24080;
    wire N__24077;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23836;
    wire N__23835;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23824;
    wire N__23823;
    wire N__23820;
    wire N__23817;
    wire N__23814;
    wire N__23805;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23719;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23711;
    wire N__23708;
    wire N__23707;
    wire N__23706;
    wire N__23705;
    wire N__23704;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23688;
    wire N__23683;
    wire N__23678;
    wire N__23675;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23656;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23645;
    wire N__23642;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23623;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23608;
    wire N__23607;
    wire N__23606;
    wire N__23603;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23570;
    wire N__23567;
    wire N__23566;
    wire N__23565;
    wire N__23562;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23554;
    wire N__23551;
    wire N__23550;
    wire N__23547;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23528;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23494;
    wire N__23491;
    wire N__23490;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23464;
    wire N__23463;
    wire N__23462;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23449;
    wire N__23446;
    wire N__23445;
    wire N__23434;
    wire N__23431;
    wire N__23428;
    wire N__23423;
    wire N__23422;
    wire N__23419;
    wire N__23418;
    wire N__23417;
    wire N__23414;
    wire N__23413;
    wire N__23410;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23354;
    wire N__23345;
    wire N__23344;
    wire N__23341;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23299;
    wire N__23298;
    wire N__23295;
    wire N__23294;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23274;
    wire N__23267;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23237;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23188;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23132;
    wire N__23129;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23117;
    wire N__23114;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23084;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23072;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23060;
    wire N__23057;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23045;
    wire N__23042;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23030;
    wire N__23027;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23015;
    wire N__23012;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23000;
    wire N__22997;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22985;
    wire N__22982;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22970;
    wire N__22967;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22955;
    wire N__22952;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22940;
    wire N__22939;
    wire N__22938;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22894;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22880;
    wire N__22877;
    wire N__22876;
    wire N__22873;
    wire N__22870;
    wire N__22867;
    wire N__22862;
    wire N__22859;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22847;
    wire N__22844;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22832;
    wire N__22829;
    wire N__22828;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22813;
    wire N__22810;
    wire N__22807;
    wire N__22802;
    wire N__22799;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22762;
    wire N__22759;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22716;
    wire N__22711;
    wire N__22708;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22663;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22625;
    wire N__22622;
    wire N__22621;
    wire N__22616;
    wire N__22613;
    wire N__22612;
    wire N__22611;
    wire N__22610;
    wire N__22609;
    wire N__22604;
    wire N__22599;
    wire N__22596;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22555;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22529;
    wire N__22526;
    wire N__22523;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22469;
    wire N__22466;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22454;
    wire N__22451;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22439;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22427;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22415;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22403;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21994;
    wire N__21993;
    wire N__21992;
    wire N__21991;
    wire N__21988;
    wire N__21983;
    wire N__21978;
    wire N__21971;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21959;
    wire N__21958;
    wire N__21955;
    wire N__21952;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21919;
    wire N__21918;
    wire N__21917;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21889;
    wire N__21888;
    wire N__21881;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21845;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21570;
    wire N__21567;
    wire N__21564;
    wire N__21563;
    wire N__21560;
    wire N__21555;
    wire N__21552;
    wire N__21545;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21530;
    wire N__21527;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21512;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21504;
    wire N__21503;
    wire N__21498;
    wire N__21495;
    wire N__21494;
    wire N__21491;
    wire N__21486;
    wire N__21483;
    wire N__21476;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21458;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21446;
    wire N__21445;
    wire N__21442;
    wire N__21439;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21421;
    wire N__21418;
    wire N__21417;
    wire N__21416;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21402;
    wire N__21401;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21387;
    wire N__21384;
    wire N__21379;
    wire N__21376;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21331;
    wire N__21328;
    wire N__21327;
    wire N__21326;
    wire N__21321;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21305;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21297;
    wire N__21296;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21284;
    wire N__21283;
    wire N__21282;
    wire N__21277;
    wire N__21274;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21254;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21194;
    wire N__21191;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21176;
    wire N__21173;
    wire N__21172;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21158;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21143;
    wire N__21140;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21089;
    wire N__21088;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21066;
    wire N__21065;
    wire N__21064;
    wire N__21059;
    wire N__21056;
    wire N__21051;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21028;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21011;
    wire N__21010;
    wire N__21007;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20983;
    wire N__20982;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20966;
    wire N__20965;
    wire N__20962;
    wire N__20961;
    wire N__20958;
    wire N__20955;
    wire N__20952;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20935;
    wire N__20932;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20919;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20905;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20864;
    wire N__20861;
    wire N__20860;
    wire N__20857;
    wire N__20854;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20842;
    wire N__20839;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20770;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20760;
    wire N__20753;
    wire N__20752;
    wire N__20751;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20739;
    wire N__20732;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20720;
    wire N__20719;
    wire N__20718;
    wire N__20711;
    wire N__20710;
    wire N__20709;
    wire N__20708;
    wire N__20707;
    wire N__20706;
    wire N__20703;
    wire N__20692;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20682;
    wire N__20677;
    wire N__20672;
    wire N__20671;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20651;
    wire N__20650;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20627;
    wire N__20626;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20582;
    wire N__20579;
    wire N__20578;
    wire N__20577;
    wire N__20572;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20559;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20545;
    wire N__20542;
    wire N__20541;
    wire N__20540;
    wire N__20539;
    wire N__20538;
    wire N__20537;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20523;
    wire N__20516;
    wire N__20507;
    wire N__20506;
    wire N__20505;
    wire N__20500;
    wire N__20497;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20425;
    wire N__20424;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20365;
    wire N__20364;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20285;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire cs_rpi2flash_c;
    wire clk_c;
    wire \pll128M2_inst.pll_clk64_0 ;
    wire \pll128M2_inst.pll_clk128 ;
    wire VCCG0;
    wire bfn_1_11_0_;
    wire sRAM_pointer_write_cry_0;
    wire sRAM_pointer_write_cry_1;
    wire sRAM_pointer_write_cry_2;
    wire sRAM_pointer_write_cry_3;
    wire sRAM_pointer_write_cry_4;
    wire sRAM_pointer_write_cry_5;
    wire sRAM_pointer_write_cry_6;
    wire sRAM_pointer_write_cry_7;
    wire bfn_1_12_0_;
    wire sRAM_pointer_write_cry_8;
    wire sRAM_pointer_write_cry_9;
    wire sRAM_pointer_write_cry_10;
    wire sRAM_pointer_write_cry_11;
    wire sRAM_pointer_write_cry_12;
    wire sRAM_pointer_write_cry_13;
    wire sRAM_pointer_write_cry_14;
    wire sRAM_pointer_write_cry_15;
    wire bfn_1_13_0_;
    wire sRAM_pointer_write_cry_16;
    wire sRAM_pointer_write_cry_17;
    wire N_1487_g;
    wire \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.N_1531_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1 ;
    wire button_mode_c;
    wire button_mode_ibuf_RNIN5KZ0Z7;
    wire DAC_cs_c;
    wire bfn_3_6_0_;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_s_1 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_s_0 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i ;
    wire \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0 ;
    wire bfn_3_8_0_;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_0 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_1 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_2 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_3 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_4 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_5 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_6 ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3 ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3 ;
    wire \spi_master_inst.sclk_gen_u0.N_1531 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_start_iZ0 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_start_i_i ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2 ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.N_48_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.N_36 ;
    wire \spi_master_inst.sclk_gen_u0.N_5 ;
    wire \spi_master_inst.sclk_gen_u0.N_150_0 ;
    wire \spi_master_inst.sclk_gen_u0.N_48 ;
    wire \spi_master_inst.spi_data_path_u1.N_1414_cascade_ ;
    wire \spi_master_inst.spi_data_path_u1.N_1415_cascade_ ;
    wire DAC_mosi_c;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_ ;
    wire \spi_master_inst.spi_data_path_u1.N_1421_cascade_ ;
    wire \spi_master_inst.spi_data_path_u1.N_1422 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4 ;
    wire \spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6 ;
    wire DAC_sclk_c;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4 ;
    wire \spi_master_inst.sclk_gen_u0.N_1737 ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4 ;
    wire \spi_master_inst.sclk_gen_u0.N_1737_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0 ;
    wire \spi_master_inst.sclk_gen_u0.N_1540 ;
    wire \spi_master_inst.ss_start_i ;
    wire \spi_master_inst.spi_data_path_u1.N_1411 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14 ;
    wire \spi_master_inst.spi_data_path_u1.N_1418 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6 ;
    wire bfn_6_7_0_;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1 ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2 ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3 ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4 ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO ;
    wire bfn_6_8_0_;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6 ;
    wire \spi_master_inst.o_sclk_RNIH6AC ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3 ;
    wire spi_mosi_ready64_prevZ0Z2;
    wire spi_mosi_ready64_prevZ0;
    wire spi_mosi_ready64_prevZ0Z3;
    wire spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_;
    wire bfn_6_12_0_;
    wire sEETrigCounterZ0Z_1;
    wire un8_trig_prev_0_cry_0;
    wire sEETrigCounterZ0Z_2;
    wire un8_trig_prev_0_cry_1;
    wire sEETrigCounterZ0Z_3;
    wire un8_trig_prev_0_cry_2;
    wire sEETrigCounterZ0Z_4;
    wire un8_trig_prev_0_cry_3;
    wire sEETrigCounterZ0Z_5;
    wire un8_trig_prev_0_cry_4;
    wire sEETrigCounterZ0Z_6;
    wire un8_trig_prev_0_cry_5;
    wire sEETrigCounterZ0Z_7;
    wire un8_trig_prev_0_cry_6;
    wire un8_trig_prev_0_cry_7;
    wire bfn_6_13_0_;
    wire un8_trig_prev_0_cry_8;
    wire un8_trig_prev_0_cry_9;
    wire un8_trig_prev_0_cry_10;
    wire un8_trig_prev_0_cry_11;
    wire un8_trig_prev_0_cry_12;
    wire un8_trig_prev_0_cry_13;
    wire un8_trig_prev_0_cry_14;
    wire sEETrigCounterZ0Z_10;
    wire sEETrigCounterZ0Z_11;
    wire sEETrigCounterZ0Z_12;
    wire sEETrigCounterZ0Z_13;
    wire sEETrigCounterZ0Z_14;
    wire sEETrigCounterZ0Z_15;
    wire sEETrigCounterZ0Z_8;
    wire sEETrigCounterZ0Z_9;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_6 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_5 ;
    wire N_316_cascade_;
    wire N_317_cascade_;
    wire sAddress_RNI8U0V1Z0Z_1_cascade_;
    wire sAddress_RNI8U0V1Z0Z_1;
    wire N_454_cascade_;
    wire N_346_i_cascade_;
    wire un1_spointer11_8_0_0_a2_1_cascade_;
    wire sAddress_RNI7G5E2Z0Z_6;
    wire sAddressZ0Z_7;
    wire sAddressZ0Z_6;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0 ;
    wire bfn_7_10_0_;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1 ;
    wire \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2 ;
    wire \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1 ;
    wire \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2 ;
    wire \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3 ;
    wire \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5 ;
    wire \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ;
    wire spi_mosi_ready;
    wire spi_mosi_ready_prevZ0;
    wire spi_mosi_ready_prevZ0Z2;
    wire spi_mosi_ready_prevZ0Z3;
    wire un8_trig_prev_0;
    wire un10_trig_prev_0;
    wire sTrigCounter_i_0;
    wire bfn_7_12_0_;
    wire un10_trig_prev_1;
    wire sTrigCounter_i_1;
    wire un10_trig_prev_cry_0;
    wire un10_trig_prev_2;
    wire sTrigCounter_i_2;
    wire un10_trig_prev_cry_1;
    wire un10_trig_prev_3;
    wire sTrigCounter_i_3;
    wire un10_trig_prev_cry_2;
    wire un10_trig_prev_4;
    wire sTrigCounter_i_4;
    wire un10_trig_prev_cry_3;
    wire un10_trig_prev_5;
    wire sTrigCounter_i_5;
    wire un10_trig_prev_cry_4;
    wire un10_trig_prev_6;
    wire sTrigCounter_i_6;
    wire un10_trig_prev_cry_5;
    wire un10_trig_prev_7;
    wire sTrigCounter_i_7;
    wire un10_trig_prev_cry_6;
    wire un10_trig_prev_cry_7;
    wire un10_trig_prev_8;
    wire sTrigCounter_i_8;
    wire bfn_7_13_0_;
    wire un10_trig_prev_9;
    wire sTrigCounter_i_9;
    wire un10_trig_prev_cry_8;
    wire un10_trig_prev_10;
    wire sTrigCounter_i_10;
    wire un10_trig_prev_cry_9;
    wire un10_trig_prev_11;
    wire sTrigCounter_i_11;
    wire un10_trig_prev_cry_10;
    wire un10_trig_prev_12;
    wire sTrigCounter_i_12;
    wire un10_trig_prev_cry_11;
    wire un10_trig_prev_13;
    wire sTrigCounter_i_13;
    wire un10_trig_prev_cry_12;
    wire un10_trig_prev_14;
    wire sTrigCounter_i_14;
    wire un10_trig_prev_cry_13;
    wire un10_trig_prev_15;
    wire sTrigCounter_i_15;
    wire un10_trig_prev_cry_14;
    wire un10_trig_prev_cry_15;
    wire bfn_7_14_0_;
    wire N_173;
    wire \INVspi_slave_inst.rx_done_neg_sclk_iC_net ;
    wire sEEADC_freqZ0Z_4;
    wire un3_trig_0;
    wire sEEADC_freqZ0Z_5;
    wire spi_mosi_rpi_c;
    wire spi_mosi_ft_c;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7 ;
    wire sDAC_mem_11_1_sqmuxa;
    wire N_344_cascade_;
    wire sDAC_mem_35_1_sqmuxa;
    wire sEESingleCont_RNOZ0Z_0;
    wire sEESingleContZ0;
    wire N_1631;
    wire sEETrigInternal_3_iv_0_0_i_0;
    wire \spi_slave_inst.rx_done_neg_sclk_iZ0 ;
    wire \spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541 ;
    wire \spi_slave_inst.rx_done_reg1_iZ0 ;
    wire N_319_cascade_;
    wire sAddress_RNI9IH12_2Z0Z_1;
    wire \spi_slave_inst.rx_done_reg2_iZ0 ;
    wire \spi_slave_inst.rx_done_reg3_iZ0 ;
    wire \spi_slave_inst.rx_ready_i_RNOZ0Z_0 ;
    wire sPointer_RNI5LBD1Z0Z_0_cascade_;
    wire sDAC_mem_17_1_sqmuxa_0_a2_0_a2_1_0;
    wire sAddressZ0Z_4;
    wire sAddress_RNIP2UK1Z0Z_4_cascade_;
    wire trig_rpi_c;
    wire trig_ext_c;
    wire trig_ft_c;
    wire trig_prevZ0;
    wire g3_0_cascade_;
    wire sAddress_RNI70I7Z0Z_1_cascade_;
    wire g1_i_a4_0_0;
    wire N_8_mux;
    wire un10_trig_prev_cry_15_THRU_CO;
    wire N_178;
    wire un1_scounter_i_0;
    wire N_178_cascade_;
    wire N_96;
    wire N_77_cascade_;
    wire sPeriod_prevZ0;
    wire un1_reset_rpi_inv_2_0;
    wire bfn_8_13_0_;
    wire un1_sTrigCounter_cry_0;
    wire sTrigCounterZ0Z_2;
    wire un1_sTrigCounter_cry_1;
    wire sTrigCounterZ0Z_3;
    wire un1_sTrigCounter_cry_2;
    wire sTrigCounterZ0Z_4;
    wire un1_sTrigCounter_cry_3;
    wire sTrigCounterZ0Z_5;
    wire un1_sTrigCounter_cry_4;
    wire sTrigCounterZ0Z_6;
    wire un1_sTrigCounter_cry_5;
    wire sTrigCounterZ0Z_7;
    wire un1_sTrigCounter_cry_6;
    wire un1_sTrigCounter_cry_7;
    wire sTrigCounterZ0Z_8;
    wire bfn_8_14_0_;
    wire sTrigCounterZ0Z_9;
    wire un1_sTrigCounter_cry_8;
    wire sTrigCounterZ0Z_10;
    wire un1_sTrigCounter_cry_9;
    wire sTrigCounterZ0Z_11;
    wire un1_sTrigCounter_cry_10;
    wire sTrigCounterZ0Z_12;
    wire un1_sTrigCounter_cry_11;
    wire sTrigCounterZ0Z_13;
    wire un1_sTrigCounter_cry_12;
    wire sTrigCounterZ0Z_14;
    wire un1_sTrigCounter_cry_13;
    wire un1_sTrigCounter_cry_14;
    wire sTrigCounterZ0Z_15;
    wire N_82_i;
    wire sDAC_mem_29_1_sqmuxa;
    wire sEEPon_1_sqmuxa;
    wire \spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0 ;
    wire \spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0 ;
    wire \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0 ;
    wire \spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10 ;
    wire sDAC_mem_38_1_sqmuxa;
    wire sAddress_RNI6VH7_3Z0Z_1;
    wire sAddress_RNI6VH7_3Z0Z_1_cascade_;
    wire sDAC_mem_10_1_sqmuxa;
    wire N_326_cascade_;
    wire LED_ACQ_obuf_RNOZ0;
    wire sAddress_RNIAM2A_0Z0Z_1_cascade_;
    wire N_445_cascade_;
    wire sAddress_RNI6VH7_5Z0Z_1;
    wire N_445;
    wire N_316;
    wire un1_spointer11_0;
    wire sAddress_RNI6VH7_2Z0Z_1;
    wire sEETrigInternalZ0;
    wire g3_0;
    wire sEETrigInternal_prevZ0;
    wire LED_MODE_c;
    wire N_831_16_cascade_;
    wire N_319;
    wire g0_13_cascade_;
    wire g0_1_0;
    wire g0_15_0;
    wire g0_13_1;
    wire g0_17_0;
    wire N_326;
    wire g0_16_0;
    wire g1_i_a4_6;
    wire g1_i_a4_5_cascade_;
    wire un1_reset_rpi_inv_2_0_o2_5;
    wire g1_i_a4_9_cascade_;
    wire sEETrigInternal_prev_RNIH3OJZ0Z1;
    wire g0_0_1;
    wire g0_16;
    wire g0_11;
    wire g0_14;
    wire sDAC_mem_30_1_sqmuxa;
    wire sEEPonZ0Z_0;
    wire sEEPon_i_0;
    wire bfn_9_17_0_;
    wire sEEPonZ0Z_1;
    wire sEEPon_i_1;
    wire un7_spon_cry_0;
    wire sEEPonZ0Z_2;
    wire sEEPon_i_2;
    wire un7_spon_cry_1;
    wire sEEPonZ0Z_3;
    wire sEEPon_i_3;
    wire un7_spon_cry_2;
    wire sEEPonZ0Z_4;
    wire sEEPon_i_4;
    wire un7_spon_cry_3;
    wire sEEPonZ0Z_5;
    wire sEEPon_i_5;
    wire un7_spon_cry_4;
    wire sEEPonZ0Z_6;
    wire sEEPon_i_6;
    wire un7_spon_cry_5;
    wire sEEPonZ0Z_7;
    wire sEEPon_i_7;
    wire un7_spon_cry_6;
    wire un7_spon_cry_7;
    wire bfn_9_18_0_;
    wire un7_spon_cry_8;
    wire un7_spon_cry_9;
    wire un7_spon_cry_10;
    wire un7_spon_cry_11;
    wire un7_spon_cry_12;
    wire un7_spon_cry_13;
    wire un7_spon_cry_14;
    wire un7_spon_cry_15;
    wire bfn_9_19_0_;
    wire un7_spon_cry_16;
    wire un7_spon_cry_17;
    wire un7_spon_cry_18;
    wire un7_spon_cry_19;
    wire un7_spon_cry_20;
    wire un7_spon_cry_21;
    wire un7_spon_cry_22;
    wire un7_spon_cry_23;
    wire bfn_9_20_0_;
    wire pon_obuf_RNOZ0;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_0 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_1 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_10 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_11 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_13 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_14 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_15 ;
    wire sDAC_mem_42_1_sqmuxa;
    wire sDAC_mem_14_1_sqmuxa;
    wire sAddress_RNI9IH12Z0Z_0;
    wire sAddress_RNI9IH12_1Z0Z_2;
    wire sDAC_mem_15_1_sqmuxa;
    wire un21_trig_prev_21_5;
    wire op_gt_op_gt_un13_striginternallto23_5_cascade_;
    wire un1_reset_rpi_inv_2_0_o2_2;
    wire g0_13_0;
    wire un21_trig_prev_21_4;
    wire g0_6;
    wire N_99;
    wire op_gt_op_gt_un13_striginternallto23_3;
    wire N_831_16;
    wire op_gt_op_gt_un13_striginternallto23_6;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2 ;
    wire \spi_master_inst.sclk_gen_u0.N_158_7 ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ;
    wire \spi_master_inst.sclk_gen_u0.spi_start_iZ0 ;
    wire \spi_master_inst.sclk_gen_u0.N_158_7_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ;
    wire \spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0 ;
    wire g2_6;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_i6_3 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_i6 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_ ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_3 ;
    wire \spi_slave_inst.un23_i_ssn_3_cascade_ ;
    wire \spi_slave_inst.un23_i_ssn_cascade_ ;
    wire g0_10;
    wire g0_10_0;
    wire sDAC_mem_31_1_sqmuxa;
    wire sAddress_RNIA6242_4Z0Z_0;
    wire sAddress_RNIA6242Z0Z_0;
    wire LED3_c_i;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15 ;
    wire sDAC_dataZ0Z_0;
    wire sDAC_dataZ0Z_1;
    wire sDAC_dataZ0Z_11;
    wire sDAC_dataZ0Z_12;
    wire sDAC_dataZ0Z_13;
    wire sDAC_dataZ0Z_14;
    wire sDAC_dataZ0Z_15;
    wire sAddress_RNIETI62Z0Z_1;
    wire sEEPeriodZ0Z_0;
    wire sEEPeriod_i_0;
    wire bfn_11_6_0_;
    wire sEEPeriodZ0Z_1;
    wire sEEPeriod_i_1;
    wire un4_speriod_cry_0;
    wire sEEPeriodZ0Z_2;
    wire sEEPeriod_i_2;
    wire un4_speriod_cry_1;
    wire sEEPeriodZ0Z_3;
    wire sEEPeriod_i_3;
    wire un4_speriod_cry_2;
    wire sEEPeriodZ0Z_4;
    wire sEEPeriod_i_4;
    wire un4_speriod_cry_3;
    wire sEEPeriodZ0Z_5;
    wire sEEPeriod_i_5;
    wire un4_speriod_cry_4;
    wire sEEPeriodZ0Z_6;
    wire sEEPeriod_i_6;
    wire un4_speriod_cry_5;
    wire sEEPeriodZ0Z_7;
    wire sEEPeriod_i_7;
    wire un4_speriod_cry_6;
    wire un4_speriod_cry_7;
    wire sEEPeriodZ0Z_8;
    wire sEEPeriod_i_8;
    wire bfn_11_7_0_;
    wire sEEPeriodZ0Z_9;
    wire sEEPeriod_i_9;
    wire un4_speriod_cry_8;
    wire sEEPeriodZ0Z_10;
    wire sEEPeriod_i_10;
    wire un4_speriod_cry_9;
    wire sEEPeriodZ0Z_11;
    wire sEEPeriod_i_11;
    wire un4_speriod_cry_10;
    wire sEEPeriodZ0Z_12;
    wire sEEPeriod_i_12;
    wire un4_speriod_cry_11;
    wire sEEPeriodZ0Z_13;
    wire sEEPeriod_i_13;
    wire un4_speriod_cry_12;
    wire sEEPeriodZ0Z_14;
    wire sEEPeriod_i_14;
    wire un4_speriod_cry_13;
    wire sEEPeriodZ0Z_15;
    wire sEEPeriod_i_15;
    wire un4_speriod_cry_14;
    wire un4_speriod_cry_15;
    wire sEEPeriodZ0Z_16;
    wire sEEPeriod_i_16;
    wire bfn_11_8_0_;
    wire sEEPeriodZ0Z_17;
    wire sEEPeriod_i_17;
    wire un4_speriod_cry_16;
    wire sEEPeriodZ0Z_18;
    wire sEEPeriod_i_18;
    wire un4_speriod_cry_17;
    wire sEEPeriodZ0Z_19;
    wire sEEPeriod_i_19;
    wire un4_speriod_cry_18;
    wire sEEPeriodZ0Z_20;
    wire sEEPeriod_i_20;
    wire un4_speriod_cry_19;
    wire sEEPeriodZ0Z_21;
    wire sEEPeriod_i_21;
    wire un4_speriod_cry_20;
    wire sEEPeriodZ0Z_22;
    wire sEEPeriod_i_22;
    wire un4_speriod_cry_21;
    wire sEEPeriodZ0Z_23;
    wire sEEPeriod_i_23;
    wire un4_speriod_cry_22;
    wire un4_speriod_cry_23;
    wire bfn_11_9_0_;
    wire un1_spointer11_2_0_0_a2_6;
    wire un1_spointer11_2_0_0_a2_1;
    wire sTrigInternalZ0;
    wire op_gt_op_gt_un13_striginternal_0;
    wire un4_speriod_cry_23_THRU_CO;
    wire bfn_11_10_0_;
    wire sCounter_cry_0;
    wire sCounter_cry_1;
    wire sCounter_cry_2;
    wire sCounter_cry_3;
    wire sCounter_cry_4;
    wire sCounter_cry_5;
    wire sCounter_cry_6;
    wire sCounter_cry_7;
    wire bfn_11_11_0_;
    wire sCounter_cry_8;
    wire sCounter_cry_9;
    wire sCounter_cry_10;
    wire sCounter_cry_11;
    wire sCounter_cry_12;
    wire sCounter_cry_13;
    wire sCounter_cry_14;
    wire sCounter_cry_15;
    wire bfn_11_12_0_;
    wire sCounter_cry_16;
    wire sCounter_cry_17;
    wire sCounter_cry_18;
    wire sCounter_cry_19;
    wire sCounter_cry_20;
    wire sCounter_cry_21;
    wire LED_ACQ_c_i;
    wire sCounter_cry_22;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0 ;
    wire bfn_11_13_0_;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7 ;
    wire un1_spointer11_5_0_2;
    wire sAddress_RNIA6242_3Z0Z_0;
    wire sEEDelayACQZ0Z_0;
    wire sEEDelayACQ_i_0;
    wire bfn_11_17_0_;
    wire sEEDelayACQZ0Z_1;
    wire sEEDelayACQ_i_1;
    wire un4_sacqtime_cry_0;
    wire sEEDelayACQZ0Z_2;
    wire sEEDelayACQ_i_2;
    wire un4_sacqtime_cry_1;
    wire sEEDelayACQZ0Z_3;
    wire sEEDelayACQ_i_3;
    wire un4_sacqtime_cry_2;
    wire sEEDelayACQZ0Z_4;
    wire sEEDelayACQ_i_4;
    wire un4_sacqtime_cry_3;
    wire sEEDelayACQZ0Z_5;
    wire sEEDelayACQ_i_5;
    wire un4_sacqtime_cry_4;
    wire sEEDelayACQZ0Z_6;
    wire sEEDelayACQ_i_6;
    wire un4_sacqtime_cry_5;
    wire sEEDelayACQZ0Z_7;
    wire sEEDelayACQ_i_7;
    wire un4_sacqtime_cry_6;
    wire un4_sacqtime_cry_7;
    wire sEEDelayACQZ0Z_8;
    wire sEEDelayACQ_i_8;
    wire bfn_11_18_0_;
    wire sEEDelayACQZ0Z_9;
    wire sEEDelayACQ_i_9;
    wire un4_sacqtime_cry_8;
    wire sEEDelayACQZ0Z_10;
    wire sEEDelayACQ_i_10;
    wire un4_sacqtime_cry_9;
    wire sEEDelayACQZ0Z_11;
    wire sEEDelayACQ_i_11;
    wire un4_sacqtime_cry_10;
    wire sEEDelayACQZ0Z_12;
    wire sEEDelayACQ_i_12;
    wire un4_sacqtime_cry_11;
    wire sEEDelayACQZ0Z_13;
    wire sEEDelayACQ_i_13;
    wire un4_sacqtime_cry_12;
    wire sEEDelayACQZ0Z_14;
    wire sEEDelayACQ_i_14;
    wire un4_sacqtime_cry_13;
    wire sEEDelayACQZ0Z_15;
    wire sEEDelayACQ_i_15;
    wire un4_sacqtime_cry_14;
    wire un4_sacqtime_cry_15;
    wire bfn_11_19_0_;
    wire un4_sacqtime_cry_16;
    wire un4_sacqtime_cry_17;
    wire un4_sacqtime_cry_18;
    wire un4_sacqtime_cry_19;
    wire g1_i_a4_4;
    wire un4_sacqtime_cry_20;
    wire un4_sacqtime_cry_21;
    wire g0_4_0;
    wire un4_sacqtime_cry_22;
    wire un4_sacqtime_cry_23;
    wire bfn_11_20_0_;
    wire spi_sclk_ft_c;
    wire spi_sclk_rpi_c;
    wire spi_sclk;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_12 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9 ;
    wire sDAC_mem_35Z0Z_3;
    wire sDAC_data_2_6_bm_1_6_cascade_;
    wire sDAC_mem_3Z0Z_3;
    wire sDAC_mem_8Z0Z_3;
    wire sDAC_data_2_20_am_1_6_cascade_;
    wire sDAC_mem_10Z0Z_3;
    wire sDAC_mem_42Z0Z_3;
    wire sDAC_data_RNO_17Z0Z_6_cascade_;
    wire sDAC_mem_11Z0Z_3;
    wire sDAC_data_RNO_8Z0Z_6_cascade_;
    wire sDAC_data_RNO_7Z0Z_6;
    wire sDAC_mem_2Z0Z_3;
    wire sDAC_mem_7Z0Z_1;
    wire un1_spointer11_2_0_0_a2_5;
    wire N_183;
    wire sPointerZ0Z_1;
    wire sPointerZ0Z_0;
    wire spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1;
    wire N_1624;
    wire sDAC_mem_34Z0Z_3;
    wire sDAC_mem_34_1_sqmuxa;
    wire sDAC_mem_39Z0Z_1;
    wire sDAC_mem_39_1_sqmuxa;
    wire sEEPoffZ0Z_0;
    wire bfn_12_10_0_;
    wire sEEPoffZ0Z_1;
    wire un1_spoff_cry_0;
    wire sEEPoffZ0Z_2;
    wire un1_spoff_cry_1;
    wire sEEPoffZ0Z_3;
    wire un1_spoff_cry_2;
    wire sEEPoffZ0Z_4;
    wire un1_spoff_cry_3;
    wire sEEPoffZ0Z_5;
    wire un1_spoff_cry_4;
    wire sEEPoffZ0Z_6;
    wire un1_spoff_cry_5;
    wire sEEPoffZ0Z_7;
    wire un1_spoff_cry_6;
    wire un1_spoff_cry_7;
    wire bfn_12_11_0_;
    wire un1_spoff_cry_8;
    wire sEEPoffZ0Z_10;
    wire un1_spoff_cry_9;
    wire un1_spoff_cry_10;
    wire un1_spoff_cry_11;
    wire un1_spoff_cry_12;
    wire un1_spoff_cry_13;
    wire un1_spoff_cry_14;
    wire un1_spoff_cry_15;
    wire sCounter_i_16;
    wire bfn_12_12_0_;
    wire sCounter_i_17;
    wire un1_spoff_cry_16;
    wire sCounter_i_18;
    wire un1_spoff_cry_17;
    wire sCounter_i_19;
    wire un1_spoff_cry_18;
    wire sCounter_i_20;
    wire un1_spoff_cry_19;
    wire sCounter_i_21;
    wire un1_spoff_cry_20;
    wire sCounter_i_22;
    wire un1_spoff_cry_21;
    wire sCounter_i_23;
    wire un1_spoff_cry_22;
    wire un1_spoff_cry_23;
    wire bfn_12_13_0_;
    wire N_1683_i;
    wire sbuttonModeStatusZ0;
    wire sbuttonModeStatus_0_sqmuxa_0;
    wire sbuttonModeStatus_0_sqmuxa_18;
    wire sAddress_RNIA6242_1Z0Z_0;
    wire sAddress_RNIA6242_0Z0Z_0;
    wire sEEPoffZ0Z_11;
    wire sEEPoffZ0Z_12;
    wire sEEPoffZ0Z_13;
    wire sEEPoffZ0Z_14;
    wire sEEPoffZ0Z_15;
    wire sEEPoffZ0Z_8;
    wire sEEPoffZ0Z_9;
    wire sAddress_RNIA6242_2Z0Z_0;
    wire un4_sacqtime_cry_23_c_RNI2CQMZ0;
    wire ADC5_c;
    wire RAM_DATA_1Z0Z_5;
    wire ADC1_c;
    wire RAM_DATA_1Z0Z_1;
    wire ADC9_c;
    wire RAM_DATA_1Z0Z_10;
    wire top_tour1_c;
    wire RAM_DATA_1Z0Z_11;
    wire sTrigCounterZ0Z_0;
    wire RAM_DATA_1Z0Z_13;
    wire sTrigCounterZ0Z_1;
    wire RAM_DATA_1Z0Z_14;
    wire ADC2_c;
    wire RAM_DATA_1Z0Z_2;
    wire ADC6_c;
    wire RAM_DATA_1Z0Z_6;
    wire ADC0_c;
    wire RAM_DATA_1Z0Z_0;
    wire sDAC_mem_40Z0Z_3;
    wire sDAC_mem_40_1_sqmuxa;
    wire sDAC_mem_8_1_sqmuxa;
    wire N_317;
    wire sAddress_RNI6VH7_4Z0Z_1;
    wire sAddress_RNI70I7Z0Z_1;
    wire sAddress_RNIAM2A_0Z0Z_1;
    wire sDAC_data_2_32_ns_1_6_cascade_;
    wire sDAC_data_RNO_15Z0Z_6;
    wire sDAC_data_2_14_ns_1_6_cascade_;
    wire sDAC_data_RNO_10Z0Z_6;
    wire sDAC_data_RNO_2Z0Z_6;
    wire sDAC_data_2_41_ns_1_6_cascade_;
    wire sDAC_data_RNO_1Z0Z_6;
    wire sDAC_data_2_6_cascade_;
    wire sDAC_dataZ0Z_6;
    wire sDAC_mem_34Z0Z_5;
    wire sDAC_mem_2Z0Z_5;
    wire sDAC_mem_35Z0Z_5;
    wire sDAC_data_2_6_bm_1_8_cascade_;
    wire sDAC_mem_3Z0Z_5;
    wire sDAC_mem_42Z0Z_5;
    wire sDAC_mem_10Z0Z_5;
    wire sDAC_data_RNO_17Z0Z_8_cascade_;
    wire sDAC_mem_11Z0Z_5;
    wire sDAC_mem_40Z0Z_5;
    wire sDAC_mem_8Z0Z_5;
    wire sDAC_data_2_20_am_1_8_cascade_;
    wire sDAC_data_RNO_7Z0Z_8_cascade_;
    wire sDAC_data_RNO_8Z0Z_8;
    wire sDAC_data_RNO_15Z0Z_8;
    wire sDAC_data_2_14_ns_1_8_cascade_;
    wire sDAC_data_RNO_2Z0Z_8;
    wire sDAC_data_RNO_1Z0Z_8_cascade_;
    wire sDAC_data_2_8_cascade_;
    wire sDAC_data_2_32_ns_1_8_cascade_;
    wire sDAC_data_RNO_10Z0Z_8_cascade_;
    wire sDAC_data_2_41_ns_1_8;
    wire sDAC_mem_34Z0Z_1;
    wire sDAC_mem_2Z0Z_1;
    wire sDAC_mem_3Z0Z_1;
    wire sDAC_mem_35Z0Z_1;
    wire sDAC_data_2_6_bm_1_4_cascade_;
    wire sDAC_mem_42Z0Z_1;
    wire sDAC_mem_10Z0Z_1;
    wire sDAC_data_RNO_17Z0Z_4_cascade_;
    wire sDAC_mem_11Z0Z_1;
    wire sDAC_mem_40Z0Z_1;
    wire sDAC_mem_8Z0Z_1;
    wire sDAC_data_2_20_am_1_4_cascade_;
    wire sDAC_data_RNO_7Z0Z_4_cascade_;
    wire sDAC_data_RNO_8Z0Z_4;
    wire sDAC_mem_15Z0Z_0;
    wire sDAC_mem_14Z0Z_0;
    wire sDAC_data_RNO_18Z0Z_3_cascade_;
    wire sDAC_data_RNO_19Z0Z_3;
    wire sDAC_data_RNO_18Z0Z_4_cascade_;
    wire sDAC_data_2_24_ns_1_4;
    wire sDAC_mem_15Z0Z_1;
    wire sDAC_mem_14Z0Z_1;
    wire sDAC_data_RNO_19Z0Z_4;
    wire sDAC_mem_12Z0Z_0;
    wire sDAC_mem_12Z0Z_1;
    wire sDAC_mem_31Z0Z_5;
    wire sDAC_mem_30Z0Z_5;
    wire sDAC_mem_29Z0Z_5;
    wire sDAC_data_RNO_24Z0Z_8;
    wire sDAC_data_RNO_23Z0Z_8_cascade_;
    wire sDAC_data_RNO_11Z0Z_8;
    wire sDAC_mem_28Z0Z_5;
    wire sDAC_mem_24Z0Z_6;
    wire sDAC_data_RNO_30Z0Z_9_cascade_;
    wire sDAC_data_2_39_ns_1_9_cascade_;
    wire sDAC_mem_26Z0Z_6;
    wire sDAC_data_RNO_31Z0Z_9;
    wire sDAC_data_RNO_30Z0Z_7_cascade_;
    wire sDAC_data_2_39_ns_1_7_cascade_;
    wire sDAC_mem_26Z0Z_4;
    wire sDAC_data_RNO_31Z0Z_7;
    wire sDAC_mem_29Z0Z_4;
    wire sDAC_mem_28Z0Z_4;
    wire sDAC_data_RNO_23Z0Z_7;
    wire sDAC_mem_30Z0Z_4;
    wire sDAC_mem_31Z0Z_4;
    wire sDAC_data_RNO_24Z0Z_7;
    wire sDAC_mem_24Z0Z_4;
    wire sDAC_data_2_39_ns_1_8;
    wire sDAC_mem_26Z0Z_1;
    wire sDAC_data_RNO_30Z0Z_4_cascade_;
    wire sDAC_data_RNO_31Z0Z_4;
    wire sDAC_data_2_39_ns_1_4_cascade_;
    wire sDAC_mem_28Z0Z_1;
    wire sDAC_mem_29Z0Z_1;
    wire sDAC_data_RNO_23Z0Z_4;
    wire sDAC_mem_31Z0Z_1;
    wire sDAC_mem_30Z0Z_1;
    wire sDAC_data_RNO_24Z0Z_4;
    wire sDAC_mem_24Z0Z_1;
    wire sDAC_mem_24_1_sqmuxa;
    wire sDAC_data_RNO_31Z0Z_5;
    wire sDAC_mem_26Z0Z_2;
    wire sDAC_data_RNO_31Z0Z_8;
    wire sDAC_mem_26Z0Z_5;
    wire sDAC_mem_26_1_sqmuxa;
    wire \spi_master_inst.sclk_gen_u0.delay_clk_iZ0 ;
    wire \spi_master_inst.sclk_gen_u0.div_clk_iZ0 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i ;
    wire \spi_master_inst.sclk_gen_u0.falling_count_start_iZ0 ;
    wire \spi_master_inst.sclk_gen_u0.falling_count_start_i_i ;
    wire sCounter_i_0;
    wire bfn_13_14_0_;
    wire sCounter_i_1;
    wire un1_sacqtime_cry_0;
    wire sCounter_i_2;
    wire un1_sacqtime_cry_1;
    wire sCounter_i_3;
    wire un1_sacqtime_cry_2;
    wire sCounter_i_4;
    wire un1_sacqtime_cry_3;
    wire sCounter_i_5;
    wire un1_sacqtime_cry_4;
    wire sCounter_i_6;
    wire un1_sacqtime_cry_5;
    wire sCounter_i_7;
    wire un1_sacqtime_cry_6;
    wire un1_sacqtime_cry_7;
    wire sCounter_i_8;
    wire bfn_13_15_0_;
    wire sCounter_i_9;
    wire un1_sacqtime_cry_8;
    wire sCounter_i_10;
    wire un1_sacqtime_cry_9;
    wire sCounter_i_11;
    wire un1_sacqtime_cry_10;
    wire sCounter_i_12;
    wire un1_sacqtime_cry_11;
    wire sCounter_i_13;
    wire un1_sacqtime_cry_12;
    wire sCounter_i_14;
    wire un1_sacqtime_cry_13;
    wire sCounter_i_15;
    wire un1_sacqtime_cry_14;
    wire un1_sacqtime_cry_15;
    wire un1_sacqtime_cry_16_sf;
    wire bfn_13_16_0_;
    wire un1_sacqtime_cry_17_sf;
    wire un1_sacqtime_cry_16;
    wire un1_sacqtime_cry_18_sf;
    wire un1_sacqtime_cry_17;
    wire un1_sacqtime_cry_19_sf;
    wire un1_sacqtime_cry_18;
    wire un1_sacqtime_cry_20_sf;
    wire un1_sacqtime_cry_19;
    wire un1_sacqtime_cry_21_sf;
    wire un1_sacqtime_cry_20;
    wire un1_sacqtime_cry_22_sf;
    wire un1_sacqtime_cry_21;
    wire un1_sacqtime_cry_23_sf;
    wire un1_sacqtime_cry_22;
    wire un1_sacqtime_cry_23;
    wire bfn_13_17_0_;
    wire sADC_clk_prevZ0;
    wire N_71_cascade_;
    wire bfn_13_18_0_;
    wire sRAM_pointer_read_cry_0;
    wire sRAM_pointer_read_cry_1;
    wire sRAM_pointer_read_cry_2;
    wire sRAM_pointer_read_cry_3;
    wire sRAM_pointer_read_cry_4;
    wire sRAM_pointer_read_cry_5;
    wire sRAM_pointer_read_cry_6;
    wire sRAM_pointer_read_cry_7;
    wire bfn_13_19_0_;
    wire sRAM_pointer_read_cry_8;
    wire sRAM_pointer_read_cry_9;
    wire sRAM_pointer_read_cry_10;
    wire sRAM_pointer_read_cry_11;
    wire sRAM_pointer_read_cry_12;
    wire sRAM_pointer_read_cry_13;
    wire sRAM_pointer_read_cry_14;
    wire sRAM_pointer_read_cry_15;
    wire bfn_13_20_0_;
    wire sRAM_pointer_read_cry_16;
    wire sRAM_pointer_read_cry_17;
    wire N_28_g;
    wire sDAC_mem_36_1_sqmuxa;
    wire sDAC_data_RNO_29Z0Z_6;
    wire sDAC_mem_18Z0Z_3;
    wire sDAC_mem_18Z0Z_4;
    wire sDAC_data_RNO_29Z0Z_8;
    wire sDAC_mem_18Z0Z_5;
    wire sDAC_mem_18Z0Z_6;
    wire sDAC_mem_18_1_sqmuxa;
    wire sDAC_mem_15Z0Z_4;
    wire sDAC_mem_14Z0Z_4;
    wire sDAC_data_RNO_18Z0Z_7_cascade_;
    wire sDAC_data_RNO_19Z0Z_7;
    wire sDAC_data_RNO_18Z0Z_8_cascade_;
    wire sDAC_data_2_24_ns_1_8;
    wire sDAC_mem_15Z0Z_5;
    wire sDAC_mem_14Z0Z_5;
    wire sDAC_data_RNO_19Z0Z_8;
    wire sDAC_mem_12Z0Z_4;
    wire sDAC_mem_12Z0Z_5;
    wire sDAC_mem_38Z0Z_2;
    wire sDAC_mem_39Z0Z_2;
    wire sDAC_data_2_13_bm_1_5_cascade_;
    wire sDAC_mem_6Z0Z_2;
    wire sDAC_mem_38Z0Z_3;
    wire sDAC_mem_39Z0Z_3;
    wire sDAC_data_2_13_bm_1_6_cascade_;
    wire sDAC_data_RNO_5Z0Z_6;
    wire sDAC_mem_6Z0Z_3;
    wire sDAC_mem_38Z0Z_4;
    wire sDAC_mem_39Z0Z_4;
    wire sDAC_data_2_13_bm_1_7_cascade_;
    wire sDAC_data_RNO_28Z0Z_6;
    wire sDAC_mem_16Z0Z_3;
    wire sDAC_mem_16Z0Z_4;
    wire sDAC_data_RNO_28Z0Z_8;
    wire sDAC_mem_16Z0Z_5;
    wire sDAC_mem_16Z0Z_6;
    wire sDAC_data_RNO_10Z0Z_4_cascade_;
    wire sDAC_data_RNO_11Z0Z_4;
    wire sDAC_data_RNO_5Z0Z_4;
    wire sDAC_data_RNO_2Z0Z_4;
    wire sDAC_data_RNO_1Z0Z_4_cascade_;
    wire sDAC_data_2_41_ns_1_4;
    wire sDAC_data_2_4_cascade_;
    wire sDAC_data_RNO_15Z0Z_4;
    wire sDAC_data_2_14_ns_1_4;
    wire sDAC_data_2_32_ns_1_4;
    wire sDAC_mem_15Z0Z_2;
    wire sDAC_mem_14Z0Z_2;
    wire sDAC_data_RNO_18Z0Z_5_cascade_;
    wire sDAC_data_RNO_19Z0Z_5;
    wire sDAC_data_RNO_18Z0Z_6_cascade_;
    wire sDAC_data_2_24_ns_1_6;
    wire sDAC_mem_15Z0Z_3;
    wire sDAC_mem_14Z0Z_3;
    wire sDAC_data_RNO_19Z0Z_6;
    wire sDAC_mem_12Z0Z_2;
    wire sDAC_mem_12Z0Z_3;
    wire sEEACQZ0Z_0;
    wire sEEACQ_i_0;
    wire bfn_14_10_0_;
    wire sEEACQZ0Z_1;
    wire sEEACQ_i_1;
    wire un5_sdacdyn_cry_0;
    wire sEEACQZ0Z_2;
    wire sEEACQ_i_2;
    wire un5_sdacdyn_cry_1;
    wire sEEACQZ0Z_3;
    wire sEEACQ_i_3;
    wire un5_sdacdyn_cry_2;
    wire sEEACQZ0Z_4;
    wire sEEACQ_i_4;
    wire un5_sdacdyn_cry_3;
    wire sEEACQZ0Z_5;
    wire sEEACQ_i_5;
    wire un5_sdacdyn_cry_4;
    wire sEEACQZ0Z_6;
    wire sEEACQ_i_6;
    wire un5_sdacdyn_cry_5;
    wire sEEACQZ0Z_7;
    wire sEEACQ_i_7;
    wire un5_sdacdyn_cry_6;
    wire un5_sdacdyn_cry_7;
    wire sEEACQZ0Z_8;
    wire sEEACQ_i_8;
    wire bfn_14_11_0_;
    wire sEEACQZ0Z_9;
    wire sEEACQ_i_9;
    wire un5_sdacdyn_cry_8;
    wire sEEACQZ0Z_10;
    wire sEEACQ_i_10;
    wire un5_sdacdyn_cry_9;
    wire sEEACQZ0Z_11;
    wire sEEACQ_i_11;
    wire un5_sdacdyn_cry_10;
    wire sEEACQZ0Z_12;
    wire sEEACQ_i_12;
    wire un5_sdacdyn_cry_11;
    wire sEEACQZ0Z_13;
    wire sEEACQ_i_13;
    wire un5_sdacdyn_cry_12;
    wire sEEACQZ0Z_14;
    wire sEEACQ_i_14;
    wire un5_sdacdyn_cry_13;
    wire sEEACQZ0Z_15;
    wire sEEACQ_i_15;
    wire un5_sdacdyn_cry_14;
    wire un5_sdacdyn_cry_15;
    wire bfn_14_12_0_;
    wire un5_sdacdyn_cry_16;
    wire un5_sdacdyn_cry_17;
    wire un5_sdacdyn_cry_18;
    wire un5_sdacdyn_cry_19;
    wire un5_sdacdyn_cry_20;
    wire un5_sdacdyn_cry_21;
    wire un5_sdacdyn_cry_22;
    wire un5_sdacdyn_cry_23;
    wire N_106;
    wire bfn_14_13_0_;
    wire sDAC_mem_24Z0Z_7;
    wire sDAC_mem_26Z0Z_7;
    wire sDAC_dataZ0Z_10;
    wire sDAC_mem_24Z0Z_2;
    wire sDAC_data_RNO_30Z0Z_5;
    wire sDAC_mem_24Z0Z_5;
    wire sDAC_data_RNO_30Z0Z_8;
    wire sDAC_mem_29Z0Z_6;
    wire sDAC_data_RNO_23Z0Z_9;
    wire sDAC_mem_28Z0Z_6;
    wire sDAC_mem_31Z0Z_0;
    wire sDAC_mem_30Z0Z_0;
    wire sDAC_mem_31Z0Z_3;
    wire sDAC_mem_30Z0Z_3;
    wire sDAC_mem_31Z0Z_6;
    wire sDAC_mem_30Z0Z_6;
    wire sDAC_data_RNO_24Z0Z_9;
    wire sDAC_mem_16Z0Z_0;
    wire sDAC_mem_16Z0Z_1;
    wire sDAC_data_RNO_28Z0Z_4;
    wire sDAC_mem_16Z0Z_2;
    wire sDAC_mem_27Z0Z_1;
    wire sDAC_mem_27Z0Z_2;
    wire sDAC_mem_27Z0Z_4;
    wire sDAC_mem_27Z0Z_5;
    wire sDAC_mem_27Z0Z_6;
    wire sDAC_mem_27Z0Z_7;
    wire sDAC_mem_27_1_sqmuxa;
    wire sEEPonPoffZ0Z_0;
    wire un7_spon_0;
    wire sEEPonPoff_i_0;
    wire bfn_14_17_0_;
    wire un7_spon_1;
    wire sEEPonPoffZ0Z_1;
    wire sEEPonPoff_i_1;
    wire un4_spoff_cry_0;
    wire sEEPonPoffZ0Z_2;
    wire un7_spon_2;
    wire sEEPonPoff_i_2;
    wire un4_spoff_cry_1;
    wire sEEPonPoffZ0Z_3;
    wire un7_spon_3;
    wire sEEPonPoff_i_3;
    wire un4_spoff_cry_2;
    wire sEEPonPoffZ0Z_4;
    wire un7_spon_4;
    wire sEEPonPoff_i_4;
    wire un4_spoff_cry_3;
    wire sEEPonPoffZ0Z_5;
    wire un7_spon_5;
    wire sEEPonPoff_i_5;
    wire un4_spoff_cry_4;
    wire sEEPonPoffZ0Z_6;
    wire un7_spon_6;
    wire sEEPonPoff_i_6;
    wire un4_spoff_cry_5;
    wire un7_spon_7;
    wire sEEPonPoffZ0Z_7;
    wire sEEPonPoff_i_7;
    wire un4_spoff_cry_6;
    wire un4_spoff_cry_7;
    wire un7_spon_8;
    wire bfn_14_18_0_;
    wire un7_spon_9;
    wire un4_spoff_cry_8;
    wire un7_spon_10;
    wire un4_spoff_cry_9;
    wire un4_spoff_cry_10;
    wire un7_spon_12;
    wire un4_spoff_cry_11;
    wire un7_spon_13;
    wire un4_spoff_cry_12;
    wire un7_spon_14;
    wire un4_spoff_cry_13;
    wire un7_spon_15;
    wire un4_spoff_cry_14;
    wire un4_spoff_cry_15;
    wire un7_spon_16;
    wire bfn_14_19_0_;
    wire un7_spon_17;
    wire un4_spoff_cry_16;
    wire un7_spon_18;
    wire un4_spoff_cry_17;
    wire un4_spoff_cry_18;
    wire un4_spoff_cry_19;
    wire un4_spoff_cry_20;
    wire un7_spon_22;
    wire un4_spoff_cry_21;
    wire un7_spon_23;
    wire un4_spoff_cry_22;
    wire un4_spoff_cry_23;
    wire bfn_14_20_0_;
    wire un4_spoff_cry_23_THRU_CO;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_3 ;
    wire sDAC_dataZ0Z_4;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_4 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_7 ;
    wire sDAC_dataZ0Z_8;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_9 ;
    wire sEEDACZ0Z_1;
    wire sEEDACZ0Z_3;
    wire sEEDACZ0Z_5;
    wire sEEDACZ0Z_7;
    wire sEEDAC_1_sqmuxa;
    wire sDAC_data_RNO_29Z0Z_7;
    wire sDAC_data_RNO_28Z0Z_7;
    wire sDAC_data_2_32_ns_1_7;
    wire sDAC_data_2_14_ns_1_7_cascade_;
    wire sDAC_data_RNO_5Z0Z_7;
    wire sDAC_data_RNO_11Z0Z_7;
    wire sDAC_data_RNO_10Z0Z_7;
    wire sDAC_data_2_41_ns_1_7_cascade_;
    wire sDAC_data_RNO_1Z0Z_7;
    wire sEEDACZ0Z_4;
    wire sDAC_data_2_7_cascade_;
    wire sDAC_dataZ0Z_7;
    wire sDAC_data_RNO_1Z0Z_9_cascade_;
    wire sEEDACZ0Z_6;
    wire sDAC_data_2_9_cascade_;
    wire sDAC_dataZ0Z_9;
    wire sDAC_data_2_14_ns_1_9;
    wire sDAC_data_RNO_29Z0Z_9;
    wire sDAC_data_RNO_28Z0Z_9;
    wire sDAC_data_2_32_ns_1_9_cascade_;
    wire sDAC_data_RNO_10Z0Z_9_cascade_;
    wire sDAC_data_RNO_11Z0Z_9;
    wire sDAC_data_2_41_ns_1_9;
    wire sDAC_data_RNO_20Z0Z_8;
    wire sDAC_mem_20Z0Z_5;
    wire sDAC_data_RNO_20Z0Z_9;
    wire sDAC_mem_20Z0Z_6;
    wire sDAC_mem_22Z0Z_0;
    wire sDAC_mem_22Z0Z_1;
    wire sDAC_data_RNO_21Z0Z_4;
    wire sDAC_mem_22Z0Z_2;
    wire sDAC_mem_22Z0Z_3;
    wire sDAC_data_RNO_21Z0Z_6;
    wire sDAC_mem_36Z0Z_4;
    wire sDAC_data_2_13_am_1_7_cascade_;
    wire sDAC_data_RNO_4Z0Z_7;
    wire sDAC_mem_4Z0Z_4;
    wire sDAC_mem_36Z0Z_5;
    wire sDAC_data_2_13_am_1_8_cascade_;
    wire sDAC_data_RNO_4Z0Z_8;
    wire sDAC_mem_38Z0Z_5;
    wire sDAC_mem_39Z0Z_5;
    wire sDAC_data_2_13_bm_1_8_cascade_;
    wire sDAC_mem_7Z0Z_5;
    wire sDAC_data_RNO_5Z0Z_8;
    wire sDAC_mem_6Z0Z_5;
    wire sDAC_mem_38Z0Z_6;
    wire sDAC_data_2_13_bm_1_9_cascade_;
    wire sDAC_mem_39Z0Z_6;
    wire sDAC_data_RNO_5Z0Z_9;
    wire sDAC_mem_6Z0Z_6;
    wire sDAC_mem_40Z0Z_7;
    wire sDAC_mem_8Z0Z_7;
    wire sDAC_data_2_20_am_1_10_cascade_;
    wire sDAC_mem_36Z0Z_6;
    wire sDAC_data_2_13_am_1_9_cascade_;
    wire sDAC_data_RNO_4Z0Z_9;
    wire sDAC_mem_4Z0Z_6;
    wire sDAC_mem_38Z0Z_7;
    wire sDAC_mem_39Z0Z_7;
    wire sDAC_data_2_13_bm_1_10_cascade_;
    wire sDAC_mem_7Z0Z_7;
    wire sDAC_mem_38Z0Z_0;
    wire sDAC_mem_39Z0Z_0;
    wire sDAC_data_2_13_bm_1_3_cascade_;
    wire sDAC_mem_7Z0Z_0;
    wire sDAC_mem_38Z0Z_1;
    wire sDAC_data_2_13_bm_1_4;
    wire sDAC_mem_34Z0Z_7;
    wire sDAC_mem_2Z0Z_7;
    wire sDAC_mem_2_1_sqmuxa;
    wire sDAC_mem_12Z0Z_7;
    wire sDAC_data_RNO_18Z0Z_10_cascade_;
    wire sDAC_mem_15Z0Z_7;
    wire sDAC_mem_14Z0Z_7;
    wire sDAC_data_RNO_19Z0Z_10;
    wire sDAC_mem_42Z0Z_7;
    wire sDAC_mem_10Z0Z_7;
    wire sDAC_data_RNO_17Z0Z_10_cascade_;
    wire sDAC_mem_11Z0Z_7;
    wire sDAC_data_2_24_ns_1_10;
    wire sDAC_data_RNO_8Z0Z_10_cascade_;
    wire sDAC_data_RNO_7Z0Z_10;
    wire un7_spon_20;
    wire un7_spon_19;
    wire un7_spon_21;
    wire un7_spon_11;
    wire g0_12;
    wire sDAC_data_RNO_2Z0Z_10;
    wire sDAC_data_2_41_ns_1_10_cascade_;
    wire sDAC_data_2_10;
    wire sbuttonModeStatus_0_sqmuxa_17;
    wire sDAC_mem_22Z0Z_7;
    wire sDAC_data_RNO_28Z0Z_10_cascade_;
    wire sDAC_data_RNO_21Z0Z_10;
    wire sDAC_data_2_32_ns_1_10_cascade_;
    wire sDAC_data_RNO_10Z0Z_10;
    wire sDAC_data_RNO_20Z0Z_10;
    wire sDAC_mem_18Z0Z_7;
    wire sDAC_data_RNO_29Z0Z_10;
    wire sDAC_mem_16Z0Z_7;
    wire sDAC_mem_16_1_sqmuxa;
    wire sDAC_data_RNO_31Z0Z_10;
    wire sDAC_data_RNO_30Z0Z_10;
    wire sDAC_mem_31Z0Z_7;
    wire sDAC_mem_30Z0Z_7;
    wire sDAC_mem_29Z0Z_7;
    wire sDAC_data_RNO_24Z0Z_10;
    wire sDAC_data_RNO_23Z0Z_10_cascade_;
    wire sDAC_data_2_39_ns_1_10;
    wire sDAC_data_RNO_11Z0Z_10;
    wire sDAC_mem_28Z0Z_7;
    wire sDAC_mem_27Z0Z_0;
    wire sDAC_mem_26Z0Z_0;
    wire sDAC_mem_24Z0Z_0;
    wire sDAC_data_RNO_30Z0Z_3_cascade_;
    wire sDAC_data_RNO_31Z0Z_3;
    wire sDAC_data_RNO_24Z0Z_3;
    wire sDAC_data_2_39_ns_1_3_cascade_;
    wire sDAC_data_RNO_21Z0Z_7;
    wire sDAC_mem_22Z0Z_4;
    wire sDAC_data_RNO_21Z0Z_8;
    wire sDAC_mem_22Z0Z_5;
    wire sDAC_data_RNO_21Z0Z_9;
    wire sDAC_mem_22Z0Z_6;
    wire sDAC_mem_22_1_sqmuxa;
    wire sDAC_mem_29Z0Z_0;
    wire sDAC_mem_28Z0Z_0;
    wire sDAC_data_RNO_23Z0Z_3;
    wire sDAC_mem_29Z0Z_3;
    wire sDAC_mem_28Z0Z_3;
    wire sbuttonModeStatus_0_sqmuxa_14_cascade_;
    wire sbuttonModeStatus_0_sqmuxa_13;
    wire sbuttonModeStatus_0_sqmuxa_22;
    wire sEEPonPoff_1_sqmuxa_0_a3_0_a2_1;
    wire sPointer_RNI5LBD1Z0Z_0;
    wire sEEPonPoff_1_sqmuxa;
    wire RAM_nWE_0_i;
    wire sRead_data_RNOZ0Z_0_cascade_;
    wire ADC_clk_c;
    wire sRead_dataZ0;
    wire spi_data_miso_0_sqmuxa_2_i_o2_4;
    wire spi_data_miso_0_sqmuxa_2_i_o2_5;
    wire ADC3_c;
    wire RAM_DATA_1Z0Z_3;
    wire sDAC_mem_19Z0Z_4;
    wire sDAC_mem_19Z0Z_5;
    wire sDAC_mem_19Z0Z_6;
    wire sDAC_mem_19Z0Z_7;
    wire sDAC_mem_21Z0Z_5;
    wire sDAC_mem_21Z0Z_6;
    wire sDAC_mem_21Z0Z_7;
    wire sDAC_mem_21_1_sqmuxa;
    wire sDAC_mem_34Z0Z_4;
    wire sDAC_mem_2Z0Z_4;
    wire sDAC_mem_35Z0Z_4;
    wire sDAC_data_2_6_bm_1_7_cascade_;
    wire sDAC_mem_3Z0Z_4;
    wire sDAC_data_RNO_15Z0Z_7;
    wire sDAC_mem_40Z0Z_4;
    wire sDAC_mem_8Z0Z_4;
    wire sDAC_data_2_20_am_1_7_cascade_;
    wire sDAC_data_2_24_ns_1_7;
    wire sDAC_data_RNO_7Z0Z_7_cascade_;
    wire sDAC_data_RNO_2Z0Z_7;
    wire sDAC_mem_11Z0Z_4;
    wire sDAC_data_RNO_8Z0Z_7;
    wire sDAC_mem_42Z0Z_4;
    wire sDAC_mem_10Z0Z_4;
    wire sDAC_data_RNO_17Z0Z_7;
    wire sDAC_mem_34Z0Z_6;
    wire sDAC_mem_2Z0Z_6;
    wire sDAC_mem_35Z0Z_6;
    wire sDAC_data_2_6_bm_1_9_cascade_;
    wire sDAC_mem_3Z0Z_6;
    wire sDAC_data_RNO_15Z0Z_9;
    wire sDAC_mem_42Z0Z_6;
    wire sDAC_mem_10Z0Z_6;
    wire sDAC_data_RNO_17Z0Z_9_cascade_;
    wire sDAC_mem_11Z0Z_6;
    wire sDAC_mem_40Z0Z_6;
    wire sDAC_mem_8Z0Z_6;
    wire sDAC_data_2_20_am_1_9_cascade_;
    wire sDAC_data_RNO_7Z0Z_9_cascade_;
    wire sDAC_data_RNO_8Z0Z_9;
    wire sDAC_data_RNO_2Z0Z_9;
    wire sDAC_data_RNO_26Z0Z_9_cascade_;
    wire sDAC_mem_32Z0Z_6;
    wire sDAC_data_RNO_14Z0Z_9;
    wire sDAC_mem_21Z0Z_0;
    wire sDAC_mem_21Z0Z_1;
    wire sDAC_data_RNO_20Z0Z_4;
    wire sDAC_mem_21Z0Z_2;
    wire sDAC_mem_21Z0Z_3;
    wire sDAC_data_RNO_20Z0Z_6;
    wire sDAC_mem_21Z0Z_4;
    wire sDAC_data_RNO_20Z0Z_7;
    wire bfn_16_8_0_;
    wire sDAC_mem_pointer_0_cry_1;
    wire sDAC_mem_pointer_0_cry_2;
    wire sDAC_mem_pointer_0_cry_3;
    wire sDAC_mem_pointer_0_cry_4;
    wire sDAC_mem_34Z0Z_2;
    wire sDAC_mem_2Z0Z_2;
    wire sDAC_mem_35Z0Z_2;
    wire sDAC_data_2_6_bm_1_5_cascade_;
    wire sDAC_mem_3Z0Z_2;
    wire sDAC_mem_42Z0Z_2;
    wire sDAC_mem_10Z0Z_2;
    wire sDAC_data_RNO_17Z0Z_5_cascade_;
    wire sDAC_mem_11Z0Z_2;
    wire sDAC_mem_40Z0Z_2;
    wire sDAC_mem_8Z0Z_2;
    wire sDAC_data_2_20_am_1_5_cascade_;
    wire sDAC_data_2_24_ns_1_5;
    wire sDAC_data_RNO_7Z0Z_5_cascade_;
    wire sDAC_data_RNO_8Z0Z_5;
    wire sDAC_mem_34Z0Z_0;
    wire sDAC_mem_2Z0Z_0;
    wire sDAC_mem_35Z0Z_0;
    wire sDAC_data_2_6_bm_1_3_cascade_;
    wire sDAC_mem_3Z0Z_0;
    wire sDAC_mem_42Z0Z_0;
    wire sDAC_mem_10Z0Z_0;
    wire sDAC_data_RNO_17Z0Z_3_cascade_;
    wire sDAC_mem_11Z0Z_0;
    wire sDAC_mem_40Z0Z_0;
    wire sDAC_mem_8Z0Z_0;
    wire sDAC_data_2_20_am_1_3_cascade_;
    wire sDAC_data_2_24_ns_1_3;
    wire sDAC_data_RNO_7Z0Z_3_cascade_;
    wire sDAC_data_RNO_8Z0Z_3;
    wire N_333;
    wire sDAC_mem_19Z0Z_0;
    wire sDAC_mem_18Z0Z_0;
    wire sDAC_mem_19Z0Z_1;
    wire sDAC_mem_18Z0Z_1;
    wire sDAC_data_RNO_29Z0Z_4;
    wire sDAC_mem_19Z0Z_2;
    wire sDAC_mem_18Z0Z_2;
    wire sDAC_mem_19Z0Z_3;
    wire sDAC_mem_19_1_sqmuxa;
    wire sDAC_mem_35Z0Z_7;
    wire sDAC_data_2_6_bm_1_10;
    wire sDAC_data_RNO_15Z0Z_10_cascade_;
    wire sDAC_data_RNO_5Z0Z_10;
    wire sDAC_data_2_14_ns_1_10_cascade_;
    wire sDAC_data_RNO_1Z0Z_10;
    wire sDAC_mem_36Z0Z_7;
    wire sDAC_data_2_13_am_1_10_cascade_;
    wire sDAC_data_RNO_4Z0Z_10;
    wire sDAC_data_RNO_26Z0Z_10;
    wire sDAC_data_RNO_14Z0Z_10;
    wire bfn_16_13_0_;
    wire button_debounce_counterZ0Z_2;
    wire un1_button_debounce_counter_cry_1;
    wire button_debounce_counterZ0Z_3;
    wire un1_button_debounce_counter_cry_2;
    wire button_debounce_counterZ0Z_4;
    wire un1_button_debounce_counter_cry_3;
    wire button_debounce_counterZ0Z_5;
    wire un1_button_debounce_counter_cry_4;
    wire button_debounce_counterZ0Z_6;
    wire un1_button_debounce_counter_cry_5;
    wire un1_button_debounce_counter_cry_6;
    wire un1_button_debounce_counter_cry_7;
    wire un1_button_debounce_counter_cry_8;
    wire bfn_16_14_0_;
    wire un1_button_debounce_counter_cry_9;
    wire un1_button_debounce_counter_cry_10;
    wire un1_button_debounce_counter_cry_11;
    wire un1_button_debounce_counter_cry_12;
    wire un1_button_debounce_counter_cry_13;
    wire button_debounce_counterZ0Z_15;
    wire un1_button_debounce_counter_cry_14;
    wire button_debounce_counterZ0Z_16;
    wire un1_button_debounce_counter_cry_15;
    wire un1_button_debounce_counter_cry_16;
    wire button_debounce_counterZ0Z_17;
    wire bfn_16_15_0_;
    wire button_debounce_counterZ0Z_18;
    wire un1_button_debounce_counter_cry_17;
    wire button_debounce_counterZ0Z_19;
    wire un1_button_debounce_counter_cry_18;
    wire button_debounce_counterZ0Z_20;
    wire un1_button_debounce_counter_cry_19;
    wire button_debounce_counterZ0Z_21;
    wire un1_button_debounce_counter_cry_20;
    wire button_debounce_counterZ0Z_22;
    wire un1_button_debounce_counter_cry_21;
    wire un1_button_debounce_counter_cry_22;
    wire un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO;
    wire un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO;
    wire bfn_16_16_0_;
    wire button_debounce_counterZ0Z_23;
    wire LED3_c_0;
    wire sRAM_pointer_readZ0Z_5;
    wire sRAM_pointer_writeZ0Z_5;
    wire RAM_ADD_c_5;
    wire sRAM_pointer_readZ0Z_0;
    wire sRAM_pointer_writeZ0Z_0;
    wire RAM_ADD_c_0;
    wire sRAM_pointer_readZ0Z_10;
    wire sRAM_pointer_writeZ0Z_10;
    wire RAM_ADD_c_10;
    wire sRAM_pointer_readZ0Z_11;
    wire sRAM_pointer_writeZ0Z_11;
    wire RAM_ADD_c_11;
    wire sRAM_pointer_writeZ0Z_12;
    wire sRAM_pointer_readZ0Z_12;
    wire RAM_ADD_c_12;
    wire sRAM_pointer_readZ0Z_13;
    wire sRAM_pointer_writeZ0Z_13;
    wire RAM_ADD_c_13;
    wire sRAM_pointer_writeZ0Z_14;
    wire sRAM_pointer_readZ0Z_14;
    wire RAM_ADD_c_14;
    wire sRAM_pointer_readZ0Z_15;
    wire sRAM_pointer_writeZ0Z_15;
    wire RAM_ADD_c_15;
    wire sRAM_pointer_readZ0Z_16;
    wire sRAM_pointer_writeZ0Z_16;
    wire RAM_ADD_c_16;
    wire sRAM_pointer_writeZ0Z_17;
    wire sRAM_pointer_readZ0Z_17;
    wire RAM_ADD_c_17;
    wire sRAM_pointer_writeZ0Z_18;
    wire sRAM_pointer_readZ0Z_18;
    wire RAM_ADD_c_18;
    wire sRAM_pointer_writeZ0Z_9;
    wire sRAM_pointer_readZ0Z_9;
    wire RAM_ADD_c_9;
    wire sRAM_pointer_writeZ0Z_7;
    wire sRAM_pointer_readZ0Z_7;
    wire RAM_ADD_c_7;
    wire sRAM_pointer_readZ0Z_2;
    wire sRAM_pointer_writeZ0Z_2;
    wire RAM_ADD_c_2;
    wire sRAM_pointer_writeZ0Z_1;
    wire sRAM_pointer_readZ0Z_1;
    wire RAM_ADD_c_1;
    wire sRAM_pointer_writeZ0Z_6;
    wire sRAM_pointer_readZ0Z_6;
    wire RAM_ADD_c_6;
    wire ADC4_c;
    wire RAM_DATA_1Z0Z_4;
    wire sDAC_mem_4Z0Z_5;
    wire sDAC_mem_4Z0Z_7;
    wire sDAC_mem_20Z0Z_0;
    wire sDAC_mem_20Z0Z_1;
    wire sDAC_mem_20Z0Z_2;
    wire sDAC_mem_20Z0Z_3;
    wire sDAC_mem_20Z0Z_4;
    wire sDAC_mem_20Z0Z_7;
    wire sDAC_mem_20_1_sqmuxa;
    wire sDAC_mem_6Z0Z_0;
    wire sDAC_mem_6Z0Z_1;
    wire sDAC_mem_6Z0Z_4;
    wire sDAC_mem_6Z0Z_7;
    wire sDAC_mem_6_1_sqmuxa;
    wire sDAC_mem_23Z0Z_0;
    wire sDAC_mem_23Z0Z_1;
    wire sDAC_mem_23Z0Z_2;
    wire sDAC_mem_23Z0Z_3;
    wire sDAC_mem_23Z0Z_4;
    wire sDAC_mem_23Z0Z_5;
    wire sDAC_mem_23Z0Z_6;
    wire sDAC_mem_23Z0Z_7;
    wire sDAC_mem_23_1_sqmuxa;
    wire sDAC_data_RNO_26Z0Z_6_cascade_;
    wire sDAC_mem_32Z0Z_3;
    wire sDAC_data_RNO_14Z0Z_6;
    wire sDAC_data_RNO_26Z0Z_7_cascade_;
    wire sDAC_data_RNO_14Z0Z_7;
    wire sDAC_mem_32Z0Z_4;
    wire sDAC_data_RNO_26Z0Z_8_cascade_;
    wire sDAC_data_RNO_14Z0Z_8;
    wire sDAC_mem_9Z0Z_0;
    wire sDAC_mem_9Z0Z_1;
    wire sDAC_mem_9Z0Z_2;
    wire sDAC_mem_9Z0Z_3;
    wire sDAC_mem_9Z0Z_4;
    wire sDAC_mem_9Z0Z_5;
    wire sDAC_mem_9Z0Z_6;
    wire sDAC_mem_9Z0Z_7;
    wire sDAC_mem_15Z0Z_6;
    wire sDAC_mem_14Z0Z_6;
    wire sDAC_data_RNO_18Z0Z_9_cascade_;
    wire sDAC_data_RNO_19Z0Z_9;
    wire sDAC_data_2_24_ns_1_9;
    wire sDAC_mem_12Z0Z_6;
    wire sDAC_mem_12_1_sqmuxa;
    wire op_le_op_le_un15_sdacdynlt4_cascade_;
    wire un17_sdacdyn_1;
    wire sDAC_mem_pointerZ0Z_7;
    wire sDAC_mem_pointerZ0Z_6;
    wire un17_sdacdyn_0;
    wire sDAC_data_RNO_5Z0Z_5;
    wire sDAC_data_RNO_2Z0Z_5;
    wire sDAC_data_RNO_1Z0Z_5_cascade_;
    wire sEEDACZ0Z_2;
    wire sDAC_data_2_5_cascade_;
    wire sDAC_dataZ0Z_5;
    wire sDAC_data_RNO_15Z0Z_5;
    wire sDAC_data_2_14_ns_1_5;
    wire sDAC_data_RNO_29Z0Z_5;
    wire sDAC_data_RNO_28Z0Z_5;
    wire sDAC_data_RNO_20Z0Z_5;
    wire sDAC_data_2_32_ns_1_5_cascade_;
    wire sDAC_data_RNO_21Z0Z_5;
    wire sDAC_data_RNO_10Z0Z_5_cascade_;
    wire sDAC_data_2_41_ns_1_5;
    wire sDAC_data_RNO_5Z0Z_3;
    wire sDAC_data_RNO_2Z0Z_3;
    wire sDAC_data_RNO_1Z0Z_3_cascade_;
    wire sEEDACZ0Z_0;
    wire sDAC_data_2_3_cascade_;
    wire un5_sdacdyn_cry_23_c_RNIELGZ0Z28;
    wire sDAC_dataZ0Z_3;
    wire sDAC_data_RNO_21Z0Z_3;
    wire sDAC_data_RNO_20Z0Z_3;
    wire sDAC_mem_pointerZ0Z_4;
    wire sDAC_mem_pointerZ0Z_3;
    wire sDAC_data_RNO_10Z0Z_3_cascade_;
    wire sDAC_data_RNO_11Z0Z_3;
    wire sDAC_data_2_41_ns_1_3;
    wire sDAC_data_RNO_15Z0Z_3;
    wire sDAC_data_2_14_ns_1_3;
    wire sDAC_data_RNO_28Z0Z_3;
    wire sDAC_data_RNO_29Z0Z_3;
    wire sDAC_data_2_32_ns_1_3;
    wire sDAC_data_2_39_ns_1_5;
    wire sDAC_data_RNO_11Z0Z_5;
    wire sDAC_mem_29Z0Z_2;
    wire sDAC_data_RNO_23Z0Z_5;
    wire sDAC_mem_24Z0Z_3;
    wire sDAC_mem_pointerZ0Z_1;
    wire sDAC_data_RNO_30Z0Z_6_cascade_;
    wire sDAC_mem_pointerZ0Z_2;
    wire sDAC_data_RNO_24Z0Z_6;
    wire sDAC_data_2_39_ns_1_6_cascade_;
    wire sDAC_data_RNO_23Z0Z_6;
    wire sDAC_data_RNO_11Z0Z_6;
    wire sDAC_mem_28Z0Z_2;
    wire sDAC_mem_28_1_sqmuxa;
    wire sDAC_mem_30Z0Z_2;
    wire sDAC_mem_31Z0Z_2;
    wire sDAC_data_RNO_24Z0Z_5;
    wire sDAC_mem_26Z0Z_3;
    wire sDAC_mem_27Z0Z_3;
    wire sDAC_data_RNO_31Z0Z_6;
    wire bfn_17_13_0_;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0 ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1 ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2 ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3 ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4 ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5 ;
    wire sDAC_mem_17Z0Z_0;
    wire sDAC_mem_17Z0Z_1;
    wire sDAC_mem_17Z0Z_2;
    wire sDAC_mem_17Z0Z_3;
    wire sDAC_mem_17Z0Z_4;
    wire sDAC_mem_17Z0Z_5;
    wire sDAC_mem_17Z0Z_6;
    wire sDAC_mem_17Z0Z_7;
    wire RAM_DATA_in_14;
    wire RAM_DATA_in_6;
    wire button_debounce_counterZ0Z_13;
    wire button_debounce_counterZ0Z_12;
    wire button_debounce_counterZ0Z_14;
    wire button_debounce_counterZ0Z_11;
    wire sbuttonModeStatus_0_sqmuxa_15;
    wire button_debounce_counterZ0Z_9;
    wire button_debounce_counterZ0Z_7;
    wire button_debounce_counterZ0Z_10;
    wire button_debounce_counterZ0Z_8;
    wire sbuttonModeStatus_0_sqmuxa_16;
    wire RAM_DATA_in_0;
    wire RAM_DATA_in_8;
    wire RAM_DATA_in_12;
    wire RAM_DATA_in_4;
    wire sEEPointerResetZ0;
    wire un4_sacqtime_cry_23_c_RNITTSZ0Z3_cascade_;
    wire N_28;
    wire sSPI_MSB0LSBZ0Z1;
    wire spi_mosi_ready_prev3_RNILKERZ0;
    wire RAM_DATA_cl_11Z0Z_15;
    wire RAM_DATA_cl_12Z0Z_15;
    wire sCounterRAMZ0Z_0;
    wire bfn_17_18_0_;
    wire sCounterRAMZ0Z_1;
    wire sCounterRAM_cry_0;
    wire sCounterRAMZ0Z_2;
    wire sCounterRAM_cry_1;
    wire sCounterRAMZ0Z_3;
    wire sCounterRAM_cry_2;
    wire sCounterRAMZ0Z_4;
    wire sCounterRAM_cry_3;
    wire sCounterRAMZ0Z_5;
    wire sCounterRAM_cry_4;
    wire sCounterRAMZ0Z_6;
    wire sCounterRAM_cry_5;
    wire N_70_i;
    wire sCounterRAM_cry_6;
    wire sCounterRAMZ0Z_7;
    wire RAM_DATA_cl_6Z0Z_15;
    wire RAM_DATA_cl_7Z0Z_15;
    wire RAM_DATA_cl_8Z0Z_15;
    wire RAM_DATA_cl_9Z0Z_15;
    wire RAM_DATA_clZ0Z_15;
    wire RAM_DATA_1Z0Z_7;
    wire sDAC_mem_41Z0Z_4;
    wire sDAC_mem_36Z0Z_3;
    wire sDAC_mem_4Z0Z_3;
    wire sDAC_data_2_13_am_1_6_cascade_;
    wire sDAC_data_RNO_4Z0Z_6;
    wire sDAC_mem_32Z0Z_5;
    wire sDAC_mem_32Z0Z_7;
    wire sDAC_mem_41Z0Z_0;
    wire sDAC_mem_41Z0Z_1;
    wire sDAC_mem_41Z0Z_2;
    wire sDAC_mem_41Z0Z_3;
    wire sDAC_mem_41Z0Z_5;
    wire sDAC_mem_41Z0Z_6;
    wire sDAC_mem_41Z0Z_7;
    wire sDAC_mem_9_1_sqmuxa;
    wire sDAC_mem_41_1_sqmuxa;
    wire sAddress_RNI6VH7_6Z0Z_1;
    wire sAddress_RNI6VH7_6Z0Z_1_cascade_;
    wire sAddressZ0Z_5;
    wire sAddress_RNIP2UK1Z0Z_4;
    wire sAddressZ0Z_2;
    wire sAddressZ0Z_1;
    wire sAddressZ0Z_3;
    wire sAddressZ0Z_0;
    wire sAddress_RNIAM2A_1Z0Z_1;
    wire sAddress_RNIAM2A_1Z0Z_1_cascade_;
    wire sAddress_RNIVREN1Z0Z_4;
    wire sDAC_mem_17_1_sqmuxa;
    wire sDAC_mem_37Z0Z_3;
    wire sDAC_mem_37Z0Z_4;
    wire sDAC_mem_37Z0Z_5;
    wire sDAC_mem_37Z0Z_6;
    wire sDAC_mem_37Z0Z_7;
    wire sDAC_mem_37_1_sqmuxa;
    wire sDAC_data_RNO_26Z0Z_3;
    wire sDAC_data_RNO_14Z0Z_3;
    wire sDAC_data_RNO_26Z0Z_4_cascade_;
    wire sDAC_data_RNO_14Z0Z_4;
    wire sDAC_mem_32Z0Z_0;
    wire sDAC_mem_32Z0Z_1;
    wire sDAC_data_RNO_26Z0Z_5_cascade_;
    wire sDAC_data_RNO_14Z0Z_5;
    wire sDAC_mem_32Z0Z_2;
    wire sDAC_mem_32_1_sqmuxa;
    wire sDAC_mem_36Z0Z_0;
    wire sDAC_mem_37Z0Z_0;
    wire sDAC_data_2_13_am_1_3_cascade_;
    wire sDAC_data_RNO_4Z0Z_3;
    wire sDAC_mem_4Z0Z_0;
    wire sDAC_mem_36Z0Z_1;
    wire sDAC_data_2_13_am_1_4_cascade_;
    wire sDAC_mem_37Z0Z_1;
    wire sDAC_data_RNO_4Z0Z_4;
    wire sDAC_mem_4Z0Z_1;
    wire sDAC_mem_4_1_sqmuxa;
    wire sDAC_mem_pointerZ0Z_5;
    wire sDAC_mem_36Z0Z_2;
    wire sDAC_mem_4Z0Z_2;
    wire sDAC_mem_pointerZ0Z_0;
    wire sDAC_mem_37Z0Z_2;
    wire sDAC_data_2_13_am_1_5_cascade_;
    wire sDAC_data_RNO_4Z0Z_5;
    wire sDAC_mem_25Z0Z_5;
    wire sDAC_mem_25Z0Z_2;
    wire sDAC_mem_25Z0Z_3;
    wire sDAC_mem_25Z0Z_4;
    wire sDAC_mem_25Z0Z_0;
    wire sDAC_mem_25Z0Z_6;
    wire sDAC_mem_25Z0Z_7;
    wire \spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0 ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1 ;
    wire \spi_slave_inst.un23_i_ssn ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2 ;
    wire spi_data_misoZ0Z_0;
    wire spi_data_misoZ0Z_4;
    wire spi_data_misoZ0Z_6;
    wire \spi_slave_inst.un4_i_wr ;
    wire bfn_18_15_0_;
    wire sCounterADC_cry_0;
    wire sCounterADC_cry_1;
    wire sCounterADC_cry_2;
    wire sCounterADCZ0Z_4;
    wire sCounterADC_cry_3;
    wire sCounterADCZ0Z_5;
    wire sCounterADC_cry_4;
    wire sCounterADC_cry_5;
    wire sCounterADC_cry_6;
    wire RAM_DATA_in_5;
    wire RAM_DATA_in_13;
    wire spi_data_misoZ0Z_5;
    wire RAM_DATA_in_15;
    wire RAM_DATA_in_7;
    wire spi_data_misoZ0Z_7;
    wire RAM_DATA_in_3;
    wire RAM_DATA_in_11;
    wire spi_data_misoZ0Z_3;
    wire RAM_DATA_in_10;
    wire RAM_DATA_in_2;
    wire spi_data_misoZ0Z_2;
    wire RAM_DATA_in_1;
    wire RAM_DATA_in_9;
    wire N_75;
    wire spi_data_misoZ0Z_1;
    wire sSPI_MSB0LSB1_RNIGRPGZ0Z4;
    wire sRAM_pointer_writeZ0Z_8;
    wire sRAM_pointer_readZ0Z_8;
    wire RAM_ADD_c_8;
    wire sRAM_pointer_writeZ0Z_4;
    wire sRAM_pointer_readZ0Z_4;
    wire RAM_ADD_c_4;
    wire sRAM_pointer_writeZ0Z_3;
    wire un1_sacqtime_cry_23_THRU_CO;
    wire sRAM_pointer_readZ0Z_3;
    wire un4_sacqtime_cry_23_THRU_CO;
    wire RAM_ADD_c_3;
    wire N_67_i;
    wire RAM_DATA_cl_13Z0Z_15;
    wire RAM_DATA_cl_14Z0Z_15;
    wire RAM_DATA_cl_15Z0Z_15;
    wire RAM_DATA_cl_1Z0Z_15;
    wire RAM_DATA_cl_10Z0Z_15;
    wire RAM_DATA_cl_3Z0Z_15;
    wire RAM_DATA_cl_4Z0Z_15;
    wire RAM_DATA_cl_2Z0Z_15;
    wire GNDG0;
    wire op_eq_scounterdac10_g;
    wire sDAC_dataZ0Z_2;
    wire \spi_master_inst.spi_data_path_u1.tx_ready_iZ0 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_2 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2 ;
    wire sDAC_mem_7Z0Z_2;
    wire sDAC_mem_7Z0Z_3;
    wire sDAC_mem_7Z0Z_4;
    wire sDAC_mem_7Z0Z_6;
    wire sDAC_mem_7_1_sqmuxa;
    wire sDAC_mem_3Z0Z_7;
    wire sDAC_mem_3_1_sqmuxa;
    wire sDAC_mem_1Z0Z_0;
    wire sDAC_mem_1Z0Z_1;
    wire sDAC_mem_1Z0Z_2;
    wire sDAC_mem_1Z0Z_3;
    wire sDAC_mem_1Z0Z_4;
    wire sDAC_mem_1Z0Z_5;
    wire sDAC_mem_1Z0Z_6;
    wire sDAC_mem_1Z0Z_7;
    wire sDAC_mem_1_1_sqmuxa;
    wire sDAC_mem_33Z0Z_0;
    wire sDAC_mem_33Z0Z_1;
    wire sDAC_mem_33Z0Z_2;
    wire sDAC_mem_33Z0Z_3;
    wire sDAC_mem_33Z0Z_4;
    wire sDAC_mem_33Z0Z_5;
    wire sDAC_mem_33Z0Z_6;
    wire sDAC_mem_33Z0Z_7;
    wire sDAC_mem_33_1_sqmuxa;
    wire sDAC_mem_5Z0Z_0;
    wire sDAC_mem_5Z0Z_1;
    wire sDAC_mem_5Z0Z_2;
    wire sDAC_mem_5Z0Z_3;
    wire sDAC_mem_5Z0Z_4;
    wire sDAC_mem_5Z0Z_5;
    wire sDAC_mem_5Z0Z_6;
    wire sDAC_mem_5Z0Z_7;
    wire sDAC_mem_5_1_sqmuxa;
    wire sDAC_mem_13Z0Z_0;
    wire sDAC_mem_13Z0Z_1;
    wire sDAC_mem_13Z0Z_2;
    wire sDAC_mem_13Z0Z_3;
    wire spi_data_mosi_4;
    wire sDAC_mem_13Z0Z_4;
    wire spi_data_mosi_5;
    wire sDAC_mem_13Z0Z_5;
    wire sDAC_mem_13Z0Z_6;
    wire sDAC_mem_13Z0Z_7;
    wire sDAC_mem_13_1_sqmuxa;
    wire \spi_slave_inst.tx_ready_iZ0 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_4 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_0 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_2 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_2 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_1 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_1 ;
    wire button_debounce_counterZ0Z_1;
    wire button_debounce_counterZ0Z_0;
    wire N_3154_g;
    wire \spi_slave_inst.data_in_reg_iZ0Z_3 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_3 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_6 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_6 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_5 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_5 ;
    wire spi_data_mosi_2;
    wire sCounterADCZ0Z_2;
    wire sEEADC_freqZ0Z_2;
    wire sCounterADCZ0Z_3;
    wire un11_sacqtime_NE_3;
    wire un11_sacqtime_NE_0_0_cascade_;
    wire un11_sacqtime_NE_0;
    wire spi_data_mosi_3;
    wire sEEADC_freqZ0Z_3;
    wire sCounterADCZ0Z_1;
    wire sCounterADCZ0Z_0;
    wire un11_sacqtime_NE_1;
    wire spi_data_mosi_0;
    wire sEEADC_freqZ0Z_0;
    wire sEEADC_freqZ0Z_1;
    wire sCounterADCZ0Z_7;
    wire sCounterADCZ0Z_6;
    wire un11_sacqtime_NE_2;
    wire ADC7_c;
    wire RAM_DATA_1Z0Z_8;
    wire ADC8_c;
    wire RAM_DATA_1Z0Z_9;
    wire top_tour2_c;
    wire RAM_DATA_1Z0Z_12;
    wire spi_miso_ft_c;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_8 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8 ;
    wire sDAC_spi_startZ0;
    wire \spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_ ;
    wire spi_select_c;
    wire spi_cs_ft_c;
    wire \spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_ ;
    wire spi_cs_rpi_c;
    wire \spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1 ;
    wire \spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3 ;
    wire \spi_slave_inst.N_1393_cascade_ ;
    wire spi_miso;
    wire \spi_slave_inst.txdata_reg_iZ0Z_0 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_4 ;
    wire \spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0_cascade_ ;
    wire \spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2 ;
    wire \spi_slave_inst.N_1396 ;
    wire N_23_mux_cascade_;
    wire N_25_mux_cascade_;
    wire m15_1;
    wire op_eq_scounterdac10;
    wire m8_2;
    wire N_23_mux;
    wire N_30_mux_cascade_;
    wire N_25_mux;
    wire N_32_mux;
    wire sCounterDACZ0Z_0;
    wire sCounterDACZ0Z_1;
    wire bfn_20_10_0_;
    wire sCounterDACZ0Z_2;
    wire un2_scounterdac_cry_1;
    wire sCounterDACZ0Z_3;
    wire un2_scounterdac_cry_2;
    wire sCounterDACZ0Z_4;
    wire un2_scounterdac_cry_3;
    wire sCounterDACZ0Z_5;
    wire un2_scounterdac_cry_4;
    wire sCounterDACZ0Z_6;
    wire un2_scounterdac_cry_5_THRU_CO;
    wire un2_scounterdac_cry_5;
    wire sCounterDACZ0Z_7;
    wire un2_scounterdac_cry_6;
    wire N_30_mux;
    wire sCounterDACZ0Z_8;
    wire un2_scounterdac_cry_7;
    wire un2_scounterdac_cry_8;
    wire bfn_20_11_0_;
    wire sCounterDACZ0Z_9;
    wire pll_clk64_0_g;
    wire \spi_slave_inst.un23_i_ssn_3 ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4 ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3 ;
    wire \spi_slave_inst.rx_done_pos_sclk_iZ0 ;
    wire spi_sclk_g;
    wire \spi_slave_inst.spi_cs_iZ0 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_7 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_7 ;
    wire spi_data_mosi_6;
    wire sEEADC_freqZ0Z_6;
    wire spi_data_mosi_7;
    wire sEEADC_freqZ0Z_7;
    wire sEEADC_freq_1_sqmuxa;
    wire N_71;
    wire LED3_c;
    wire un4_sacqtime_cry_23_c_RNITTSZ0Z3;
    wire RAM_DATA_cl_5Z0Z_15;
    wire \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0 ;
    wire bfn_22_7_0_;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1 ;
    wire \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2 ;
    wire \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3 ;
    wire \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4 ;
    wire \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3 ;
    wire \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5 ;
    wire \spi_slave_inst.spi_csZ0 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_i6 ;
    wire \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ;
    wire \spi_slave_inst.tx_done_neg_sclk_iZ0 ;
    wire \spi_slave_inst.tx_done_reg1_iZ0 ;
    wire \spi_slave_inst.tx_done_reg3_iZ0 ;
    wire \spi_slave_inst.tx_done_reg2_iZ0 ;
    wire \spi_slave_inst.un4_tx_done_reg2_i ;
    wire spi_data_mosi_1;
    wire sDAC_mem_25Z0Z_1;
    wire sDAC_mem_25_1_sqmuxa;
    wire CONSTANT_ONE_NET;
    wire RAM_DATA_1Z0Z_15;
    wire _gnd_net_;
    wire pll_clk128_g;
    wire N_31_i;
    wire LED3_c_i_g;

    defparam \pll128M2_inst.pll128M2_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll128M2_inst.pll128M2_inst .TEST_MODE=1'b0;
    defparam \pll128M2_inst.pll128M2_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll128M2_inst.pll128M2_inst .PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam \pll128M2_inst.pll128M2_inst .PLLOUT_SELECT_PORTA="GENCLK";
    defparam \pll128M2_inst.pll128M2_inst .FILTER_RANGE=3'b001;
    defparam \pll128M2_inst.pll128M2_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll128M2_inst.pll128M2_inst .FDA_RELATIVE=4'b0000;
    defparam \pll128M2_inst.pll128M2_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll128M2_inst.pll128M2_inst .ENABLE_ICEGATE_PORTB=1'b0;
    defparam \pll128M2_inst.pll128M2_inst .ENABLE_ICEGATE_PORTA=1'b0;
    defparam \pll128M2_inst.pll128M2_inst .DIVR=4'b0000;
    defparam \pll128M2_inst.pll128M2_inst .DIVQ=3'b011;
    defparam \pll128M2_inst.pll128M2_inst .DIVF=7'b1010100;
    defparam \pll128M2_inst.pll128M2_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE \pll128M2_inst.pll128M2_inst  (
            .EXTFEEDBACK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(\pll128M2_inst.pll_clk64_0 ),
            .REFERENCECLK(N__20270),
            .RESETB(N__49049),
            .BYPASS(GNDG0),
            .PLLOUTCOREA(\pll128M2_inst.pll_clk128 ),
            .SDI(GNDG0),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(GNDG0),
            .PLLOUTGLOBALA(),
            .SCLK(GNDG0));
    IO_PAD RAM_ADD_obuf_5_iopad (
            .OE(N__53520),
            .DIN(N__53519),
            .DOUT(N__53518),
            .PACKAGEPIN(RAM_ADD[5]));
    defparam RAM_ADD_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_5_preio (
            .PADOEN(N__53520),
            .PADOUT(N__53519),
            .PADIN(N__53518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35216),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_mosi_rpi_ibuf_iopad (
            .OE(N__53511),
            .DIN(N__53510),
            .DOUT(N__53509),
            .PACKAGEPIN(spi_mosi_rpi));
    defparam spi_mosi_rpi_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_mosi_rpi_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_mosi_rpi_ibuf_preio (
            .PADOEN(N__53511),
            .PADOUT(N__53510),
            .PADIN(N__53509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_mosi_rpi_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_sclk_rpi_ibuf_iopad (
            .OE(N__53502),
            .DIN(N__53501),
            .DOUT(N__53500),
            .PACKAGEPIN(spi_sclk_rpi));
    defparam spi_sclk_rpi_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_sclk_rpi_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_sclk_rpi_ibuf_preio (
            .PADOEN(N__53502),
            .PADOUT(N__53501),
            .PADIN(N__53500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_sclk_rpi_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_miso_ft_obuf_iopad (
            .OE(N__53493),
            .DIN(N__53492),
            .DOUT(N__53491),
            .PACKAGEPIN(spi_miso_ft));
    defparam spi_miso_ft_obuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_miso_ft_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO spi_miso_ft_obuf_preio (
            .PADOEN(N__53493),
            .PADOUT(N__53492),
            .PADIN(N__53491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__47600),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC5_ibuf_iopad (
            .OE(N__53484),
            .DIN(N__53483),
            .DOUT(N__53482),
            .PACKAGEPIN(ADC5));
    defparam ADC5_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC5_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC5_ibuf_preio (
            .PADOEN(N__53484),
            .PADOUT(N__53483),
            .PADIN(N__53482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC5_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_ACQ_obuf_iopad (
            .OE(N__53475),
            .DIN(N__53474),
            .DOUT(N__53473),
            .PACKAGEPIN(LED_ACQ));
    defparam LED_ACQ_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED_ACQ_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_ACQ_obuf_preio (
            .PADOEN(N__53475),
            .PADOUT(N__53474),
            .PADIN(N__53473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23318),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD reset_rpi_ibuf_iopad (
            .OE(N__53466),
            .DIN(N__53465),
            .DOUT(N__53464),
            .PACKAGEPIN(reset_rpi));
    defparam reset_rpi_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam reset_rpi_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_rpi_ibuf_preio (
            .PADOEN(N__53466),
            .PADOUT(N__53465),
            .PADIN(N__53464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(LED3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_6_iopad (
            .OE(N__53457),
            .DIN(N__53456),
            .DOUT(N__53455),
            .PACKAGEPIN(RAM_DATA[6]));
    defparam RAM_DATA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_6_preio (
            .PADOEN(N__53457),
            .PADOUT(N__53456),
            .PADIN(N__53455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__43172),
            .DIN0(RAM_DATA_in_6),
            .DOUT0(N__26861),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_9_iopad (
            .OE(N__53448),
            .DIN(N__53447),
            .DOUT(N__53446),
            .PACKAGEPIN(RAM_ADD[9]));
    defparam RAM_ADD_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_9_preio (
            .PADOEN(N__53448),
            .PADOUT(N__53447),
            .PADIN(N__53446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36218),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_11_iopad (
            .OE(N__53439),
            .DIN(N__53438),
            .DOUT(N__53437),
            .PACKAGEPIN(RAM_DATA[11]));
    defparam RAM_DATA_iobuf_11_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_11_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_11_preio (
            .PADOEN(N__53439),
            .PADOUT(N__53438),
            .PADIN(N__53437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__39428),
            .DIN0(RAM_DATA_in_11),
            .DOUT0(N__26594),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD trig_rpi_ibuf_iopad (
            .OE(N__53430),
            .DIN(N__53429),
            .DOUT(N__53428),
            .PACKAGEPIN(trig_rpi));
    defparam trig_rpi_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam trig_rpi_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO trig_rpi_ibuf_preio (
            .PADOEN(N__53430),
            .PADOUT(N__53429),
            .PADIN(N__53428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(trig_rpi_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_0_iopad (
            .OE(N__53421),
            .DIN(N__53420),
            .DOUT(N__53419),
            .PACKAGEPIN(RAM_DATA[0]));
    defparam RAM_DATA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_0_preio (
            .PADOEN(N__53421),
            .PADOUT(N__53420),
            .PADIN(N__53419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__39071),
            .DIN0(RAM_DATA_in_0),
            .DOUT0(N__26822),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC2_ibuf_iopad (
            .OE(N__53412),
            .DIN(N__53411),
            .DOUT(N__53410),
            .PACKAGEPIN(ADC2));
    defparam ADC2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC2_ibuf_preio (
            .PADOEN(N__53412),
            .PADOUT(N__53411),
            .PADIN(N__53410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_18_iopad (
            .OE(N__53403),
            .DIN(N__53402),
            .DOUT(N__53401),
            .PACKAGEPIN(RAM_ADD[18]));
    defparam RAM_ADD_obuf_18_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_18_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_18_preio (
            .PADOEN(N__53403),
            .PADOUT(N__53402),
            .PADIN(N__53401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36290),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_2_iopad (
            .OE(N__53394),
            .DIN(N__53393),
            .DOUT(N__53392),
            .PACKAGEPIN(RAM_ADD[2]));
    defparam RAM_ADD_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_2_preio (
            .PADOEN(N__53394),
            .PADOUT(N__53393),
            .PADIN(N__53392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36089),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DAC_mosi_obuf_iopad (
            .OE(N__53385),
            .DIN(N__53384),
            .DOUT(N__53383),
            .PACKAGEPIN(DAC_mosi));
    defparam DAC_mosi_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DAC_mosi_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DAC_mosi_obuf_preio (
            .PADOEN(N__53385),
            .PADOUT(N__53384),
            .PADIN(N__53383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20810),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_13_iopad (
            .OE(N__53376),
            .DIN(N__53375),
            .DOUT(N__53374),
            .PACKAGEPIN(RAM_ADD[13]));
    defparam RAM_ADD_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_13_preio (
            .PADOEN(N__53376),
            .PADOUT(N__53375),
            .PADIN(N__53374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35594),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_nWE_obuf_iopad (
            .OE(N__53367),
            .DIN(N__53366),
            .DOUT(N__53365),
            .PACKAGEPIN(RAM_nWE));
    defparam RAM_nWE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAM_nWE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_nWE_obuf_preio (
            .PADOEN(N__53367),
            .PADOUT(N__53366),
            .PADIN(N__53365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33671),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_7_iopad (
            .OE(N__53358),
            .DIN(N__53357),
            .DOUT(N__53356),
            .PACKAGEPIN(RAM_DATA[7]));
    defparam RAM_DATA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_7_preio (
            .PADOEN(N__53358),
            .PADOUT(N__53357),
            .PADIN(N__53356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__39755),
            .DIN0(RAM_DATA_in_7),
            .DOUT0(N__39701),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC0_ibuf_iopad (
            .OE(N__53349),
            .DIN(N__53348),
            .DOUT(N__53347),
            .PACKAGEPIN(ADC0));
    defparam ADC0_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC0_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC0_ibuf_preio (
            .PADOEN(N__53349),
            .PADOUT(N__53348),
            .PADIN(N__53347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC0_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_nLB_obuf_iopad (
            .OE(N__53340),
            .DIN(N__53339),
            .DOUT(N__53338),
            .PACKAGEPIN(RAM_nLB));
    defparam RAM_nLB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAM_nLB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_nLB_obuf_preio (
            .PADOEN(N__53340),
            .PADOUT(N__53339),
            .PADIN(N__53338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_10_iopad (
            .OE(N__53331),
            .DIN(N__53330),
            .DOUT(N__53329),
            .PACKAGEPIN(RAM_DATA[10]));
    defparam RAM_DATA_iobuf_10_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_10_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_10_preio (
            .PADOEN(N__53331),
            .PADOUT(N__53330),
            .PADIN(N__53329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__39461),
            .DIN0(RAM_DATA_in_10),
            .DOUT0(N__26627),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_1_iopad (
            .OE(N__53322),
            .DIN(N__53321),
            .DOUT(N__53320),
            .PACKAGEPIN(RAM_DATA[1]));
    defparam RAM_DATA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_1_preio (
            .PADOEN(N__53322),
            .PADOUT(N__53321),
            .PADIN(N__53320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__44015),
            .DIN0(RAM_DATA_in_1),
            .DOUT0(N__26660),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_select_ibuf_iopad (
            .OE(N__53313),
            .DIN(N__53312),
            .DOUT(N__53311),
            .PACKAGEPIN(spi_select));
    defparam spi_select_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_select_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_select_ibuf_preio (
            .PADOEN(N__53313),
            .PADOUT(N__53312),
            .PADIN(N__53311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_select_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_nCE_obuf_iopad (
            .OE(N__53304),
            .DIN(N__53303),
            .DOUT(N__53302),
            .PACKAGEPIN(RAM_nCE));
    defparam RAM_nCE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAM_nCE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_nCE_obuf_preio (
            .PADOEN(N__53304),
            .PADOUT(N__53303),
            .PADIN(N__53302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_sclk_flash_obuf_iopad (
            .OE(N__53295),
            .DIN(N__53294),
            .DOUT(N__53293),
            .PACKAGEPIN(spi_sclk_flash));
    defparam spi_sclk_flash_obuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_sclk_flash_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO spi_sclk_flash_obuf_preio (
            .PADOEN(N__53295),
            .PADOUT(N__53294),
            .PADIN(N__53293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_3_iopad (
            .OE(N__53286),
            .DIN(N__53285),
            .DOUT(N__53284),
            .PACKAGEPIN(RAM_ADD[3]));
    defparam RAM_ADD_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_3_preio (
            .PADOEN(N__53286),
            .PADOUT(N__53285),
            .PADIN(N__53284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__43244),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_12_iopad (
            .OE(N__53277),
            .DIN(N__53276),
            .DOUT(N__53275),
            .PACKAGEPIN(RAM_ADD[12]));
    defparam RAM_ADD_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_12_preio (
            .PADOEN(N__53277),
            .PADOUT(N__53276),
            .PADIN(N__53275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35660),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC3_ibuf_iopad (
            .OE(N__53268),
            .DIN(N__53267),
            .DOUT(N__53266),
            .PACKAGEPIN(ADC3));
    defparam ADC3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC3_ibuf_preio (
            .PADOEN(N__53268),
            .PADOUT(N__53267),
            .PADIN(N__53266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_15_iopad (
            .OE(N__53259),
            .DIN(N__53258),
            .DOUT(N__53257),
            .PACKAGEPIN(RAM_DATA[15]));
    defparam RAM_DATA_iobuf_15_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_15_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_15_preio (
            .PADOEN(N__53259),
            .PADOUT(N__53258),
            .PADIN(N__53257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__43142),
            .DIN0(RAM_DATA_in_15),
            .DOUT0(N__52367),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pon_obuf_iopad (
            .OE(N__53250),
            .DIN(N__53249),
            .DOUT(N__53248),
            .PACKAGEPIN(pon));
    defparam pon_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pon_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pon_obuf_preio (
            .PADOEN(N__53250),
            .PADOUT(N__53249),
            .PADIN(N__53248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24014),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DAC_sclk_obuf_iopad (
            .OE(N__53241),
            .DIN(N__53240),
            .DOUT(N__53239),
            .PACKAGEPIN(DAC_sclk));
    defparam DAC_sclk_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DAC_sclk_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DAC_sclk_obuf_preio (
            .PADOEN(N__53241),
            .PADOUT(N__53240),
            .PADIN(N__53239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20888),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_4_iopad (
            .OE(N__53232),
            .DIN(N__53231),
            .DOUT(N__53230),
            .PACKAGEPIN(RAM_DATA[4]));
    defparam RAM_DATA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_4_preio (
            .PADOEN(N__53232),
            .PADOUT(N__53231),
            .PADIN(N__53230),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__39785),
            .DIN0(RAM_DATA_in_4),
            .DOUT0(N__35930),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC1_ibuf_iopad (
            .OE(N__53223),
            .DIN(N__53222),
            .DOUT(N__53221),
            .PACKAGEPIN(ADC1));
    defparam ADC1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC1_ibuf_preio (
            .PADOEN(N__53223),
            .PADOUT(N__53222),
            .PADIN(N__53221),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_cs_flash_obuf_iopad (
            .OE(N__53214),
            .DIN(N__53213),
            .DOUT(N__53212),
            .PACKAGEPIN(spi_cs_flash));
    defparam spi_cs_flash_obuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_cs_flash_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO spi_cs_flash_obuf_preio (
            .PADOEN(N__53214),
            .PADOUT(N__53213),
            .PADIN(N__53212),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD trig_ext_ibuf_iopad (
            .OE(N__53205),
            .DIN(N__53204),
            .DOUT(N__53203),
            .PACKAGEPIN(trig_ext));
    defparam trig_ext_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam trig_ext_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO trig_ext_ibuf_preio (
            .PADOEN(N__53205),
            .PADOUT(N__53204),
            .PADIN(N__53203),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(trig_ext_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_6_iopad (
            .OE(N__53196),
            .DIN(N__53195),
            .DOUT(N__53194),
            .PACKAGEPIN(RAM_ADD[6]));
    defparam RAM_ADD_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_6_preio (
            .PADOEN(N__53196),
            .PADOUT(N__53195),
            .PADIN(N__53194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35972),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD top_tour1_ibuf_iopad (
            .OE(N__53187),
            .DIN(N__53186),
            .DOUT(N__53185),
            .PACKAGEPIN(top_tour1));
    defparam top_tour1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam top_tour1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO top_tour1_ibuf_preio (
            .PADOEN(N__53187),
            .PADOUT(N__53186),
            .PADIN(N__53185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(top_tour1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_17_iopad (
            .OE(N__53178),
            .DIN(N__53177),
            .DOUT(N__53176),
            .PACKAGEPIN(RAM_ADD[17]));
    defparam RAM_ADD_obuf_17_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_17_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_17_preio (
            .PADOEN(N__53178),
            .PADOUT(N__53177),
            .PADIN(N__53176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36356),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_0_iopad (
            .OE(N__53169),
            .DIN(N__53168),
            .DOUT(N__53167),
            .PACKAGEPIN(RAM_ADD[0]));
    defparam RAM_ADD_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_0_preio (
            .PADOEN(N__53169),
            .PADOUT(N__53168),
            .PADIN(N__53167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35861),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_MODE_obuf_iopad (
            .OE(N__53160),
            .DIN(N__53159),
            .DOUT(N__53158),
            .PACKAGEPIN(LED_MODE));
    defparam LED_MODE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED_MODE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_MODE_obuf_preio (
            .PADOEN(N__53160),
            .PADOUT(N__53159),
            .PADIN(N__53158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23618),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_nUB_obuf_iopad (
            .OE(N__53151),
            .DIN(N__53150),
            .DOUT(N__53149),
            .PACKAGEPIN(RAM_nUB));
    defparam RAM_nUB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAM_nUB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_nUB_obuf_preio (
            .PADOEN(N__53151),
            .PADOUT(N__53150),
            .PADIN(N__53149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_11_iopad (
            .OE(N__53142),
            .DIN(N__53141),
            .DOUT(N__53140),
            .PACKAGEPIN(RAM_ADD[11]));
    defparam RAM_ADD_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_11_preio (
            .PADOEN(N__53142),
            .PADOUT(N__53141),
            .PADIN(N__53140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35726),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_14_iopad (
            .OE(N__53133),
            .DIN(N__53132),
            .DOUT(N__53131),
            .PACKAGEPIN(RAM_DATA[14]));
    defparam RAM_DATA_iobuf_14_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_14_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_14_preio (
            .PADOEN(N__53133),
            .PADOUT(N__53132),
            .PADIN(N__53131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__43988),
            .DIN0(RAM_DATA_in_14),
            .DOUT0(N__26933),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DAC_cs_obuf_iopad (
            .OE(N__53124),
            .DIN(N__53123),
            .DOUT(N__53122),
            .PACKAGEPIN(DAC_cs));
    defparam DAC_cs_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DAC_cs_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DAC_cs_obuf_preio (
            .PADOEN(N__53124),
            .PADOUT(N__53123),
            .PADIN(N__53122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20471),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC8_ibuf_iopad (
            .OE(N__53115),
            .DIN(N__53114),
            .DOUT(N__53113),
            .PACKAGEPIN(ADC8));
    defparam ADC8_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC8_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC8_ibuf_preio (
            .PADOEN(N__53115),
            .PADOUT(N__53114),
            .PADIN(N__53113),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC8_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_5_iopad (
            .OE(N__53106),
            .DIN(N__53105),
            .DOUT(N__53104),
            .PACKAGEPIN(RAM_DATA[5]));
    defparam RAM_DATA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_5_preio (
            .PADOEN(N__53106),
            .PADOUT(N__53105),
            .PADIN(N__53104),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__43190),
            .DIN0(RAM_DATA_in_5),
            .DOUT0(N__26702),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC_clk_obuf_iopad (
            .OE(N__53097),
            .DIN(N__53096),
            .DOUT(N__53095),
            .PACKAGEPIN(ADC_clk));
    defparam ADC_clk_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC_clk_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ADC_clk_obuf_preio (
            .PADOEN(N__53097),
            .PADOUT(N__53096),
            .PADIN(N__53095),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34028),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_miso_rpi_obuft_iopad (
            .OE(N__53088),
            .DIN(N__53087),
            .DOUT(N__53086),
            .PACKAGEPIN(spi_miso_rpi));
    defparam spi_miso_rpi_obuft_preio.NEG_TRIGGER=1'b0;
    defparam spi_miso_rpi_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO spi_miso_rpi_obuft_preio (
            .PADOEN(N__53088),
            .PADOUT(N__53087),
            .PADIN(N__53086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__20294),
            .DIN0(),
            .DOUT0(N__47798),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_7_iopad (
            .OE(N__53079),
            .DIN(N__53078),
            .DOUT(N__53077),
            .PACKAGEPIN(RAM_ADD[7]));
    defparam RAM_ADD_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_7_preio (
            .PADOEN(N__53079),
            .PADOUT(N__53078),
            .PADIN(N__53077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36152),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD poff_obuf_iopad (
            .OE(N__53070),
            .DIN(N__53069),
            .DOUT(N__53068),
            .PACKAGEPIN(poff));
    defparam poff_obuf_preio.NEG_TRIGGER=1'b0;
    defparam poff_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO poff_obuf_preio (
            .PADOEN(N__53070),
            .PADOUT(N__53069),
            .PADIN(N__53068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26423),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC4_ibuf_iopad (
            .OE(N__53061),
            .DIN(N__53060),
            .DOUT(N__53059),
            .PACKAGEPIN(ADC4));
    defparam ADC4_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC4_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC4_ibuf_preio (
            .PADOEN(N__53061),
            .PADOUT(N__53060),
            .PADIN(N__53059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC4_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC6_ibuf_iopad (
            .OE(N__53052),
            .DIN(N__53051),
            .DOUT(N__53050),
            .PACKAGEPIN(ADC6));
    defparam ADC6_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC6_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC6_ibuf_preio (
            .PADOEN(N__53052),
            .PADOUT(N__53051),
            .PADIN(N__53050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC6_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_16_iopad (
            .OE(N__53043),
            .DIN(N__53042),
            .DOUT(N__53041),
            .PACKAGEPIN(RAM_ADD[16]));
    defparam RAM_ADD_obuf_16_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_16_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_16_preio (
            .PADOEN(N__53043),
            .PADOUT(N__53042),
            .PADIN(N__53041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35381),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_1_iopad (
            .OE(N__53034),
            .DIN(N__53033),
            .DOUT(N__53032),
            .PACKAGEPIN(RAM_ADD[1]));
    defparam RAM_ADD_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_1_preio (
            .PADOEN(N__53034),
            .PADOUT(N__53033),
            .PADIN(N__53032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36029),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC7_ibuf_iopad (
            .OE(N__53025),
            .DIN(N__53024),
            .DOUT(N__53023),
            .PACKAGEPIN(ADC7));
    defparam ADC7_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC7_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC7_ibuf_preio (
            .PADOEN(N__53025),
            .PADOUT(N__53024),
            .PADIN(N__53023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC7_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD button_mode_ibuf_iopad (
            .OE(N__53016),
            .DIN(N__53015),
            .DOUT(N__53014),
            .PACKAGEPIN(button_mode));
    defparam button_mode_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam button_mode_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO button_mode_ibuf_preio (
            .PADOEN(N__53016),
            .PADOUT(N__53015),
            .PADIN(N__53014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(button_mode_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_sclk_ft_ibuf_iopad (
            .OE(N__53007),
            .DIN(N__53006),
            .DOUT(N__53005),
            .PACKAGEPIN(spi_sclk_ft));
    defparam spi_sclk_ft_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_sclk_ft_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_sclk_ft_ibuf_preio (
            .PADOEN(N__53007),
            .PADOUT(N__53006),
            .PADIN(N__53005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_sclk_ft_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_8_iopad (
            .OE(N__52998),
            .DIN(N__52997),
            .DOUT(N__52996),
            .PACKAGEPIN(RAM_DATA[8]));
    defparam RAM_DATA_iobuf_8_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_8_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_8_preio (
            .PADOEN(N__52998),
            .PADOUT(N__52997),
            .PADIN(N__52996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__39101),
            .DIN0(RAM_DATA_in_8),
            .DOUT0(N__47702),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_10_iopad (
            .OE(N__52989),
            .DIN(N__52988),
            .DOUT(N__52987),
            .PACKAGEPIN(RAM_ADD[10]));
    defparam RAM_ADD_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_10_preio (
            .PADOEN(N__52989),
            .PADOUT(N__52988),
            .PADIN(N__52987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35798),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_13_iopad (
            .OE(N__52980),
            .DIN(N__52979),
            .DOUT(N__52978),
            .PACKAGEPIN(RAM_DATA[13]));
    defparam RAM_DATA_iobuf_13_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_13_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_13_preio (
            .PADOEN(N__52980),
            .PADOUT(N__52979),
            .PADIN(N__52978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__48815),
            .DIN0(RAM_DATA_in_13),
            .DOUT0(N__26546),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD trig_ft_ibuf_iopad (
            .OE(N__52971),
            .DIN(N__52970),
            .DOUT(N__52969),
            .PACKAGEPIN(trig_ft));
    defparam trig_ft_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam trig_ft_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO trig_ft_ibuf_preio (
            .PADOEN(N__52971),
            .PADOUT(N__52970),
            .PADIN(N__52969),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(trig_ft_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC9_ibuf_iopad (
            .OE(N__52962),
            .DIN(N__52961),
            .DOUT(N__52960),
            .PACKAGEPIN(ADC9));
    defparam ADC9_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC9_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC9_ibuf_preio (
            .PADOEN(N__52962),
            .PADOUT(N__52961),
            .PADIN(N__52960),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC9_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_2_iopad (
            .OE(N__52953),
            .DIN(N__52952),
            .DOUT(N__52951),
            .PACKAGEPIN(RAM_DATA[2]));
    defparam RAM_DATA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_2_preio (
            .PADOEN(N__52953),
            .PADOUT(N__52952),
            .PADIN(N__52951),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__39725),
            .DIN0(RAM_DATA_in_2),
            .DOUT0(N__26894),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD cs_rpi2flash_ibuf_iopad (
            .OE(N__52944),
            .DIN(N__52943),
            .DOUT(N__52942),
            .PACKAGEPIN(cs_rpi2flash));
    defparam cs_rpi2flash_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam cs_rpi2flash_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO cs_rpi2flash_ibuf_preio (
            .PADOEN(N__52944),
            .PADOUT(N__52943),
            .PADIN(N__52942),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(cs_rpi2flash_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED3_obuf_iopad (
            .OE(N__52935),
            .DIN(N__52934),
            .DOUT(N__52933),
            .PACKAGEPIN(LED3));
    defparam LED3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED3_obuf_preio (
            .PADOEN(N__52935),
            .PADOUT(N__52934),
            .PADIN(N__52933),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__49419),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_mosi_ft_ibuf_iopad (
            .OE(N__52926),
            .DIN(N__52925),
            .DOUT(N__52924),
            .PACKAGEPIN(spi_mosi_ft));
    defparam spi_mosi_ft_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_mosi_ft_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_mosi_ft_ibuf_preio (
            .PADOEN(N__52926),
            .PADOUT(N__52925),
            .PADIN(N__52924),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_mosi_ft_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_nOE_obuf_iopad (
            .OE(N__52917),
            .DIN(N__52916),
            .DOUT(N__52915),
            .PACKAGEPIN(RAM_nOE));
    defparam RAM_nOE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAM_nOE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_nOE_obuf_preio (
            .PADOEN(N__52917),
            .PADOUT(N__52916),
            .PADIN(N__52915),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_4_iopad (
            .OE(N__52908),
            .DIN(N__52907),
            .DOUT(N__52906),
            .PACKAGEPIN(RAM_ADD[4]));
    defparam RAM_ADD_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_4_preio (
            .PADOEN(N__52908),
            .PADOUT(N__52907),
            .PADIN(N__52906),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__43538),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_ibuf_iopad (
            .OE(N__52899),
            .DIN(N__52898),
            .DOUT(N__52897),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_preio (
            .PADOEN(N__52899),
            .PADOUT(N__52898),
            .PADIN(N__52897),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD top_tour2_ibuf_iopad (
            .OE(N__52890),
            .DIN(N__52889),
            .DOUT(N__52888),
            .PACKAGEPIN(top_tour2));
    defparam top_tour2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam top_tour2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO top_tour2_ibuf_preio (
            .PADOEN(N__52890),
            .PADOUT(N__52889),
            .PADIN(N__52888),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(top_tour2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_cs_rpi_ibuf_iopad (
            .OE(N__52881),
            .DIN(N__52880),
            .DOUT(N__52879),
            .PACKAGEPIN(spi_cs_rpi));
    defparam spi_cs_rpi_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_cs_rpi_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_cs_rpi_ibuf_preio (
            .PADOEN(N__52881),
            .PADOUT(N__52880),
            .PADIN(N__52879),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_cs_rpi_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_15_iopad (
            .OE(N__52872),
            .DIN(N__52871),
            .DOUT(N__52870),
            .PACKAGEPIN(RAM_ADD[15]));
    defparam RAM_ADD_obuf_15_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_15_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_15_preio (
            .PADOEN(N__52872),
            .PADOUT(N__52871),
            .PADIN(N__52870),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35453),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_9_iopad (
            .OE(N__52863),
            .DIN(N__52862),
            .DOUT(N__52861),
            .PACKAGEPIN(RAM_DATA[9]));
    defparam RAM_DATA_iobuf_9_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_9_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_9_preio (
            .PADOEN(N__52863),
            .PADOUT(N__52862),
            .PADIN(N__52861),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__43115),
            .DIN0(RAM_DATA_in_9),
            .DOUT0(N__47657),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_8_iopad (
            .OE(N__52854),
            .DIN(N__52853),
            .DOUT(N__52852),
            .PACKAGEPIN(RAM_ADD[8]));
    defparam RAM_ADD_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_8_preio (
            .PADOEN(N__52854),
            .PADOUT(N__52853),
            .PADIN(N__52852),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__43610),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_12_iopad (
            .OE(N__52845),
            .DIN(N__52844),
            .DOUT(N__52843),
            .PACKAGEPIN(RAM_DATA[12]));
    defparam RAM_DATA_iobuf_12_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_12_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_12_preio (
            .PADOEN(N__52845),
            .PADOUT(N__52844),
            .PADIN(N__52843),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__44075),
            .DIN0(RAM_DATA_in_12),
            .DOUT0(N__47618),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_3_iopad (
            .OE(N__52836),
            .DIN(N__52835),
            .DOUT(N__52834),
            .PACKAGEPIN(RAM_DATA[3]));
    defparam RAM_DATA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_3_preio (
            .PADOEN(N__52836),
            .PADOUT(N__52835),
            .PADIN(N__52834),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__44045),
            .DIN0(RAM_DATA_in_3),
            .DOUT0(N__33944),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_cs_ft_ibuf_iopad (
            .OE(N__52827),
            .DIN(N__52826),
            .DOUT(N__52825),
            .PACKAGEPIN(spi_cs_ft));
    defparam spi_cs_ft_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_cs_ft_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_cs_ft_ibuf_preio (
            .PADOEN(N__52827),
            .PADOUT(N__52826),
            .PADIN(N__52825),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_cs_ft_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_mosi_flash_obuf_iopad (
            .OE(N__52818),
            .DIN(N__52817),
            .DOUT(N__52816),
            .PACKAGEPIN(spi_mosi_flash));
    defparam spi_mosi_flash_obuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_mosi_flash_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO spi_mosi_flash_obuf_preio (
            .PADOEN(N__52818),
            .PADOUT(N__52817),
            .PADIN(N__52816),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_14_iopad (
            .OE(N__52809),
            .DIN(N__52808),
            .DOUT(N__52807),
            .PACKAGEPIN(RAM_ADD[14]));
    defparam RAM_ADD_obuf_14_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_14_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_14_preio (
            .PADOEN(N__52809),
            .PADOUT(N__52808),
            .PADIN(N__52807),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35528),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__12567 (
            .O(N__52790),
            .I(N__52770));
    InMux I__12566 (
            .O(N__52789),
            .I(N__52770));
    InMux I__12565 (
            .O(N__52788),
            .I(N__52770));
    InMux I__12564 (
            .O(N__52787),
            .I(N__52770));
    CascadeMux I__12563 (
            .O(N__52786),
            .I(N__52760));
    CascadeMux I__12562 (
            .O(N__52785),
            .I(N__52756));
    CascadeMux I__12561 (
            .O(N__52784),
            .I(N__52752));
    CascadeMux I__12560 (
            .O(N__52783),
            .I(N__52748));
    CascadeMux I__12559 (
            .O(N__52782),
            .I(N__52739));
    InMux I__12558 (
            .O(N__52781),
            .I(N__52731));
    InMux I__12557 (
            .O(N__52780),
            .I(N__52731));
    InMux I__12556 (
            .O(N__52779),
            .I(N__52731));
    LocalMux I__12555 (
            .O(N__52770),
            .I(N__52728));
    InMux I__12554 (
            .O(N__52769),
            .I(N__52721));
    InMux I__12553 (
            .O(N__52768),
            .I(N__52721));
    InMux I__12552 (
            .O(N__52767),
            .I(N__52721));
    InMux I__12551 (
            .O(N__52766),
            .I(N__52712));
    InMux I__12550 (
            .O(N__52765),
            .I(N__52712));
    InMux I__12549 (
            .O(N__52764),
            .I(N__52712));
    InMux I__12548 (
            .O(N__52763),
            .I(N__52712));
    InMux I__12547 (
            .O(N__52760),
            .I(N__52688));
    InMux I__12546 (
            .O(N__52759),
            .I(N__52688));
    InMux I__12545 (
            .O(N__52756),
            .I(N__52688));
    InMux I__12544 (
            .O(N__52755),
            .I(N__52688));
    InMux I__12543 (
            .O(N__52752),
            .I(N__52688));
    InMux I__12542 (
            .O(N__52751),
            .I(N__52688));
    InMux I__12541 (
            .O(N__52748),
            .I(N__52688));
    InMux I__12540 (
            .O(N__52747),
            .I(N__52688));
    CascadeMux I__12539 (
            .O(N__52746),
            .I(N__52685));
    CascadeMux I__12538 (
            .O(N__52745),
            .I(N__52681));
    CascadeMux I__12537 (
            .O(N__52744),
            .I(N__52677));
    CascadeMux I__12536 (
            .O(N__52743),
            .I(N__52673));
    InMux I__12535 (
            .O(N__52742),
            .I(N__52661));
    InMux I__12534 (
            .O(N__52739),
            .I(N__52661));
    InMux I__12533 (
            .O(N__52738),
            .I(N__52661));
    LocalMux I__12532 (
            .O(N__52731),
            .I(N__52658));
    Span4Mux_h I__12531 (
            .O(N__52728),
            .I(N__52651));
    LocalMux I__12530 (
            .O(N__52721),
            .I(N__52651));
    LocalMux I__12529 (
            .O(N__52712),
            .I(N__52651));
    CascadeMux I__12528 (
            .O(N__52711),
            .I(N__52646));
    CascadeMux I__12527 (
            .O(N__52710),
            .I(N__52643));
    CascadeMux I__12526 (
            .O(N__52709),
            .I(N__52640));
    CascadeMux I__12525 (
            .O(N__52708),
            .I(N__52636));
    CascadeMux I__12524 (
            .O(N__52707),
            .I(N__52633));
    CascadeMux I__12523 (
            .O(N__52706),
            .I(N__52630));
    CascadeMux I__12522 (
            .O(N__52705),
            .I(N__52627));
    LocalMux I__12521 (
            .O(N__52688),
            .I(N__52620));
    InMux I__12520 (
            .O(N__52685),
            .I(N__52603));
    InMux I__12519 (
            .O(N__52684),
            .I(N__52603));
    InMux I__12518 (
            .O(N__52681),
            .I(N__52603));
    InMux I__12517 (
            .O(N__52680),
            .I(N__52603));
    InMux I__12516 (
            .O(N__52677),
            .I(N__52603));
    InMux I__12515 (
            .O(N__52676),
            .I(N__52603));
    InMux I__12514 (
            .O(N__52673),
            .I(N__52603));
    InMux I__12513 (
            .O(N__52672),
            .I(N__52603));
    CascadeMux I__12512 (
            .O(N__52671),
            .I(N__52599));
    CascadeMux I__12511 (
            .O(N__52670),
            .I(N__52595));
    CascadeMux I__12510 (
            .O(N__52669),
            .I(N__52591));
    CascadeMux I__12509 (
            .O(N__52668),
            .I(N__52587));
    LocalMux I__12508 (
            .O(N__52661),
            .I(N__52579));
    Span4Mux_v I__12507 (
            .O(N__52658),
            .I(N__52579));
    Span4Mux_v I__12506 (
            .O(N__52651),
            .I(N__52579));
    InMux I__12505 (
            .O(N__52650),
            .I(N__52574));
    InMux I__12504 (
            .O(N__52649),
            .I(N__52574));
    InMux I__12503 (
            .O(N__52646),
            .I(N__52563));
    InMux I__12502 (
            .O(N__52643),
            .I(N__52563));
    InMux I__12501 (
            .O(N__52640),
            .I(N__52563));
    InMux I__12500 (
            .O(N__52639),
            .I(N__52552));
    InMux I__12499 (
            .O(N__52636),
            .I(N__52552));
    InMux I__12498 (
            .O(N__52633),
            .I(N__52552));
    InMux I__12497 (
            .O(N__52630),
            .I(N__52552));
    InMux I__12496 (
            .O(N__52627),
            .I(N__52552));
    CascadeMux I__12495 (
            .O(N__52626),
            .I(N__52549));
    CascadeMux I__12494 (
            .O(N__52625),
            .I(N__52545));
    CascadeMux I__12493 (
            .O(N__52624),
            .I(N__52541));
    CascadeMux I__12492 (
            .O(N__52623),
            .I(N__52537));
    Span4Mux_v I__12491 (
            .O(N__52620),
            .I(N__52531));
    LocalMux I__12490 (
            .O(N__52603),
            .I(N__52531));
    InMux I__12489 (
            .O(N__52602),
            .I(N__52514));
    InMux I__12488 (
            .O(N__52599),
            .I(N__52514));
    InMux I__12487 (
            .O(N__52598),
            .I(N__52514));
    InMux I__12486 (
            .O(N__52595),
            .I(N__52514));
    InMux I__12485 (
            .O(N__52594),
            .I(N__52514));
    InMux I__12484 (
            .O(N__52591),
            .I(N__52514));
    InMux I__12483 (
            .O(N__52590),
            .I(N__52514));
    InMux I__12482 (
            .O(N__52587),
            .I(N__52514));
    CascadeMux I__12481 (
            .O(N__52586),
            .I(N__52511));
    Span4Mux_v I__12480 (
            .O(N__52579),
            .I(N__52507));
    LocalMux I__12479 (
            .O(N__52574),
            .I(N__52504));
    CascadeMux I__12478 (
            .O(N__52573),
            .I(N__52500));
    CascadeMux I__12477 (
            .O(N__52572),
            .I(N__52496));
    CascadeMux I__12476 (
            .O(N__52571),
            .I(N__52492));
    CascadeMux I__12475 (
            .O(N__52570),
            .I(N__52488));
    LocalMux I__12474 (
            .O(N__52563),
            .I(N__52485));
    LocalMux I__12473 (
            .O(N__52552),
            .I(N__52482));
    InMux I__12472 (
            .O(N__52549),
            .I(N__52465));
    InMux I__12471 (
            .O(N__52548),
            .I(N__52465));
    InMux I__12470 (
            .O(N__52545),
            .I(N__52465));
    InMux I__12469 (
            .O(N__52544),
            .I(N__52465));
    InMux I__12468 (
            .O(N__52541),
            .I(N__52465));
    InMux I__12467 (
            .O(N__52540),
            .I(N__52465));
    InMux I__12466 (
            .O(N__52537),
            .I(N__52465));
    InMux I__12465 (
            .O(N__52536),
            .I(N__52465));
    Span4Mux_h I__12464 (
            .O(N__52531),
            .I(N__52460));
    LocalMux I__12463 (
            .O(N__52514),
            .I(N__52460));
    InMux I__12462 (
            .O(N__52511),
            .I(N__52455));
    InMux I__12461 (
            .O(N__52510),
            .I(N__52455));
    Span4Mux_h I__12460 (
            .O(N__52507),
            .I(N__52450));
    Span4Mux_v I__12459 (
            .O(N__52504),
            .I(N__52450));
    InMux I__12458 (
            .O(N__52503),
            .I(N__52433));
    InMux I__12457 (
            .O(N__52500),
            .I(N__52433));
    InMux I__12456 (
            .O(N__52499),
            .I(N__52433));
    InMux I__12455 (
            .O(N__52496),
            .I(N__52433));
    InMux I__12454 (
            .O(N__52495),
            .I(N__52433));
    InMux I__12453 (
            .O(N__52492),
            .I(N__52433));
    InMux I__12452 (
            .O(N__52491),
            .I(N__52433));
    InMux I__12451 (
            .O(N__52488),
            .I(N__52433));
    Span4Mux_v I__12450 (
            .O(N__52485),
            .I(N__52428));
    Span4Mux_v I__12449 (
            .O(N__52482),
            .I(N__52428));
    LocalMux I__12448 (
            .O(N__52465),
            .I(N__52425));
    Span4Mux_h I__12447 (
            .O(N__52460),
            .I(N__52420));
    LocalMux I__12446 (
            .O(N__52455),
            .I(N__52420));
    Span4Mux_h I__12445 (
            .O(N__52450),
            .I(N__52417));
    LocalMux I__12444 (
            .O(N__52433),
            .I(N__52414));
    Span4Mux_h I__12443 (
            .O(N__52428),
            .I(N__52409));
    Span4Mux_v I__12442 (
            .O(N__52425),
            .I(N__52409));
    Span4Mux_v I__12441 (
            .O(N__52420),
            .I(N__52405));
    Span4Mux_h I__12440 (
            .O(N__52417),
            .I(N__52402));
    Span4Mux_v I__12439 (
            .O(N__52414),
            .I(N__52399));
    Span4Mux_h I__12438 (
            .O(N__52409),
            .I(N__52396));
    InMux I__12437 (
            .O(N__52408),
            .I(N__52393));
    Span4Mux_v I__12436 (
            .O(N__52405),
            .I(N__52390));
    Span4Mux_v I__12435 (
            .O(N__52402),
            .I(N__52385));
    Span4Mux_h I__12434 (
            .O(N__52399),
            .I(N__52385));
    Span4Mux_h I__12433 (
            .O(N__52396),
            .I(N__52380));
    LocalMux I__12432 (
            .O(N__52393),
            .I(N__52380));
    Span4Mux_h I__12431 (
            .O(N__52390),
            .I(N__52377));
    Span4Mux_h I__12430 (
            .O(N__52385),
            .I(N__52372));
    Span4Mux_v I__12429 (
            .O(N__52380),
            .I(N__52372));
    Odrv4 I__12428 (
            .O(N__52377),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12427 (
            .O(N__52372),
            .I(CONSTANT_ONE_NET));
    IoInMux I__12426 (
            .O(N__52367),
            .I(N__52364));
    LocalMux I__12425 (
            .O(N__52364),
            .I(N__52361));
    IoSpan4Mux I__12424 (
            .O(N__52361),
            .I(N__52358));
    Span4Mux_s3_h I__12423 (
            .O(N__52358),
            .I(N__52355));
    Span4Mux_v I__12422 (
            .O(N__52355),
            .I(N__52352));
    Odrv4 I__12421 (
            .O(N__52352),
            .I(RAM_DATA_1Z0Z_15));
    ClkMux I__12420 (
            .O(N__52349),
            .I(N__51902));
    ClkMux I__12419 (
            .O(N__52348),
            .I(N__51902));
    ClkMux I__12418 (
            .O(N__52347),
            .I(N__51902));
    ClkMux I__12417 (
            .O(N__52346),
            .I(N__51902));
    ClkMux I__12416 (
            .O(N__52345),
            .I(N__51902));
    ClkMux I__12415 (
            .O(N__52344),
            .I(N__51902));
    ClkMux I__12414 (
            .O(N__52343),
            .I(N__51902));
    ClkMux I__12413 (
            .O(N__52342),
            .I(N__51902));
    ClkMux I__12412 (
            .O(N__52341),
            .I(N__51902));
    ClkMux I__12411 (
            .O(N__52340),
            .I(N__51902));
    ClkMux I__12410 (
            .O(N__52339),
            .I(N__51902));
    ClkMux I__12409 (
            .O(N__52338),
            .I(N__51902));
    ClkMux I__12408 (
            .O(N__52337),
            .I(N__51902));
    ClkMux I__12407 (
            .O(N__52336),
            .I(N__51902));
    ClkMux I__12406 (
            .O(N__52335),
            .I(N__51902));
    ClkMux I__12405 (
            .O(N__52334),
            .I(N__51902));
    ClkMux I__12404 (
            .O(N__52333),
            .I(N__51902));
    ClkMux I__12403 (
            .O(N__52332),
            .I(N__51902));
    ClkMux I__12402 (
            .O(N__52331),
            .I(N__51902));
    ClkMux I__12401 (
            .O(N__52330),
            .I(N__51902));
    ClkMux I__12400 (
            .O(N__52329),
            .I(N__51902));
    ClkMux I__12399 (
            .O(N__52328),
            .I(N__51902));
    ClkMux I__12398 (
            .O(N__52327),
            .I(N__51902));
    ClkMux I__12397 (
            .O(N__52326),
            .I(N__51902));
    ClkMux I__12396 (
            .O(N__52325),
            .I(N__51902));
    ClkMux I__12395 (
            .O(N__52324),
            .I(N__51902));
    ClkMux I__12394 (
            .O(N__52323),
            .I(N__51902));
    ClkMux I__12393 (
            .O(N__52322),
            .I(N__51902));
    ClkMux I__12392 (
            .O(N__52321),
            .I(N__51902));
    ClkMux I__12391 (
            .O(N__52320),
            .I(N__51902));
    ClkMux I__12390 (
            .O(N__52319),
            .I(N__51902));
    ClkMux I__12389 (
            .O(N__52318),
            .I(N__51902));
    ClkMux I__12388 (
            .O(N__52317),
            .I(N__51902));
    ClkMux I__12387 (
            .O(N__52316),
            .I(N__51902));
    ClkMux I__12386 (
            .O(N__52315),
            .I(N__51902));
    ClkMux I__12385 (
            .O(N__52314),
            .I(N__51902));
    ClkMux I__12384 (
            .O(N__52313),
            .I(N__51902));
    ClkMux I__12383 (
            .O(N__52312),
            .I(N__51902));
    ClkMux I__12382 (
            .O(N__52311),
            .I(N__51902));
    ClkMux I__12381 (
            .O(N__52310),
            .I(N__51902));
    ClkMux I__12380 (
            .O(N__52309),
            .I(N__51902));
    ClkMux I__12379 (
            .O(N__52308),
            .I(N__51902));
    ClkMux I__12378 (
            .O(N__52307),
            .I(N__51902));
    ClkMux I__12377 (
            .O(N__52306),
            .I(N__51902));
    ClkMux I__12376 (
            .O(N__52305),
            .I(N__51902));
    ClkMux I__12375 (
            .O(N__52304),
            .I(N__51902));
    ClkMux I__12374 (
            .O(N__52303),
            .I(N__51902));
    ClkMux I__12373 (
            .O(N__52302),
            .I(N__51902));
    ClkMux I__12372 (
            .O(N__52301),
            .I(N__51902));
    ClkMux I__12371 (
            .O(N__52300),
            .I(N__51902));
    ClkMux I__12370 (
            .O(N__52299),
            .I(N__51902));
    ClkMux I__12369 (
            .O(N__52298),
            .I(N__51902));
    ClkMux I__12368 (
            .O(N__52297),
            .I(N__51902));
    ClkMux I__12367 (
            .O(N__52296),
            .I(N__51902));
    ClkMux I__12366 (
            .O(N__52295),
            .I(N__51902));
    ClkMux I__12365 (
            .O(N__52294),
            .I(N__51902));
    ClkMux I__12364 (
            .O(N__52293),
            .I(N__51902));
    ClkMux I__12363 (
            .O(N__52292),
            .I(N__51902));
    ClkMux I__12362 (
            .O(N__52291),
            .I(N__51902));
    ClkMux I__12361 (
            .O(N__52290),
            .I(N__51902));
    ClkMux I__12360 (
            .O(N__52289),
            .I(N__51902));
    ClkMux I__12359 (
            .O(N__52288),
            .I(N__51902));
    ClkMux I__12358 (
            .O(N__52287),
            .I(N__51902));
    ClkMux I__12357 (
            .O(N__52286),
            .I(N__51902));
    ClkMux I__12356 (
            .O(N__52285),
            .I(N__51902));
    ClkMux I__12355 (
            .O(N__52284),
            .I(N__51902));
    ClkMux I__12354 (
            .O(N__52283),
            .I(N__51902));
    ClkMux I__12353 (
            .O(N__52282),
            .I(N__51902));
    ClkMux I__12352 (
            .O(N__52281),
            .I(N__51902));
    ClkMux I__12351 (
            .O(N__52280),
            .I(N__51902));
    ClkMux I__12350 (
            .O(N__52279),
            .I(N__51902));
    ClkMux I__12349 (
            .O(N__52278),
            .I(N__51902));
    ClkMux I__12348 (
            .O(N__52277),
            .I(N__51902));
    ClkMux I__12347 (
            .O(N__52276),
            .I(N__51902));
    ClkMux I__12346 (
            .O(N__52275),
            .I(N__51902));
    ClkMux I__12345 (
            .O(N__52274),
            .I(N__51902));
    ClkMux I__12344 (
            .O(N__52273),
            .I(N__51902));
    ClkMux I__12343 (
            .O(N__52272),
            .I(N__51902));
    ClkMux I__12342 (
            .O(N__52271),
            .I(N__51902));
    ClkMux I__12341 (
            .O(N__52270),
            .I(N__51902));
    ClkMux I__12340 (
            .O(N__52269),
            .I(N__51902));
    ClkMux I__12339 (
            .O(N__52268),
            .I(N__51902));
    ClkMux I__12338 (
            .O(N__52267),
            .I(N__51902));
    ClkMux I__12337 (
            .O(N__52266),
            .I(N__51902));
    ClkMux I__12336 (
            .O(N__52265),
            .I(N__51902));
    ClkMux I__12335 (
            .O(N__52264),
            .I(N__51902));
    ClkMux I__12334 (
            .O(N__52263),
            .I(N__51902));
    ClkMux I__12333 (
            .O(N__52262),
            .I(N__51902));
    ClkMux I__12332 (
            .O(N__52261),
            .I(N__51902));
    ClkMux I__12331 (
            .O(N__52260),
            .I(N__51902));
    ClkMux I__12330 (
            .O(N__52259),
            .I(N__51902));
    ClkMux I__12329 (
            .O(N__52258),
            .I(N__51902));
    ClkMux I__12328 (
            .O(N__52257),
            .I(N__51902));
    ClkMux I__12327 (
            .O(N__52256),
            .I(N__51902));
    ClkMux I__12326 (
            .O(N__52255),
            .I(N__51902));
    ClkMux I__12325 (
            .O(N__52254),
            .I(N__51902));
    ClkMux I__12324 (
            .O(N__52253),
            .I(N__51902));
    ClkMux I__12323 (
            .O(N__52252),
            .I(N__51902));
    ClkMux I__12322 (
            .O(N__52251),
            .I(N__51902));
    ClkMux I__12321 (
            .O(N__52250),
            .I(N__51902));
    ClkMux I__12320 (
            .O(N__52249),
            .I(N__51902));
    ClkMux I__12319 (
            .O(N__52248),
            .I(N__51902));
    ClkMux I__12318 (
            .O(N__52247),
            .I(N__51902));
    ClkMux I__12317 (
            .O(N__52246),
            .I(N__51902));
    ClkMux I__12316 (
            .O(N__52245),
            .I(N__51902));
    ClkMux I__12315 (
            .O(N__52244),
            .I(N__51902));
    ClkMux I__12314 (
            .O(N__52243),
            .I(N__51902));
    ClkMux I__12313 (
            .O(N__52242),
            .I(N__51902));
    ClkMux I__12312 (
            .O(N__52241),
            .I(N__51902));
    ClkMux I__12311 (
            .O(N__52240),
            .I(N__51902));
    ClkMux I__12310 (
            .O(N__52239),
            .I(N__51902));
    ClkMux I__12309 (
            .O(N__52238),
            .I(N__51902));
    ClkMux I__12308 (
            .O(N__52237),
            .I(N__51902));
    ClkMux I__12307 (
            .O(N__52236),
            .I(N__51902));
    ClkMux I__12306 (
            .O(N__52235),
            .I(N__51902));
    ClkMux I__12305 (
            .O(N__52234),
            .I(N__51902));
    ClkMux I__12304 (
            .O(N__52233),
            .I(N__51902));
    ClkMux I__12303 (
            .O(N__52232),
            .I(N__51902));
    ClkMux I__12302 (
            .O(N__52231),
            .I(N__51902));
    ClkMux I__12301 (
            .O(N__52230),
            .I(N__51902));
    ClkMux I__12300 (
            .O(N__52229),
            .I(N__51902));
    ClkMux I__12299 (
            .O(N__52228),
            .I(N__51902));
    ClkMux I__12298 (
            .O(N__52227),
            .I(N__51902));
    ClkMux I__12297 (
            .O(N__52226),
            .I(N__51902));
    ClkMux I__12296 (
            .O(N__52225),
            .I(N__51902));
    ClkMux I__12295 (
            .O(N__52224),
            .I(N__51902));
    ClkMux I__12294 (
            .O(N__52223),
            .I(N__51902));
    ClkMux I__12293 (
            .O(N__52222),
            .I(N__51902));
    ClkMux I__12292 (
            .O(N__52221),
            .I(N__51902));
    ClkMux I__12291 (
            .O(N__52220),
            .I(N__51902));
    ClkMux I__12290 (
            .O(N__52219),
            .I(N__51902));
    ClkMux I__12289 (
            .O(N__52218),
            .I(N__51902));
    ClkMux I__12288 (
            .O(N__52217),
            .I(N__51902));
    ClkMux I__12287 (
            .O(N__52216),
            .I(N__51902));
    ClkMux I__12286 (
            .O(N__52215),
            .I(N__51902));
    ClkMux I__12285 (
            .O(N__52214),
            .I(N__51902));
    ClkMux I__12284 (
            .O(N__52213),
            .I(N__51902));
    ClkMux I__12283 (
            .O(N__52212),
            .I(N__51902));
    ClkMux I__12282 (
            .O(N__52211),
            .I(N__51902));
    ClkMux I__12281 (
            .O(N__52210),
            .I(N__51902));
    ClkMux I__12280 (
            .O(N__52209),
            .I(N__51902));
    ClkMux I__12279 (
            .O(N__52208),
            .I(N__51902));
    ClkMux I__12278 (
            .O(N__52207),
            .I(N__51902));
    ClkMux I__12277 (
            .O(N__52206),
            .I(N__51902));
    ClkMux I__12276 (
            .O(N__52205),
            .I(N__51902));
    ClkMux I__12275 (
            .O(N__52204),
            .I(N__51902));
    ClkMux I__12274 (
            .O(N__52203),
            .I(N__51902));
    ClkMux I__12273 (
            .O(N__52202),
            .I(N__51902));
    ClkMux I__12272 (
            .O(N__52201),
            .I(N__51902));
    GlobalMux I__12271 (
            .O(N__51902),
            .I(N__51899));
    gio2CtrlBuf I__12270 (
            .O(N__51899),
            .I(pll_clk128_g));
    CEMux I__12269 (
            .O(N__51896),
            .I(N__51891));
    CEMux I__12268 (
            .O(N__51895),
            .I(N__51886));
    CEMux I__12267 (
            .O(N__51894),
            .I(N__51883));
    LocalMux I__12266 (
            .O(N__51891),
            .I(N__51879));
    CEMux I__12265 (
            .O(N__51890),
            .I(N__51876));
    CEMux I__12264 (
            .O(N__51889),
            .I(N__51873));
    LocalMux I__12263 (
            .O(N__51886),
            .I(N__51869));
    LocalMux I__12262 (
            .O(N__51883),
            .I(N__51866));
    CEMux I__12261 (
            .O(N__51882),
            .I(N__51863));
    Span4Mux_h I__12260 (
            .O(N__51879),
            .I(N__51858));
    LocalMux I__12259 (
            .O(N__51876),
            .I(N__51858));
    LocalMux I__12258 (
            .O(N__51873),
            .I(N__51855));
    CEMux I__12257 (
            .O(N__51872),
            .I(N__51852));
    Span4Mux_h I__12256 (
            .O(N__51869),
            .I(N__51849));
    Span12Mux_s6_h I__12255 (
            .O(N__51866),
            .I(N__51844));
    LocalMux I__12254 (
            .O(N__51863),
            .I(N__51844));
    Span4Mux_h I__12253 (
            .O(N__51858),
            .I(N__51841));
    Span4Mux_v I__12252 (
            .O(N__51855),
            .I(N__51836));
    LocalMux I__12251 (
            .O(N__51852),
            .I(N__51836));
    Odrv4 I__12250 (
            .O(N__51849),
            .I(N_31_i));
    Odrv12 I__12249 (
            .O(N__51844),
            .I(N_31_i));
    Odrv4 I__12248 (
            .O(N__51841),
            .I(N_31_i));
    Odrv4 I__12247 (
            .O(N__51836),
            .I(N_31_i));
    SRMux I__12246 (
            .O(N__51827),
            .I(N__51269));
    SRMux I__12245 (
            .O(N__51826),
            .I(N__51269));
    SRMux I__12244 (
            .O(N__51825),
            .I(N__51269));
    SRMux I__12243 (
            .O(N__51824),
            .I(N__51269));
    SRMux I__12242 (
            .O(N__51823),
            .I(N__51269));
    SRMux I__12241 (
            .O(N__51822),
            .I(N__51269));
    SRMux I__12240 (
            .O(N__51821),
            .I(N__51269));
    SRMux I__12239 (
            .O(N__51820),
            .I(N__51269));
    SRMux I__12238 (
            .O(N__51819),
            .I(N__51269));
    SRMux I__12237 (
            .O(N__51818),
            .I(N__51269));
    SRMux I__12236 (
            .O(N__51817),
            .I(N__51269));
    SRMux I__12235 (
            .O(N__51816),
            .I(N__51269));
    SRMux I__12234 (
            .O(N__51815),
            .I(N__51269));
    SRMux I__12233 (
            .O(N__51814),
            .I(N__51269));
    SRMux I__12232 (
            .O(N__51813),
            .I(N__51269));
    SRMux I__12231 (
            .O(N__51812),
            .I(N__51269));
    SRMux I__12230 (
            .O(N__51811),
            .I(N__51269));
    SRMux I__12229 (
            .O(N__51810),
            .I(N__51269));
    SRMux I__12228 (
            .O(N__51809),
            .I(N__51269));
    SRMux I__12227 (
            .O(N__51808),
            .I(N__51269));
    SRMux I__12226 (
            .O(N__51807),
            .I(N__51269));
    SRMux I__12225 (
            .O(N__51806),
            .I(N__51269));
    SRMux I__12224 (
            .O(N__51805),
            .I(N__51269));
    SRMux I__12223 (
            .O(N__51804),
            .I(N__51269));
    SRMux I__12222 (
            .O(N__51803),
            .I(N__51269));
    SRMux I__12221 (
            .O(N__51802),
            .I(N__51269));
    SRMux I__12220 (
            .O(N__51801),
            .I(N__51269));
    SRMux I__12219 (
            .O(N__51800),
            .I(N__51269));
    SRMux I__12218 (
            .O(N__51799),
            .I(N__51269));
    SRMux I__12217 (
            .O(N__51798),
            .I(N__51269));
    SRMux I__12216 (
            .O(N__51797),
            .I(N__51269));
    SRMux I__12215 (
            .O(N__51796),
            .I(N__51269));
    SRMux I__12214 (
            .O(N__51795),
            .I(N__51269));
    SRMux I__12213 (
            .O(N__51794),
            .I(N__51269));
    SRMux I__12212 (
            .O(N__51793),
            .I(N__51269));
    SRMux I__12211 (
            .O(N__51792),
            .I(N__51269));
    SRMux I__12210 (
            .O(N__51791),
            .I(N__51269));
    SRMux I__12209 (
            .O(N__51790),
            .I(N__51269));
    SRMux I__12208 (
            .O(N__51789),
            .I(N__51269));
    SRMux I__12207 (
            .O(N__51788),
            .I(N__51269));
    SRMux I__12206 (
            .O(N__51787),
            .I(N__51269));
    SRMux I__12205 (
            .O(N__51786),
            .I(N__51269));
    SRMux I__12204 (
            .O(N__51785),
            .I(N__51269));
    SRMux I__12203 (
            .O(N__51784),
            .I(N__51269));
    SRMux I__12202 (
            .O(N__51783),
            .I(N__51269));
    SRMux I__12201 (
            .O(N__51782),
            .I(N__51269));
    SRMux I__12200 (
            .O(N__51781),
            .I(N__51269));
    SRMux I__12199 (
            .O(N__51780),
            .I(N__51269));
    SRMux I__12198 (
            .O(N__51779),
            .I(N__51269));
    SRMux I__12197 (
            .O(N__51778),
            .I(N__51269));
    SRMux I__12196 (
            .O(N__51777),
            .I(N__51269));
    SRMux I__12195 (
            .O(N__51776),
            .I(N__51269));
    SRMux I__12194 (
            .O(N__51775),
            .I(N__51269));
    SRMux I__12193 (
            .O(N__51774),
            .I(N__51269));
    SRMux I__12192 (
            .O(N__51773),
            .I(N__51269));
    SRMux I__12191 (
            .O(N__51772),
            .I(N__51269));
    SRMux I__12190 (
            .O(N__51771),
            .I(N__51269));
    SRMux I__12189 (
            .O(N__51770),
            .I(N__51269));
    SRMux I__12188 (
            .O(N__51769),
            .I(N__51269));
    SRMux I__12187 (
            .O(N__51768),
            .I(N__51269));
    SRMux I__12186 (
            .O(N__51767),
            .I(N__51269));
    SRMux I__12185 (
            .O(N__51766),
            .I(N__51269));
    SRMux I__12184 (
            .O(N__51765),
            .I(N__51269));
    SRMux I__12183 (
            .O(N__51764),
            .I(N__51269));
    SRMux I__12182 (
            .O(N__51763),
            .I(N__51269));
    SRMux I__12181 (
            .O(N__51762),
            .I(N__51269));
    SRMux I__12180 (
            .O(N__51761),
            .I(N__51269));
    SRMux I__12179 (
            .O(N__51760),
            .I(N__51269));
    SRMux I__12178 (
            .O(N__51759),
            .I(N__51269));
    SRMux I__12177 (
            .O(N__51758),
            .I(N__51269));
    SRMux I__12176 (
            .O(N__51757),
            .I(N__51269));
    SRMux I__12175 (
            .O(N__51756),
            .I(N__51269));
    SRMux I__12174 (
            .O(N__51755),
            .I(N__51269));
    SRMux I__12173 (
            .O(N__51754),
            .I(N__51269));
    SRMux I__12172 (
            .O(N__51753),
            .I(N__51269));
    SRMux I__12171 (
            .O(N__51752),
            .I(N__51269));
    SRMux I__12170 (
            .O(N__51751),
            .I(N__51269));
    SRMux I__12169 (
            .O(N__51750),
            .I(N__51269));
    SRMux I__12168 (
            .O(N__51749),
            .I(N__51269));
    SRMux I__12167 (
            .O(N__51748),
            .I(N__51269));
    SRMux I__12166 (
            .O(N__51747),
            .I(N__51269));
    SRMux I__12165 (
            .O(N__51746),
            .I(N__51269));
    SRMux I__12164 (
            .O(N__51745),
            .I(N__51269));
    SRMux I__12163 (
            .O(N__51744),
            .I(N__51269));
    SRMux I__12162 (
            .O(N__51743),
            .I(N__51269));
    SRMux I__12161 (
            .O(N__51742),
            .I(N__51269));
    SRMux I__12160 (
            .O(N__51741),
            .I(N__51269));
    SRMux I__12159 (
            .O(N__51740),
            .I(N__51269));
    SRMux I__12158 (
            .O(N__51739),
            .I(N__51269));
    SRMux I__12157 (
            .O(N__51738),
            .I(N__51269));
    SRMux I__12156 (
            .O(N__51737),
            .I(N__51269));
    SRMux I__12155 (
            .O(N__51736),
            .I(N__51269));
    SRMux I__12154 (
            .O(N__51735),
            .I(N__51269));
    SRMux I__12153 (
            .O(N__51734),
            .I(N__51269));
    SRMux I__12152 (
            .O(N__51733),
            .I(N__51269));
    SRMux I__12151 (
            .O(N__51732),
            .I(N__51269));
    SRMux I__12150 (
            .O(N__51731),
            .I(N__51269));
    SRMux I__12149 (
            .O(N__51730),
            .I(N__51269));
    SRMux I__12148 (
            .O(N__51729),
            .I(N__51269));
    SRMux I__12147 (
            .O(N__51728),
            .I(N__51269));
    SRMux I__12146 (
            .O(N__51727),
            .I(N__51269));
    SRMux I__12145 (
            .O(N__51726),
            .I(N__51269));
    SRMux I__12144 (
            .O(N__51725),
            .I(N__51269));
    SRMux I__12143 (
            .O(N__51724),
            .I(N__51269));
    SRMux I__12142 (
            .O(N__51723),
            .I(N__51269));
    SRMux I__12141 (
            .O(N__51722),
            .I(N__51269));
    SRMux I__12140 (
            .O(N__51721),
            .I(N__51269));
    SRMux I__12139 (
            .O(N__51720),
            .I(N__51269));
    SRMux I__12138 (
            .O(N__51719),
            .I(N__51269));
    SRMux I__12137 (
            .O(N__51718),
            .I(N__51269));
    SRMux I__12136 (
            .O(N__51717),
            .I(N__51269));
    SRMux I__12135 (
            .O(N__51716),
            .I(N__51269));
    SRMux I__12134 (
            .O(N__51715),
            .I(N__51269));
    SRMux I__12133 (
            .O(N__51714),
            .I(N__51269));
    SRMux I__12132 (
            .O(N__51713),
            .I(N__51269));
    SRMux I__12131 (
            .O(N__51712),
            .I(N__51269));
    SRMux I__12130 (
            .O(N__51711),
            .I(N__51269));
    SRMux I__12129 (
            .O(N__51710),
            .I(N__51269));
    SRMux I__12128 (
            .O(N__51709),
            .I(N__51269));
    SRMux I__12127 (
            .O(N__51708),
            .I(N__51269));
    SRMux I__12126 (
            .O(N__51707),
            .I(N__51269));
    SRMux I__12125 (
            .O(N__51706),
            .I(N__51269));
    SRMux I__12124 (
            .O(N__51705),
            .I(N__51269));
    SRMux I__12123 (
            .O(N__51704),
            .I(N__51269));
    SRMux I__12122 (
            .O(N__51703),
            .I(N__51269));
    SRMux I__12121 (
            .O(N__51702),
            .I(N__51269));
    SRMux I__12120 (
            .O(N__51701),
            .I(N__51269));
    SRMux I__12119 (
            .O(N__51700),
            .I(N__51269));
    SRMux I__12118 (
            .O(N__51699),
            .I(N__51269));
    SRMux I__12117 (
            .O(N__51698),
            .I(N__51269));
    SRMux I__12116 (
            .O(N__51697),
            .I(N__51269));
    SRMux I__12115 (
            .O(N__51696),
            .I(N__51269));
    SRMux I__12114 (
            .O(N__51695),
            .I(N__51269));
    SRMux I__12113 (
            .O(N__51694),
            .I(N__51269));
    SRMux I__12112 (
            .O(N__51693),
            .I(N__51269));
    SRMux I__12111 (
            .O(N__51692),
            .I(N__51269));
    SRMux I__12110 (
            .O(N__51691),
            .I(N__51269));
    SRMux I__12109 (
            .O(N__51690),
            .I(N__51269));
    SRMux I__12108 (
            .O(N__51689),
            .I(N__51269));
    SRMux I__12107 (
            .O(N__51688),
            .I(N__51269));
    SRMux I__12106 (
            .O(N__51687),
            .I(N__51269));
    SRMux I__12105 (
            .O(N__51686),
            .I(N__51269));
    SRMux I__12104 (
            .O(N__51685),
            .I(N__51269));
    SRMux I__12103 (
            .O(N__51684),
            .I(N__51269));
    SRMux I__12102 (
            .O(N__51683),
            .I(N__51269));
    SRMux I__12101 (
            .O(N__51682),
            .I(N__51269));
    SRMux I__12100 (
            .O(N__51681),
            .I(N__51269));
    SRMux I__12099 (
            .O(N__51680),
            .I(N__51269));
    SRMux I__12098 (
            .O(N__51679),
            .I(N__51269));
    SRMux I__12097 (
            .O(N__51678),
            .I(N__51269));
    SRMux I__12096 (
            .O(N__51677),
            .I(N__51269));
    SRMux I__12095 (
            .O(N__51676),
            .I(N__51269));
    SRMux I__12094 (
            .O(N__51675),
            .I(N__51269));
    SRMux I__12093 (
            .O(N__51674),
            .I(N__51269));
    SRMux I__12092 (
            .O(N__51673),
            .I(N__51269));
    SRMux I__12091 (
            .O(N__51672),
            .I(N__51269));
    SRMux I__12090 (
            .O(N__51671),
            .I(N__51269));
    SRMux I__12089 (
            .O(N__51670),
            .I(N__51269));
    SRMux I__12088 (
            .O(N__51669),
            .I(N__51269));
    SRMux I__12087 (
            .O(N__51668),
            .I(N__51269));
    SRMux I__12086 (
            .O(N__51667),
            .I(N__51269));
    SRMux I__12085 (
            .O(N__51666),
            .I(N__51269));
    SRMux I__12084 (
            .O(N__51665),
            .I(N__51269));
    SRMux I__12083 (
            .O(N__51664),
            .I(N__51269));
    SRMux I__12082 (
            .O(N__51663),
            .I(N__51269));
    SRMux I__12081 (
            .O(N__51662),
            .I(N__51269));
    SRMux I__12080 (
            .O(N__51661),
            .I(N__51269));
    SRMux I__12079 (
            .O(N__51660),
            .I(N__51269));
    SRMux I__12078 (
            .O(N__51659),
            .I(N__51269));
    SRMux I__12077 (
            .O(N__51658),
            .I(N__51269));
    SRMux I__12076 (
            .O(N__51657),
            .I(N__51269));
    SRMux I__12075 (
            .O(N__51656),
            .I(N__51269));
    SRMux I__12074 (
            .O(N__51655),
            .I(N__51269));
    SRMux I__12073 (
            .O(N__51654),
            .I(N__51269));
    SRMux I__12072 (
            .O(N__51653),
            .I(N__51269));
    SRMux I__12071 (
            .O(N__51652),
            .I(N__51269));
    SRMux I__12070 (
            .O(N__51651),
            .I(N__51269));
    SRMux I__12069 (
            .O(N__51650),
            .I(N__51269));
    SRMux I__12068 (
            .O(N__51649),
            .I(N__51269));
    SRMux I__12067 (
            .O(N__51648),
            .I(N__51269));
    SRMux I__12066 (
            .O(N__51647),
            .I(N__51269));
    SRMux I__12065 (
            .O(N__51646),
            .I(N__51269));
    SRMux I__12064 (
            .O(N__51645),
            .I(N__51269));
    SRMux I__12063 (
            .O(N__51644),
            .I(N__51269));
    SRMux I__12062 (
            .O(N__51643),
            .I(N__51269));
    SRMux I__12061 (
            .O(N__51642),
            .I(N__51269));
    GlobalMux I__12060 (
            .O(N__51269),
            .I(N__51266));
    gio2CtrlBuf I__12059 (
            .O(N__51266),
            .I(LED3_c_i_g));
    InMux I__12058 (
            .O(N__51263),
            .I(N__51259));
    InMux I__12057 (
            .O(N__51262),
            .I(N__51256));
    LocalMux I__12056 (
            .O(N__51259),
            .I(N__51253));
    LocalMux I__12055 (
            .O(N__51256),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4 ));
    Odrv4 I__12054 (
            .O(N__51253),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4 ));
    InMux I__12053 (
            .O(N__51248),
            .I(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3 ));
    InMux I__12052 (
            .O(N__51245),
            .I(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4 ));
    InMux I__12051 (
            .O(N__51242),
            .I(N__51238));
    InMux I__12050 (
            .O(N__51241),
            .I(N__51235));
    LocalMux I__12049 (
            .O(N__51238),
            .I(N__51232));
    LocalMux I__12048 (
            .O(N__51235),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5 ));
    Odrv4 I__12047 (
            .O(N__51232),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5 ));
    InMux I__12046 (
            .O(N__51227),
            .I(N__51224));
    LocalMux I__12045 (
            .O(N__51224),
            .I(N__51220));
    InMux I__12044 (
            .O(N__51223),
            .I(N__51217));
    Span4Mux_v I__12043 (
            .O(N__51220),
            .I(N__51208));
    LocalMux I__12042 (
            .O(N__51217),
            .I(N__51208));
    InMux I__12041 (
            .O(N__51216),
            .I(N__51205));
    InMux I__12040 (
            .O(N__51215),
            .I(N__51198));
    InMux I__12039 (
            .O(N__51214),
            .I(N__51198));
    InMux I__12038 (
            .O(N__51213),
            .I(N__51198));
    Span4Mux_v I__12037 (
            .O(N__51208),
            .I(N__51192));
    LocalMux I__12036 (
            .O(N__51205),
            .I(N__51192));
    LocalMux I__12035 (
            .O(N__51198),
            .I(N__51188));
    InMux I__12034 (
            .O(N__51197),
            .I(N__51185));
    Span4Mux_h I__12033 (
            .O(N__51192),
            .I(N__51182));
    InMux I__12032 (
            .O(N__51191),
            .I(N__51179));
    Span4Mux_v I__12031 (
            .O(N__51188),
            .I(N__51175));
    LocalMux I__12030 (
            .O(N__51185),
            .I(N__51172));
    Span4Mux_h I__12029 (
            .O(N__51182),
            .I(N__51169));
    LocalMux I__12028 (
            .O(N__51179),
            .I(N__51166));
    InMux I__12027 (
            .O(N__51178),
            .I(N__51163));
    Span4Mux_v I__12026 (
            .O(N__51175),
            .I(N__51158));
    Span4Mux_v I__12025 (
            .O(N__51172),
            .I(N__51158));
    Span4Mux_h I__12024 (
            .O(N__51169),
            .I(N__51151));
    Span4Mux_v I__12023 (
            .O(N__51166),
            .I(N__51151));
    LocalMux I__12022 (
            .O(N__51163),
            .I(N__51151));
    Odrv4 I__12021 (
            .O(N__51158),
            .I(\spi_slave_inst.spi_csZ0 ));
    Odrv4 I__12020 (
            .O(N__51151),
            .I(\spi_slave_inst.spi_csZ0 ));
    InMux I__12019 (
            .O(N__51146),
            .I(N__51138));
    InMux I__12018 (
            .O(N__51145),
            .I(N__51138));
    InMux I__12017 (
            .O(N__51144),
            .I(N__51133));
    InMux I__12016 (
            .O(N__51143),
            .I(N__51133));
    LocalMux I__12015 (
            .O(N__51138),
            .I(N__51128));
    LocalMux I__12014 (
            .O(N__51133),
            .I(N__51128));
    Odrv4 I__12013 (
            .O(N__51128),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_i6 ));
    InMux I__12012 (
            .O(N__51125),
            .I(N__51121));
    InMux I__12011 (
            .O(N__51124),
            .I(N__51118));
    LocalMux I__12010 (
            .O(N__51121),
            .I(\spi_slave_inst.tx_done_neg_sclk_iZ0 ));
    LocalMux I__12009 (
            .O(N__51118),
            .I(\spi_slave_inst.tx_done_neg_sclk_iZ0 ));
    InMux I__12008 (
            .O(N__51113),
            .I(N__51110));
    LocalMux I__12007 (
            .O(N__51110),
            .I(\spi_slave_inst.tx_done_reg1_iZ0 ));
    InMux I__12006 (
            .O(N__51107),
            .I(N__51104));
    LocalMux I__12005 (
            .O(N__51104),
            .I(\spi_slave_inst.tx_done_reg3_iZ0 ));
    InMux I__12004 (
            .O(N__51101),
            .I(N__51097));
    InMux I__12003 (
            .O(N__51100),
            .I(N__51094));
    LocalMux I__12002 (
            .O(N__51097),
            .I(\spi_slave_inst.tx_done_reg2_iZ0 ));
    LocalMux I__12001 (
            .O(N__51094),
            .I(\spi_slave_inst.tx_done_reg2_iZ0 ));
    InMux I__12000 (
            .O(N__51089),
            .I(N__51086));
    LocalMux I__11999 (
            .O(N__51086),
            .I(N__51083));
    Span4Mux_h I__11998 (
            .O(N__51083),
            .I(N__51080));
    Odrv4 I__11997 (
            .O(N__51080),
            .I(\spi_slave_inst.un4_tx_done_reg2_i ));
    InMux I__11996 (
            .O(N__51077),
            .I(N__51071));
    InMux I__11995 (
            .O(N__51076),
            .I(N__51065));
    InMux I__11994 (
            .O(N__51075),
            .I(N__51059));
    InMux I__11993 (
            .O(N__51074),
            .I(N__51056));
    LocalMux I__11992 (
            .O(N__51071),
            .I(N__51047));
    InMux I__11991 (
            .O(N__51070),
            .I(N__51044));
    InMux I__11990 (
            .O(N__51069),
            .I(N__51034));
    InMux I__11989 (
            .O(N__51068),
            .I(N__51031));
    LocalMux I__11988 (
            .O(N__51065),
            .I(N__51026));
    InMux I__11987 (
            .O(N__51064),
            .I(N__51023));
    InMux I__11986 (
            .O(N__51063),
            .I(N__51020));
    InMux I__11985 (
            .O(N__51062),
            .I(N__51014));
    LocalMux I__11984 (
            .O(N__51059),
            .I(N__51009));
    LocalMux I__11983 (
            .O(N__51056),
            .I(N__51009));
    InMux I__11982 (
            .O(N__51055),
            .I(N__51006));
    InMux I__11981 (
            .O(N__51054),
            .I(N__51003));
    InMux I__11980 (
            .O(N__51053),
            .I(N__51000));
    InMux I__11979 (
            .O(N__51052),
            .I(N__50997));
    InMux I__11978 (
            .O(N__51051),
            .I(N__50994));
    InMux I__11977 (
            .O(N__51050),
            .I(N__50991));
    Span4Mux_h I__11976 (
            .O(N__51047),
            .I(N__50986));
    LocalMux I__11975 (
            .O(N__51044),
            .I(N__50986));
    InMux I__11974 (
            .O(N__51043),
            .I(N__50979));
    InMux I__11973 (
            .O(N__51042),
            .I(N__50976));
    InMux I__11972 (
            .O(N__51041),
            .I(N__50973));
    InMux I__11971 (
            .O(N__51040),
            .I(N__50970));
    InMux I__11970 (
            .O(N__51039),
            .I(N__50967));
    InMux I__11969 (
            .O(N__51038),
            .I(N__50964));
    InMux I__11968 (
            .O(N__51037),
            .I(N__50961));
    LocalMux I__11967 (
            .O(N__51034),
            .I(N__50956));
    LocalMux I__11966 (
            .O(N__51031),
            .I(N__50956));
    InMux I__11965 (
            .O(N__51030),
            .I(N__50953));
    InMux I__11964 (
            .O(N__51029),
            .I(N__50950));
    Span4Mux_v I__11963 (
            .O(N__51026),
            .I(N__50943));
    LocalMux I__11962 (
            .O(N__51023),
            .I(N__50943));
    LocalMux I__11961 (
            .O(N__51020),
            .I(N__50943));
    InMux I__11960 (
            .O(N__51019),
            .I(N__50940));
    InMux I__11959 (
            .O(N__51018),
            .I(N__50935));
    InMux I__11958 (
            .O(N__51017),
            .I(N__50932));
    LocalMux I__11957 (
            .O(N__51014),
            .I(N__50925));
    Span4Mux_h I__11956 (
            .O(N__51009),
            .I(N__50914));
    LocalMux I__11955 (
            .O(N__51006),
            .I(N__50914));
    LocalMux I__11954 (
            .O(N__51003),
            .I(N__50914));
    LocalMux I__11953 (
            .O(N__51000),
            .I(N__50914));
    LocalMux I__11952 (
            .O(N__50997),
            .I(N__50914));
    LocalMux I__11951 (
            .O(N__50994),
            .I(N__50907));
    LocalMux I__11950 (
            .O(N__50991),
            .I(N__50907));
    Span4Mux_v I__11949 (
            .O(N__50986),
            .I(N__50907));
    InMux I__11948 (
            .O(N__50985),
            .I(N__50904));
    InMux I__11947 (
            .O(N__50984),
            .I(N__50900));
    InMux I__11946 (
            .O(N__50983),
            .I(N__50893));
    InMux I__11945 (
            .O(N__50982),
            .I(N__50889));
    LocalMux I__11944 (
            .O(N__50979),
            .I(N__50884));
    LocalMux I__11943 (
            .O(N__50976),
            .I(N__50884));
    LocalMux I__11942 (
            .O(N__50973),
            .I(N__50872));
    LocalMux I__11941 (
            .O(N__50970),
            .I(N__50872));
    LocalMux I__11940 (
            .O(N__50967),
            .I(N__50861));
    LocalMux I__11939 (
            .O(N__50964),
            .I(N__50861));
    LocalMux I__11938 (
            .O(N__50961),
            .I(N__50861));
    Span4Mux_h I__11937 (
            .O(N__50956),
            .I(N__50861));
    LocalMux I__11936 (
            .O(N__50953),
            .I(N__50861));
    LocalMux I__11935 (
            .O(N__50950),
            .I(N__50858));
    Span4Mux_h I__11934 (
            .O(N__50943),
            .I(N__50855));
    LocalMux I__11933 (
            .O(N__50940),
            .I(N__50852));
    InMux I__11932 (
            .O(N__50939),
            .I(N__50848));
    InMux I__11931 (
            .O(N__50938),
            .I(N__50845));
    LocalMux I__11930 (
            .O(N__50935),
            .I(N__50840));
    LocalMux I__11929 (
            .O(N__50932),
            .I(N__50840));
    InMux I__11928 (
            .O(N__50931),
            .I(N__50837));
    InMux I__11927 (
            .O(N__50930),
            .I(N__50834));
    InMux I__11926 (
            .O(N__50929),
            .I(N__50831));
    InMux I__11925 (
            .O(N__50928),
            .I(N__50828));
    Span4Mux_v I__11924 (
            .O(N__50925),
            .I(N__50825));
    Span4Mux_v I__11923 (
            .O(N__50914),
            .I(N__50820));
    Span4Mux_h I__11922 (
            .O(N__50907),
            .I(N__50820));
    LocalMux I__11921 (
            .O(N__50904),
            .I(N__50817));
    InMux I__11920 (
            .O(N__50903),
            .I(N__50811));
    LocalMux I__11919 (
            .O(N__50900),
            .I(N__50808));
    InMux I__11918 (
            .O(N__50899),
            .I(N__50805));
    InMux I__11917 (
            .O(N__50898),
            .I(N__50802));
    InMux I__11916 (
            .O(N__50897),
            .I(N__50799));
    InMux I__11915 (
            .O(N__50896),
            .I(N__50796));
    LocalMux I__11914 (
            .O(N__50893),
            .I(N__50793));
    InMux I__11913 (
            .O(N__50892),
            .I(N__50790));
    LocalMux I__11912 (
            .O(N__50889),
            .I(N__50787));
    Span4Mux_v I__11911 (
            .O(N__50884),
            .I(N__50784));
    InMux I__11910 (
            .O(N__50883),
            .I(N__50781));
    InMux I__11909 (
            .O(N__50882),
            .I(N__50778));
    InMux I__11908 (
            .O(N__50881),
            .I(N__50775));
    InMux I__11907 (
            .O(N__50880),
            .I(N__50772));
    InMux I__11906 (
            .O(N__50879),
            .I(N__50769));
    InMux I__11905 (
            .O(N__50878),
            .I(N__50766));
    InMux I__11904 (
            .O(N__50877),
            .I(N__50763));
    Span4Mux_v I__11903 (
            .O(N__50872),
            .I(N__50758));
    Span4Mux_v I__11902 (
            .O(N__50861),
            .I(N__50758));
    Span4Mux_v I__11901 (
            .O(N__50858),
            .I(N__50755));
    Span4Mux_v I__11900 (
            .O(N__50855),
            .I(N__50750));
    Span4Mux_v I__11899 (
            .O(N__50852),
            .I(N__50750));
    InMux I__11898 (
            .O(N__50851),
            .I(N__50747));
    LocalMux I__11897 (
            .O(N__50848),
            .I(N__50742));
    LocalMux I__11896 (
            .O(N__50845),
            .I(N__50742));
    Span4Mux_v I__11895 (
            .O(N__50840),
            .I(N__50739));
    LocalMux I__11894 (
            .O(N__50837),
            .I(N__50724));
    LocalMux I__11893 (
            .O(N__50834),
            .I(N__50724));
    LocalMux I__11892 (
            .O(N__50831),
            .I(N__50724));
    LocalMux I__11891 (
            .O(N__50828),
            .I(N__50724));
    Span4Mux_v I__11890 (
            .O(N__50825),
            .I(N__50724));
    Span4Mux_h I__11889 (
            .O(N__50820),
            .I(N__50724));
    Span4Mux_h I__11888 (
            .O(N__50817),
            .I(N__50724));
    InMux I__11887 (
            .O(N__50816),
            .I(N__50719));
    InMux I__11886 (
            .O(N__50815),
            .I(N__50719));
    InMux I__11885 (
            .O(N__50814),
            .I(N__50712));
    LocalMux I__11884 (
            .O(N__50811),
            .I(N__50707));
    Span4Mux_v I__11883 (
            .O(N__50808),
            .I(N__50707));
    LocalMux I__11882 (
            .O(N__50805),
            .I(N__50696));
    LocalMux I__11881 (
            .O(N__50802),
            .I(N__50696));
    LocalMux I__11880 (
            .O(N__50799),
            .I(N__50696));
    LocalMux I__11879 (
            .O(N__50796),
            .I(N__50696));
    Span4Mux_v I__11878 (
            .O(N__50793),
            .I(N__50696));
    LocalMux I__11877 (
            .O(N__50790),
            .I(N__50689));
    Span4Mux_v I__11876 (
            .O(N__50787),
            .I(N__50689));
    Span4Mux_h I__11875 (
            .O(N__50784),
            .I(N__50689));
    LocalMux I__11874 (
            .O(N__50781),
            .I(N__50682));
    LocalMux I__11873 (
            .O(N__50778),
            .I(N__50682));
    LocalMux I__11872 (
            .O(N__50775),
            .I(N__50682));
    LocalMux I__11871 (
            .O(N__50772),
            .I(N__50667));
    LocalMux I__11870 (
            .O(N__50769),
            .I(N__50667));
    LocalMux I__11869 (
            .O(N__50766),
            .I(N__50667));
    LocalMux I__11868 (
            .O(N__50763),
            .I(N__50667));
    Sp12to4 I__11867 (
            .O(N__50758),
            .I(N__50667));
    Sp12to4 I__11866 (
            .O(N__50755),
            .I(N__50667));
    Sp12to4 I__11865 (
            .O(N__50750),
            .I(N__50667));
    LocalMux I__11864 (
            .O(N__50747),
            .I(N__50664));
    Span4Mux_v I__11863 (
            .O(N__50742),
            .I(N__50655));
    Span4Mux_v I__11862 (
            .O(N__50739),
            .I(N__50655));
    Span4Mux_v I__11861 (
            .O(N__50724),
            .I(N__50655));
    LocalMux I__11860 (
            .O(N__50719),
            .I(N__50655));
    InMux I__11859 (
            .O(N__50718),
            .I(N__50652));
    InMux I__11858 (
            .O(N__50717),
            .I(N__50649));
    InMux I__11857 (
            .O(N__50716),
            .I(N__50646));
    InMux I__11856 (
            .O(N__50715),
            .I(N__50643));
    LocalMux I__11855 (
            .O(N__50712),
            .I(N__50634));
    Span4Mux_v I__11854 (
            .O(N__50707),
            .I(N__50634));
    Span4Mux_v I__11853 (
            .O(N__50696),
            .I(N__50634));
    Span4Mux_h I__11852 (
            .O(N__50689),
            .I(N__50634));
    Span12Mux_v I__11851 (
            .O(N__50682),
            .I(N__50629));
    Span12Mux_h I__11850 (
            .O(N__50667),
            .I(N__50629));
    Span4Mux_v I__11849 (
            .O(N__50664),
            .I(N__50624));
    Span4Mux_h I__11848 (
            .O(N__50655),
            .I(N__50624));
    LocalMux I__11847 (
            .O(N__50652),
            .I(spi_data_mosi_1));
    LocalMux I__11846 (
            .O(N__50649),
            .I(spi_data_mosi_1));
    LocalMux I__11845 (
            .O(N__50646),
            .I(spi_data_mosi_1));
    LocalMux I__11844 (
            .O(N__50643),
            .I(spi_data_mosi_1));
    Odrv4 I__11843 (
            .O(N__50634),
            .I(spi_data_mosi_1));
    Odrv12 I__11842 (
            .O(N__50629),
            .I(spi_data_mosi_1));
    Odrv4 I__11841 (
            .O(N__50624),
            .I(spi_data_mosi_1));
    InMux I__11840 (
            .O(N__50609),
            .I(N__50606));
    LocalMux I__11839 (
            .O(N__50606),
            .I(N__50603));
    Span4Mux_h I__11838 (
            .O(N__50603),
            .I(N__50600));
    Span4Mux_h I__11837 (
            .O(N__50600),
            .I(N__50597));
    Odrv4 I__11836 (
            .O(N__50597),
            .I(sDAC_mem_25Z0Z_1));
    CEMux I__11835 (
            .O(N__50594),
            .I(N__50590));
    CEMux I__11834 (
            .O(N__50593),
            .I(N__50587));
    LocalMux I__11833 (
            .O(N__50590),
            .I(N__50584));
    LocalMux I__11832 (
            .O(N__50587),
            .I(N__50581));
    Span4Mux_v I__11831 (
            .O(N__50584),
            .I(N__50578));
    Span4Mux_v I__11830 (
            .O(N__50581),
            .I(N__50575));
    Odrv4 I__11829 (
            .O(N__50578),
            .I(sDAC_mem_25_1_sqmuxa));
    Odrv4 I__11828 (
            .O(N__50575),
            .I(sDAC_mem_25_1_sqmuxa));
    InMux I__11827 (
            .O(N__50570),
            .I(N__50567));
    LocalMux I__11826 (
            .O(N__50567),
            .I(N__50564));
    Span4Mux_h I__11825 (
            .O(N__50564),
            .I(N__50561));
    Odrv4 I__11824 (
            .O(N__50561),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_7 ));
    InMux I__11823 (
            .O(N__50558),
            .I(N__50555));
    LocalMux I__11822 (
            .O(N__50555),
            .I(N__50552));
    Span4Mux_v I__11821 (
            .O(N__50552),
            .I(N__50549));
    Odrv4 I__11820 (
            .O(N__50549),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_7 ));
    InMux I__11819 (
            .O(N__50546),
            .I(N__50538));
    InMux I__11818 (
            .O(N__50545),
            .I(N__50535));
    InMux I__11817 (
            .O(N__50544),
            .I(N__50532));
    InMux I__11816 (
            .O(N__50543),
            .I(N__50523));
    InMux I__11815 (
            .O(N__50542),
            .I(N__50520));
    InMux I__11814 (
            .O(N__50541),
            .I(N__50517));
    LocalMux I__11813 (
            .O(N__50538),
            .I(N__50513));
    LocalMux I__11812 (
            .O(N__50535),
            .I(N__50508));
    LocalMux I__11811 (
            .O(N__50532),
            .I(N__50508));
    InMux I__11810 (
            .O(N__50531),
            .I(N__50505));
    InMux I__11809 (
            .O(N__50530),
            .I(N__50502));
    InMux I__11808 (
            .O(N__50529),
            .I(N__50499));
    InMux I__11807 (
            .O(N__50528),
            .I(N__50496));
    InMux I__11806 (
            .O(N__50527),
            .I(N__50492));
    InMux I__11805 (
            .O(N__50526),
            .I(N__50489));
    LocalMux I__11804 (
            .O(N__50523),
            .I(N__50473));
    LocalMux I__11803 (
            .O(N__50520),
            .I(N__50473));
    LocalMux I__11802 (
            .O(N__50517),
            .I(N__50473));
    InMux I__11801 (
            .O(N__50516),
            .I(N__50470));
    Span4Mux_h I__11800 (
            .O(N__50513),
            .I(N__50452));
    Span4Mux_v I__11799 (
            .O(N__50508),
            .I(N__50452));
    LocalMux I__11798 (
            .O(N__50505),
            .I(N__50452));
    LocalMux I__11797 (
            .O(N__50502),
            .I(N__50452));
    LocalMux I__11796 (
            .O(N__50499),
            .I(N__50452));
    LocalMux I__11795 (
            .O(N__50496),
            .I(N__50449));
    InMux I__11794 (
            .O(N__50495),
            .I(N__50446));
    LocalMux I__11793 (
            .O(N__50492),
            .I(N__50443));
    LocalMux I__11792 (
            .O(N__50489),
            .I(N__50440));
    InMux I__11791 (
            .O(N__50488),
            .I(N__50437));
    InMux I__11790 (
            .O(N__50487),
            .I(N__50434));
    InMux I__11789 (
            .O(N__50486),
            .I(N__50431));
    InMux I__11788 (
            .O(N__50485),
            .I(N__50427));
    InMux I__11787 (
            .O(N__50484),
            .I(N__50424));
    InMux I__11786 (
            .O(N__50483),
            .I(N__50421));
    InMux I__11785 (
            .O(N__50482),
            .I(N__50417));
    InMux I__11784 (
            .O(N__50481),
            .I(N__50414));
    InMux I__11783 (
            .O(N__50480),
            .I(N__50410));
    Span4Mux_v I__11782 (
            .O(N__50473),
            .I(N__50402));
    LocalMux I__11781 (
            .O(N__50470),
            .I(N__50402));
    InMux I__11780 (
            .O(N__50469),
            .I(N__50399));
    InMux I__11779 (
            .O(N__50468),
            .I(N__50396));
    InMux I__11778 (
            .O(N__50467),
            .I(N__50393));
    InMux I__11777 (
            .O(N__50466),
            .I(N__50388));
    InMux I__11776 (
            .O(N__50465),
            .I(N__50385));
    InMux I__11775 (
            .O(N__50464),
            .I(N__50382));
    InMux I__11774 (
            .O(N__50463),
            .I(N__50375));
    Span4Mux_h I__11773 (
            .O(N__50452),
            .I(N__50367));
    Span4Mux_v I__11772 (
            .O(N__50449),
            .I(N__50367));
    LocalMux I__11771 (
            .O(N__50446),
            .I(N__50367));
    Span4Mux_v I__11770 (
            .O(N__50443),
            .I(N__50356));
    Span4Mux_h I__11769 (
            .O(N__50440),
            .I(N__50356));
    LocalMux I__11768 (
            .O(N__50437),
            .I(N__50356));
    LocalMux I__11767 (
            .O(N__50434),
            .I(N__50356));
    LocalMux I__11766 (
            .O(N__50431),
            .I(N__50356));
    InMux I__11765 (
            .O(N__50430),
            .I(N__50353));
    LocalMux I__11764 (
            .O(N__50427),
            .I(N__50346));
    LocalMux I__11763 (
            .O(N__50424),
            .I(N__50346));
    LocalMux I__11762 (
            .O(N__50421),
            .I(N__50346));
    InMux I__11761 (
            .O(N__50420),
            .I(N__50343));
    LocalMux I__11760 (
            .O(N__50417),
            .I(N__50338));
    LocalMux I__11759 (
            .O(N__50414),
            .I(N__50338));
    InMux I__11758 (
            .O(N__50413),
            .I(N__50335));
    LocalMux I__11757 (
            .O(N__50410),
            .I(N__50331));
    InMux I__11756 (
            .O(N__50409),
            .I(N__50324));
    InMux I__11755 (
            .O(N__50408),
            .I(N__50321));
    InMux I__11754 (
            .O(N__50407),
            .I(N__50318));
    Span4Mux_v I__11753 (
            .O(N__50402),
            .I(N__50310));
    LocalMux I__11752 (
            .O(N__50399),
            .I(N__50310));
    LocalMux I__11751 (
            .O(N__50396),
            .I(N__50310));
    LocalMux I__11750 (
            .O(N__50393),
            .I(N__50302));
    InMux I__11749 (
            .O(N__50392),
            .I(N__50299));
    InMux I__11748 (
            .O(N__50391),
            .I(N__50296));
    LocalMux I__11747 (
            .O(N__50388),
            .I(N__50289));
    LocalMux I__11746 (
            .O(N__50385),
            .I(N__50289));
    LocalMux I__11745 (
            .O(N__50382),
            .I(N__50289));
    InMux I__11744 (
            .O(N__50381),
            .I(N__50286));
    InMux I__11743 (
            .O(N__50380),
            .I(N__50283));
    InMux I__11742 (
            .O(N__50379),
            .I(N__50280));
    InMux I__11741 (
            .O(N__50378),
            .I(N__50277));
    LocalMux I__11740 (
            .O(N__50375),
            .I(N__50274));
    InMux I__11739 (
            .O(N__50374),
            .I(N__50271));
    Span4Mux_v I__11738 (
            .O(N__50367),
            .I(N__50268));
    Span4Mux_v I__11737 (
            .O(N__50356),
            .I(N__50261));
    LocalMux I__11736 (
            .O(N__50353),
            .I(N__50261));
    Span4Mux_v I__11735 (
            .O(N__50346),
            .I(N__50261));
    LocalMux I__11734 (
            .O(N__50343),
            .I(N__50254));
    Span4Mux_v I__11733 (
            .O(N__50338),
            .I(N__50254));
    LocalMux I__11732 (
            .O(N__50335),
            .I(N__50254));
    InMux I__11731 (
            .O(N__50334),
            .I(N__50251));
    Span12Mux_v I__11730 (
            .O(N__50331),
            .I(N__50248));
    InMux I__11729 (
            .O(N__50330),
            .I(N__50245));
    InMux I__11728 (
            .O(N__50329),
            .I(N__50242));
    InMux I__11727 (
            .O(N__50328),
            .I(N__50239));
    InMux I__11726 (
            .O(N__50327),
            .I(N__50236));
    LocalMux I__11725 (
            .O(N__50324),
            .I(N__50229));
    LocalMux I__11724 (
            .O(N__50321),
            .I(N__50229));
    LocalMux I__11723 (
            .O(N__50318),
            .I(N__50229));
    InMux I__11722 (
            .O(N__50317),
            .I(N__50226));
    Span4Mux_v I__11721 (
            .O(N__50310),
            .I(N__50221));
    InMux I__11720 (
            .O(N__50309),
            .I(N__50218));
    InMux I__11719 (
            .O(N__50308),
            .I(N__50215));
    InMux I__11718 (
            .O(N__50307),
            .I(N__50212));
    InMux I__11717 (
            .O(N__50306),
            .I(N__50209));
    InMux I__11716 (
            .O(N__50305),
            .I(N__50206));
    Span12Mux_s9_v I__11715 (
            .O(N__50302),
            .I(N__50199));
    LocalMux I__11714 (
            .O(N__50299),
            .I(N__50199));
    LocalMux I__11713 (
            .O(N__50296),
            .I(N__50199));
    Span4Mux_v I__11712 (
            .O(N__50289),
            .I(N__50196));
    LocalMux I__11711 (
            .O(N__50286),
            .I(N__50189));
    LocalMux I__11710 (
            .O(N__50283),
            .I(N__50189));
    LocalMux I__11709 (
            .O(N__50280),
            .I(N__50189));
    LocalMux I__11708 (
            .O(N__50277),
            .I(N__50186));
    Span4Mux_v I__11707 (
            .O(N__50274),
            .I(N__50183));
    LocalMux I__11706 (
            .O(N__50271),
            .I(N__50180));
    Span4Mux_v I__11705 (
            .O(N__50268),
            .I(N__50171));
    Span4Mux_h I__11704 (
            .O(N__50261),
            .I(N__50171));
    Span4Mux_v I__11703 (
            .O(N__50254),
            .I(N__50171));
    LocalMux I__11702 (
            .O(N__50251),
            .I(N__50171));
    Span12Mux_h I__11701 (
            .O(N__50248),
            .I(N__50161));
    LocalMux I__11700 (
            .O(N__50245),
            .I(N__50161));
    LocalMux I__11699 (
            .O(N__50242),
            .I(N__50161));
    LocalMux I__11698 (
            .O(N__50239),
            .I(N__50156));
    LocalMux I__11697 (
            .O(N__50236),
            .I(N__50156));
    Span4Mux_v I__11696 (
            .O(N__50229),
            .I(N__50153));
    LocalMux I__11695 (
            .O(N__50226),
            .I(N__50150));
    InMux I__11694 (
            .O(N__50225),
            .I(N__50147));
    InMux I__11693 (
            .O(N__50224),
            .I(N__50144));
    Span4Mux_h I__11692 (
            .O(N__50221),
            .I(N__50131));
    LocalMux I__11691 (
            .O(N__50218),
            .I(N__50131));
    LocalMux I__11690 (
            .O(N__50215),
            .I(N__50131));
    LocalMux I__11689 (
            .O(N__50212),
            .I(N__50131));
    LocalMux I__11688 (
            .O(N__50209),
            .I(N__50131));
    LocalMux I__11687 (
            .O(N__50206),
            .I(N__50131));
    Span12Mux_v I__11686 (
            .O(N__50199),
            .I(N__50128));
    Sp12to4 I__11685 (
            .O(N__50196),
            .I(N__50117));
    Span12Mux_v I__11684 (
            .O(N__50189),
            .I(N__50117));
    Span12Mux_v I__11683 (
            .O(N__50186),
            .I(N__50117));
    Sp12to4 I__11682 (
            .O(N__50183),
            .I(N__50117));
    Span12Mux_s10_h I__11681 (
            .O(N__50180),
            .I(N__50117));
    Span4Mux_h I__11680 (
            .O(N__50171),
            .I(N__50114));
    InMux I__11679 (
            .O(N__50170),
            .I(N__50111));
    InMux I__11678 (
            .O(N__50169),
            .I(N__50108));
    InMux I__11677 (
            .O(N__50168),
            .I(N__50105));
    Span12Mux_v I__11676 (
            .O(N__50161),
            .I(N__50100));
    Span12Mux_s11_h I__11675 (
            .O(N__50156),
            .I(N__50100));
    Span4Mux_h I__11674 (
            .O(N__50153),
            .I(N__50089));
    Span4Mux_v I__11673 (
            .O(N__50150),
            .I(N__50089));
    LocalMux I__11672 (
            .O(N__50147),
            .I(N__50089));
    LocalMux I__11671 (
            .O(N__50144),
            .I(N__50089));
    Span4Mux_v I__11670 (
            .O(N__50131),
            .I(N__50089));
    Odrv12 I__11669 (
            .O(N__50128),
            .I(spi_data_mosi_6));
    Odrv12 I__11668 (
            .O(N__50117),
            .I(spi_data_mosi_6));
    Odrv4 I__11667 (
            .O(N__50114),
            .I(spi_data_mosi_6));
    LocalMux I__11666 (
            .O(N__50111),
            .I(spi_data_mosi_6));
    LocalMux I__11665 (
            .O(N__50108),
            .I(spi_data_mosi_6));
    LocalMux I__11664 (
            .O(N__50105),
            .I(spi_data_mosi_6));
    Odrv12 I__11663 (
            .O(N__50100),
            .I(spi_data_mosi_6));
    Odrv4 I__11662 (
            .O(N__50089),
            .I(spi_data_mosi_6));
    InMux I__11661 (
            .O(N__50072),
            .I(N__50069));
    LocalMux I__11660 (
            .O(N__50069),
            .I(N__50066));
    Odrv4 I__11659 (
            .O(N__50066),
            .I(sEEADC_freqZ0Z_6));
    InMux I__11658 (
            .O(N__50063),
            .I(N__50044));
    InMux I__11657 (
            .O(N__50062),
            .I(N__50041));
    InMux I__11656 (
            .O(N__50061),
            .I(N__50038));
    InMux I__11655 (
            .O(N__50060),
            .I(N__50024));
    InMux I__11654 (
            .O(N__50059),
            .I(N__50020));
    InMux I__11653 (
            .O(N__50058),
            .I(N__50017));
    InMux I__11652 (
            .O(N__50057),
            .I(N__50013));
    InMux I__11651 (
            .O(N__50056),
            .I(N__50010));
    InMux I__11650 (
            .O(N__50055),
            .I(N__50006));
    InMux I__11649 (
            .O(N__50054),
            .I(N__50003));
    InMux I__11648 (
            .O(N__50053),
            .I(N__50000));
    InMux I__11647 (
            .O(N__50052),
            .I(N__49997));
    InMux I__11646 (
            .O(N__50051),
            .I(N__49991));
    InMux I__11645 (
            .O(N__50050),
            .I(N__49987));
    InMux I__11644 (
            .O(N__50049),
            .I(N__49984));
    InMux I__11643 (
            .O(N__50048),
            .I(N__49981));
    InMux I__11642 (
            .O(N__50047),
            .I(N__49978));
    LocalMux I__11641 (
            .O(N__50044),
            .I(N__49973));
    LocalMux I__11640 (
            .O(N__50041),
            .I(N__49973));
    LocalMux I__11639 (
            .O(N__50038),
            .I(N__49970));
    InMux I__11638 (
            .O(N__50037),
            .I(N__49967));
    InMux I__11637 (
            .O(N__50036),
            .I(N__49964));
    InMux I__11636 (
            .O(N__50035),
            .I(N__49961));
    InMux I__11635 (
            .O(N__50034),
            .I(N__49958));
    InMux I__11634 (
            .O(N__50033),
            .I(N__49955));
    InMux I__11633 (
            .O(N__50032),
            .I(N__49952));
    InMux I__11632 (
            .O(N__50031),
            .I(N__49949));
    InMux I__11631 (
            .O(N__50030),
            .I(N__49946));
    InMux I__11630 (
            .O(N__50029),
            .I(N__49943));
    InMux I__11629 (
            .O(N__50028),
            .I(N__49940));
    InMux I__11628 (
            .O(N__50027),
            .I(N__49936));
    LocalMux I__11627 (
            .O(N__50024),
            .I(N__49933));
    InMux I__11626 (
            .O(N__50023),
            .I(N__49930));
    LocalMux I__11625 (
            .O(N__50020),
            .I(N__49926));
    LocalMux I__11624 (
            .O(N__50017),
            .I(N__49923));
    InMux I__11623 (
            .O(N__50016),
            .I(N__49920));
    LocalMux I__11622 (
            .O(N__50013),
            .I(N__49915));
    LocalMux I__11621 (
            .O(N__50010),
            .I(N__49915));
    InMux I__11620 (
            .O(N__50009),
            .I(N__49912));
    LocalMux I__11619 (
            .O(N__50006),
            .I(N__49905));
    LocalMux I__11618 (
            .O(N__50003),
            .I(N__49905));
    LocalMux I__11617 (
            .O(N__50000),
            .I(N__49900));
    LocalMux I__11616 (
            .O(N__49997),
            .I(N__49900));
    InMux I__11615 (
            .O(N__49996),
            .I(N__49897));
    InMux I__11614 (
            .O(N__49995),
            .I(N__49894));
    CascadeMux I__11613 (
            .O(N__49994),
            .I(N__49889));
    LocalMux I__11612 (
            .O(N__49991),
            .I(N__49886));
    InMux I__11611 (
            .O(N__49990),
            .I(N__49883));
    LocalMux I__11610 (
            .O(N__49987),
            .I(N__49880));
    LocalMux I__11609 (
            .O(N__49984),
            .I(N__49877));
    LocalMux I__11608 (
            .O(N__49981),
            .I(N__49871));
    LocalMux I__11607 (
            .O(N__49978),
            .I(N__49868));
    Span4Mux_v I__11606 (
            .O(N__49973),
            .I(N__49848));
    Span4Mux_h I__11605 (
            .O(N__49970),
            .I(N__49848));
    LocalMux I__11604 (
            .O(N__49967),
            .I(N__49848));
    LocalMux I__11603 (
            .O(N__49964),
            .I(N__49848));
    LocalMux I__11602 (
            .O(N__49961),
            .I(N__49848));
    LocalMux I__11601 (
            .O(N__49958),
            .I(N__49848));
    LocalMux I__11600 (
            .O(N__49955),
            .I(N__49848));
    LocalMux I__11599 (
            .O(N__49952),
            .I(N__49848));
    LocalMux I__11598 (
            .O(N__49949),
            .I(N__49838));
    LocalMux I__11597 (
            .O(N__49946),
            .I(N__49838));
    LocalMux I__11596 (
            .O(N__49943),
            .I(N__49838));
    LocalMux I__11595 (
            .O(N__49940),
            .I(N__49838));
    InMux I__11594 (
            .O(N__49939),
            .I(N__49835));
    LocalMux I__11593 (
            .O(N__49936),
            .I(N__49828));
    Span4Mux_v I__11592 (
            .O(N__49933),
            .I(N__49823));
    LocalMux I__11591 (
            .O(N__49930),
            .I(N__49823));
    InMux I__11590 (
            .O(N__49929),
            .I(N__49820));
    Span4Mux_h I__11589 (
            .O(N__49926),
            .I(N__49813));
    Span4Mux_v I__11588 (
            .O(N__49923),
            .I(N__49813));
    LocalMux I__11587 (
            .O(N__49920),
            .I(N__49813));
    Span4Mux_v I__11586 (
            .O(N__49915),
            .I(N__49808));
    LocalMux I__11585 (
            .O(N__49912),
            .I(N__49808));
    InMux I__11584 (
            .O(N__49911),
            .I(N__49805));
    InMux I__11583 (
            .O(N__49910),
            .I(N__49802));
    Span4Mux_h I__11582 (
            .O(N__49905),
            .I(N__49793));
    Span4Mux_v I__11581 (
            .O(N__49900),
            .I(N__49793));
    LocalMux I__11580 (
            .O(N__49897),
            .I(N__49793));
    LocalMux I__11579 (
            .O(N__49894),
            .I(N__49793));
    InMux I__11578 (
            .O(N__49893),
            .I(N__49790));
    InMux I__11577 (
            .O(N__49892),
            .I(N__49784));
    InMux I__11576 (
            .O(N__49889),
            .I(N__49784));
    Span4Mux_h I__11575 (
            .O(N__49886),
            .I(N__49779));
    LocalMux I__11574 (
            .O(N__49883),
            .I(N__49779));
    Span4Mux_h I__11573 (
            .O(N__49880),
            .I(N__49774));
    Span4Mux_h I__11572 (
            .O(N__49877),
            .I(N__49774));
    InMux I__11571 (
            .O(N__49876),
            .I(N__49771));
    InMux I__11570 (
            .O(N__49875),
            .I(N__49768));
    InMux I__11569 (
            .O(N__49874),
            .I(N__49765));
    Span4Mux_h I__11568 (
            .O(N__49871),
            .I(N__49760));
    Span4Mux_h I__11567 (
            .O(N__49868),
            .I(N__49760));
    InMux I__11566 (
            .O(N__49867),
            .I(N__49757));
    InMux I__11565 (
            .O(N__49866),
            .I(N__49754));
    InMux I__11564 (
            .O(N__49865),
            .I(N__49751));
    Span4Mux_v I__11563 (
            .O(N__49848),
            .I(N__49748));
    InMux I__11562 (
            .O(N__49847),
            .I(N__49745));
    Span4Mux_v I__11561 (
            .O(N__49838),
            .I(N__49740));
    LocalMux I__11560 (
            .O(N__49835),
            .I(N__49740));
    InMux I__11559 (
            .O(N__49834),
            .I(N__49737));
    InMux I__11558 (
            .O(N__49833),
            .I(N__49734));
    InMux I__11557 (
            .O(N__49832),
            .I(N__49731));
    InMux I__11556 (
            .O(N__49831),
            .I(N__49728));
    Span4Mux_h I__11555 (
            .O(N__49828),
            .I(N__49719));
    Span4Mux_h I__11554 (
            .O(N__49823),
            .I(N__49719));
    LocalMux I__11553 (
            .O(N__49820),
            .I(N__49719));
    Span4Mux_v I__11552 (
            .O(N__49813),
            .I(N__49710));
    Span4Mux_h I__11551 (
            .O(N__49808),
            .I(N__49710));
    LocalMux I__11550 (
            .O(N__49805),
            .I(N__49710));
    LocalMux I__11549 (
            .O(N__49802),
            .I(N__49710));
    Span4Mux_h I__11548 (
            .O(N__49793),
            .I(N__49705));
    LocalMux I__11547 (
            .O(N__49790),
            .I(N__49705));
    InMux I__11546 (
            .O(N__49789),
            .I(N__49702));
    LocalMux I__11545 (
            .O(N__49784),
            .I(N__49699));
    Sp12to4 I__11544 (
            .O(N__49779),
            .I(N__49690));
    Sp12to4 I__11543 (
            .O(N__49774),
            .I(N__49690));
    LocalMux I__11542 (
            .O(N__49771),
            .I(N__49690));
    LocalMux I__11541 (
            .O(N__49768),
            .I(N__49690));
    LocalMux I__11540 (
            .O(N__49765),
            .I(N__49681));
    Sp12to4 I__11539 (
            .O(N__49760),
            .I(N__49681));
    LocalMux I__11538 (
            .O(N__49757),
            .I(N__49681));
    LocalMux I__11537 (
            .O(N__49754),
            .I(N__49681));
    LocalMux I__11536 (
            .O(N__49751),
            .I(N__49678));
    Sp12to4 I__11535 (
            .O(N__49748),
            .I(N__49673));
    LocalMux I__11534 (
            .O(N__49745),
            .I(N__49673));
    Span4Mux_v I__11533 (
            .O(N__49740),
            .I(N__49662));
    LocalMux I__11532 (
            .O(N__49737),
            .I(N__49662));
    LocalMux I__11531 (
            .O(N__49734),
            .I(N__49662));
    LocalMux I__11530 (
            .O(N__49731),
            .I(N__49662));
    LocalMux I__11529 (
            .O(N__49728),
            .I(N__49659));
    InMux I__11528 (
            .O(N__49727),
            .I(N__49656));
    InMux I__11527 (
            .O(N__49726),
            .I(N__49651));
    Span4Mux_v I__11526 (
            .O(N__49719),
            .I(N__49648));
    Span4Mux_v I__11525 (
            .O(N__49710),
            .I(N__49639));
    Span4Mux_v I__11524 (
            .O(N__49705),
            .I(N__49639));
    LocalMux I__11523 (
            .O(N__49702),
            .I(N__49639));
    Span4Mux_h I__11522 (
            .O(N__49699),
            .I(N__49639));
    Span12Mux_v I__11521 (
            .O(N__49690),
            .I(N__49636));
    Span12Mux_v I__11520 (
            .O(N__49681),
            .I(N__49629));
    Span12Mux_s10_v I__11519 (
            .O(N__49678),
            .I(N__49629));
    Span12Mux_s11_h I__11518 (
            .O(N__49673),
            .I(N__49629));
    InMux I__11517 (
            .O(N__49672),
            .I(N__49626));
    InMux I__11516 (
            .O(N__49671),
            .I(N__49623));
    Span4Mux_v I__11515 (
            .O(N__49662),
            .I(N__49616));
    Span4Mux_v I__11514 (
            .O(N__49659),
            .I(N__49616));
    LocalMux I__11513 (
            .O(N__49656),
            .I(N__49616));
    InMux I__11512 (
            .O(N__49655),
            .I(N__49613));
    InMux I__11511 (
            .O(N__49654),
            .I(N__49610));
    LocalMux I__11510 (
            .O(N__49651),
            .I(N__49603));
    Span4Mux_h I__11509 (
            .O(N__49648),
            .I(N__49603));
    Span4Mux_h I__11508 (
            .O(N__49639),
            .I(N__49603));
    Odrv12 I__11507 (
            .O(N__49636),
            .I(spi_data_mosi_7));
    Odrv12 I__11506 (
            .O(N__49629),
            .I(spi_data_mosi_7));
    LocalMux I__11505 (
            .O(N__49626),
            .I(spi_data_mosi_7));
    LocalMux I__11504 (
            .O(N__49623),
            .I(spi_data_mosi_7));
    Odrv4 I__11503 (
            .O(N__49616),
            .I(spi_data_mosi_7));
    LocalMux I__11502 (
            .O(N__49613),
            .I(spi_data_mosi_7));
    LocalMux I__11501 (
            .O(N__49610),
            .I(spi_data_mosi_7));
    Odrv4 I__11500 (
            .O(N__49603),
            .I(spi_data_mosi_7));
    InMux I__11499 (
            .O(N__49586),
            .I(N__49583));
    LocalMux I__11498 (
            .O(N__49583),
            .I(sEEADC_freqZ0Z_7));
    CEMux I__11497 (
            .O(N__49580),
            .I(N__49577));
    LocalMux I__11496 (
            .O(N__49577),
            .I(N__49573));
    CEMux I__11495 (
            .O(N__49576),
            .I(N__49570));
    Span4Mux_h I__11494 (
            .O(N__49573),
            .I(N__49565));
    LocalMux I__11493 (
            .O(N__49570),
            .I(N__49565));
    Span4Mux_h I__11492 (
            .O(N__49565),
            .I(N__49562));
    Span4Mux_h I__11491 (
            .O(N__49562),
            .I(N__49558));
    CEMux I__11490 (
            .O(N__49561),
            .I(N__49555));
    Span4Mux_h I__11489 (
            .O(N__49558),
            .I(N__49550));
    LocalMux I__11488 (
            .O(N__49555),
            .I(N__49550));
    Span4Mux_v I__11487 (
            .O(N__49550),
            .I(N__49547));
    Span4Mux_v I__11486 (
            .O(N__49547),
            .I(N__49544));
    Span4Mux_v I__11485 (
            .O(N__49544),
            .I(N__49541));
    Odrv4 I__11484 (
            .O(N__49541),
            .I(sEEADC_freq_1_sqmuxa));
    InMux I__11483 (
            .O(N__49538),
            .I(N__49519));
    InMux I__11482 (
            .O(N__49537),
            .I(N__49519));
    InMux I__11481 (
            .O(N__49536),
            .I(N__49519));
    InMux I__11480 (
            .O(N__49535),
            .I(N__49510));
    InMux I__11479 (
            .O(N__49534),
            .I(N__49510));
    InMux I__11478 (
            .O(N__49533),
            .I(N__49510));
    InMux I__11477 (
            .O(N__49532),
            .I(N__49510));
    InMux I__11476 (
            .O(N__49531),
            .I(N__49505));
    InMux I__11475 (
            .O(N__49530),
            .I(N__49505));
    InMux I__11474 (
            .O(N__49529),
            .I(N__49496));
    InMux I__11473 (
            .O(N__49528),
            .I(N__49496));
    InMux I__11472 (
            .O(N__49527),
            .I(N__49496));
    InMux I__11471 (
            .O(N__49526),
            .I(N__49496));
    LocalMux I__11470 (
            .O(N__49519),
            .I(N__49485));
    LocalMux I__11469 (
            .O(N__49510),
            .I(N__49485));
    LocalMux I__11468 (
            .O(N__49505),
            .I(N__49485));
    LocalMux I__11467 (
            .O(N__49496),
            .I(N__49485));
    CascadeMux I__11466 (
            .O(N__49495),
            .I(N__49480));
    InMux I__11465 (
            .O(N__49494),
            .I(N__49476));
    Span4Mux_v I__11464 (
            .O(N__49485),
            .I(N__49473));
    InMux I__11463 (
            .O(N__49484),
            .I(N__49470));
    InMux I__11462 (
            .O(N__49483),
            .I(N__49463));
    InMux I__11461 (
            .O(N__49480),
            .I(N__49463));
    InMux I__11460 (
            .O(N__49479),
            .I(N__49463));
    LocalMux I__11459 (
            .O(N__49476),
            .I(N__49453));
    Sp12to4 I__11458 (
            .O(N__49473),
            .I(N__49453));
    LocalMux I__11457 (
            .O(N__49470),
            .I(N__49453));
    LocalMux I__11456 (
            .O(N__49463),
            .I(N__49453));
    InMux I__11455 (
            .O(N__49462),
            .I(N__49450));
    Odrv12 I__11454 (
            .O(N__49453),
            .I(N_71));
    LocalMux I__11453 (
            .O(N__49450),
            .I(N_71));
    InMux I__11452 (
            .O(N__49445),
            .I(N__49442));
    LocalMux I__11451 (
            .O(N__49442),
            .I(N__49423));
    CEMux I__11450 (
            .O(N__49441),
            .I(N__49420));
    CascadeMux I__11449 (
            .O(N__49440),
            .I(N__49414));
    CascadeMux I__11448 (
            .O(N__49439),
            .I(N__49410));
    CascadeMux I__11447 (
            .O(N__49438),
            .I(N__49407));
    CascadeMux I__11446 (
            .O(N__49437),
            .I(N__49401));
    CascadeMux I__11445 (
            .O(N__49436),
            .I(N__49397));
    CascadeMux I__11444 (
            .O(N__49435),
            .I(N__49394));
    CascadeMux I__11443 (
            .O(N__49434),
            .I(N__49391));
    CascadeMux I__11442 (
            .O(N__49433),
            .I(N__49387));
    CascadeMux I__11441 (
            .O(N__49432),
            .I(N__49383));
    InMux I__11440 (
            .O(N__49431),
            .I(N__49372));
    InMux I__11439 (
            .O(N__49430),
            .I(N__49372));
    InMux I__11438 (
            .O(N__49429),
            .I(N__49372));
    InMux I__11437 (
            .O(N__49428),
            .I(N__49372));
    InMux I__11436 (
            .O(N__49427),
            .I(N__49369));
    CEMux I__11435 (
            .O(N__49426),
            .I(N__49366));
    Span4Mux_v I__11434 (
            .O(N__49423),
            .I(N__49359));
    LocalMux I__11433 (
            .O(N__49420),
            .I(N__49356));
    IoInMux I__11432 (
            .O(N__49419),
            .I(N__49349));
    InMux I__11431 (
            .O(N__49418),
            .I(N__49338));
    InMux I__11430 (
            .O(N__49417),
            .I(N__49338));
    InMux I__11429 (
            .O(N__49414),
            .I(N__49338));
    InMux I__11428 (
            .O(N__49413),
            .I(N__49338));
    InMux I__11427 (
            .O(N__49410),
            .I(N__49338));
    InMux I__11426 (
            .O(N__49407),
            .I(N__49321));
    InMux I__11425 (
            .O(N__49406),
            .I(N__49321));
    InMux I__11424 (
            .O(N__49405),
            .I(N__49321));
    InMux I__11423 (
            .O(N__49404),
            .I(N__49321));
    InMux I__11422 (
            .O(N__49401),
            .I(N__49321));
    InMux I__11421 (
            .O(N__49400),
            .I(N__49321));
    InMux I__11420 (
            .O(N__49397),
            .I(N__49321));
    InMux I__11419 (
            .O(N__49394),
            .I(N__49321));
    InMux I__11418 (
            .O(N__49391),
            .I(N__49318));
    CascadeMux I__11417 (
            .O(N__49390),
            .I(N__49315));
    InMux I__11416 (
            .O(N__49387),
            .I(N__49308));
    InMux I__11415 (
            .O(N__49386),
            .I(N__49308));
    InMux I__11414 (
            .O(N__49383),
            .I(N__49308));
    InMux I__11413 (
            .O(N__49382),
            .I(N__49299));
    InMux I__11412 (
            .O(N__49381),
            .I(N__49296));
    LocalMux I__11411 (
            .O(N__49372),
            .I(N__49283));
    LocalMux I__11410 (
            .O(N__49369),
            .I(N__49283));
    LocalMux I__11409 (
            .O(N__49366),
            .I(N__49280));
    InMux I__11408 (
            .O(N__49365),
            .I(N__49275));
    InMux I__11407 (
            .O(N__49364),
            .I(N__49275));
    CascadeMux I__11406 (
            .O(N__49363),
            .I(N__49272));
    CascadeMux I__11405 (
            .O(N__49362),
            .I(N__49269));
    Span4Mux_h I__11404 (
            .O(N__49359),
            .I(N__49264));
    Span4Mux_v I__11403 (
            .O(N__49356),
            .I(N__49264));
    CascadeMux I__11402 (
            .O(N__49355),
            .I(N__49261));
    InMux I__11401 (
            .O(N__49354),
            .I(N__49257));
    CascadeMux I__11400 (
            .O(N__49353),
            .I(N__49254));
    CascadeMux I__11399 (
            .O(N__49352),
            .I(N__49250));
    LocalMux I__11398 (
            .O(N__49349),
            .I(N__49247));
    LocalMux I__11397 (
            .O(N__49338),
            .I(N__49241));
    LocalMux I__11396 (
            .O(N__49321),
            .I(N__49241));
    LocalMux I__11395 (
            .O(N__49318),
            .I(N__49237));
    InMux I__11394 (
            .O(N__49315),
            .I(N__49234));
    LocalMux I__11393 (
            .O(N__49308),
            .I(N__49231));
    InMux I__11392 (
            .O(N__49307),
            .I(N__49224));
    InMux I__11391 (
            .O(N__49306),
            .I(N__49224));
    InMux I__11390 (
            .O(N__49305),
            .I(N__49224));
    InMux I__11389 (
            .O(N__49304),
            .I(N__49217));
    InMux I__11388 (
            .O(N__49303),
            .I(N__49217));
    InMux I__11387 (
            .O(N__49302),
            .I(N__49217));
    LocalMux I__11386 (
            .O(N__49299),
            .I(N__49212));
    LocalMux I__11385 (
            .O(N__49296),
            .I(N__49212));
    InMux I__11384 (
            .O(N__49295),
            .I(N__49203));
    InMux I__11383 (
            .O(N__49294),
            .I(N__49203));
    InMux I__11382 (
            .O(N__49293),
            .I(N__49203));
    InMux I__11381 (
            .O(N__49292),
            .I(N__49203));
    InMux I__11380 (
            .O(N__49291),
            .I(N__49194));
    InMux I__11379 (
            .O(N__49290),
            .I(N__49194));
    InMux I__11378 (
            .O(N__49289),
            .I(N__49194));
    InMux I__11377 (
            .O(N__49288),
            .I(N__49194));
    Span4Mux_v I__11376 (
            .O(N__49283),
            .I(N__49188));
    Span4Mux_h I__11375 (
            .O(N__49280),
            .I(N__49185));
    LocalMux I__11374 (
            .O(N__49275),
            .I(N__49182));
    InMux I__11373 (
            .O(N__49272),
            .I(N__49179));
    InMux I__11372 (
            .O(N__49269),
            .I(N__49176));
    Span4Mux_v I__11371 (
            .O(N__49264),
            .I(N__49173));
    InMux I__11370 (
            .O(N__49261),
            .I(N__49170));
    CascadeMux I__11369 (
            .O(N__49260),
            .I(N__49167));
    LocalMux I__11368 (
            .O(N__49257),
            .I(N__49164));
    InMux I__11367 (
            .O(N__49254),
            .I(N__49161));
    InMux I__11366 (
            .O(N__49253),
            .I(N__49158));
    InMux I__11365 (
            .O(N__49250),
            .I(N__49155));
    Span4Mux_s2_h I__11364 (
            .O(N__49247),
            .I(N__49152));
    InMux I__11363 (
            .O(N__49246),
            .I(N__49149));
    Span4Mux_v I__11362 (
            .O(N__49241),
            .I(N__49146));
    InMux I__11361 (
            .O(N__49240),
            .I(N__49142));
    Span4Mux_v I__11360 (
            .O(N__49237),
            .I(N__49137));
    LocalMux I__11359 (
            .O(N__49234),
            .I(N__49137));
    Span4Mux_h I__11358 (
            .O(N__49231),
            .I(N__49124));
    LocalMux I__11357 (
            .O(N__49224),
            .I(N__49124));
    LocalMux I__11356 (
            .O(N__49217),
            .I(N__49124));
    Span4Mux_h I__11355 (
            .O(N__49212),
            .I(N__49124));
    LocalMux I__11354 (
            .O(N__49203),
            .I(N__49124));
    LocalMux I__11353 (
            .O(N__49194),
            .I(N__49124));
    InMux I__11352 (
            .O(N__49193),
            .I(N__49117));
    InMux I__11351 (
            .O(N__49192),
            .I(N__49117));
    InMux I__11350 (
            .O(N__49191),
            .I(N__49117));
    Span4Mux_h I__11349 (
            .O(N__49188),
            .I(N__49105));
    Span4Mux_h I__11348 (
            .O(N__49185),
            .I(N__49105));
    Span4Mux_h I__11347 (
            .O(N__49182),
            .I(N__49105));
    LocalMux I__11346 (
            .O(N__49179),
            .I(N__49105));
    LocalMux I__11345 (
            .O(N__49176),
            .I(N__49105));
    Span4Mux_h I__11344 (
            .O(N__49173),
            .I(N__49102));
    LocalMux I__11343 (
            .O(N__49170),
            .I(N__49099));
    InMux I__11342 (
            .O(N__49167),
            .I(N__49096));
    Span4Mux_v I__11341 (
            .O(N__49164),
            .I(N__49088));
    LocalMux I__11340 (
            .O(N__49161),
            .I(N__49088));
    LocalMux I__11339 (
            .O(N__49158),
            .I(N__49088));
    LocalMux I__11338 (
            .O(N__49155),
            .I(N__49085));
    Sp12to4 I__11337 (
            .O(N__49152),
            .I(N__49082));
    LocalMux I__11336 (
            .O(N__49149),
            .I(N__49079));
    Span4Mux_v I__11335 (
            .O(N__49146),
            .I(N__49076));
    InMux I__11334 (
            .O(N__49145),
            .I(N__49073));
    LocalMux I__11333 (
            .O(N__49142),
            .I(N__49064));
    Span4Mux_v I__11332 (
            .O(N__49137),
            .I(N__49064));
    Span4Mux_v I__11331 (
            .O(N__49124),
            .I(N__49064));
    LocalMux I__11330 (
            .O(N__49117),
            .I(N__49064));
    InMux I__11329 (
            .O(N__49116),
            .I(N__49061));
    Span4Mux_v I__11328 (
            .O(N__49105),
            .I(N__49058));
    Span4Mux_v I__11327 (
            .O(N__49102),
            .I(N__49053));
    Span4Mux_v I__11326 (
            .O(N__49099),
            .I(N__49053));
    LocalMux I__11325 (
            .O(N__49096),
            .I(N__49050));
    InMux I__11324 (
            .O(N__49095),
            .I(N__49046));
    Span4Mux_h I__11323 (
            .O(N__49088),
            .I(N__49043));
    Span4Mux_v I__11322 (
            .O(N__49085),
            .I(N__49040));
    Span12Mux_v I__11321 (
            .O(N__49082),
            .I(N__49037));
    Sp12to4 I__11320 (
            .O(N__49079),
            .I(N__49034));
    Sp12to4 I__11319 (
            .O(N__49076),
            .I(N__49027));
    LocalMux I__11318 (
            .O(N__49073),
            .I(N__49027));
    Sp12to4 I__11317 (
            .O(N__49064),
            .I(N__49027));
    LocalMux I__11316 (
            .O(N__49061),
            .I(N__49024));
    Span4Mux_v I__11315 (
            .O(N__49058),
            .I(N__49021));
    Span4Mux_v I__11314 (
            .O(N__49053),
            .I(N__49018));
    Span4Mux_v I__11313 (
            .O(N__49050),
            .I(N__49015));
    IoInMux I__11312 (
            .O(N__49049),
            .I(N__49012));
    LocalMux I__11311 (
            .O(N__49046),
            .I(N__49007));
    Sp12to4 I__11310 (
            .O(N__49043),
            .I(N__49007));
    Span4Mux_h I__11309 (
            .O(N__49040),
            .I(N__49004));
    Span12Mux_v I__11308 (
            .O(N__49037),
            .I(N__49001));
    Span12Mux_v I__11307 (
            .O(N__49034),
            .I(N__48994));
    Span12Mux_h I__11306 (
            .O(N__49027),
            .I(N__48994));
    Span12Mux_h I__11305 (
            .O(N__49024),
            .I(N__48994));
    Sp12to4 I__11304 (
            .O(N__49021),
            .I(N__48987));
    Sp12to4 I__11303 (
            .O(N__49018),
            .I(N__48987));
    Sp12to4 I__11302 (
            .O(N__49015),
            .I(N__48987));
    LocalMux I__11301 (
            .O(N__49012),
            .I(N__48984));
    Span12Mux_v I__11300 (
            .O(N__49007),
            .I(N__48979));
    Sp12to4 I__11299 (
            .O(N__49004),
            .I(N__48979));
    Span12Mux_h I__11298 (
            .O(N__49001),
            .I(N__48972));
    Span12Mux_v I__11297 (
            .O(N__48994),
            .I(N__48972));
    Span12Mux_h I__11296 (
            .O(N__48987),
            .I(N__48972));
    IoSpan4Mux I__11295 (
            .O(N__48984),
            .I(N__48969));
    Odrv12 I__11294 (
            .O(N__48979),
            .I(LED3_c));
    Odrv12 I__11293 (
            .O(N__48972),
            .I(LED3_c));
    Odrv4 I__11292 (
            .O(N__48969),
            .I(LED3_c));
    InMux I__11291 (
            .O(N__48962),
            .I(N__48957));
    InMux I__11290 (
            .O(N__48961),
            .I(N__48953));
    CEMux I__11289 (
            .O(N__48960),
            .I(N__48943));
    LocalMux I__11288 (
            .O(N__48957),
            .I(N__48940));
    InMux I__11287 (
            .O(N__48956),
            .I(N__48937));
    LocalMux I__11286 (
            .O(N__48953),
            .I(N__48926));
    InMux I__11285 (
            .O(N__48952),
            .I(N__48923));
    InMux I__11284 (
            .O(N__48951),
            .I(N__48912));
    InMux I__11283 (
            .O(N__48950),
            .I(N__48912));
    InMux I__11282 (
            .O(N__48949),
            .I(N__48912));
    InMux I__11281 (
            .O(N__48948),
            .I(N__48912));
    InMux I__11280 (
            .O(N__48947),
            .I(N__48912));
    InMux I__11279 (
            .O(N__48946),
            .I(N__48904));
    LocalMux I__11278 (
            .O(N__48943),
            .I(N__48894));
    Span4Mux_h I__11277 (
            .O(N__48940),
            .I(N__48889));
    LocalMux I__11276 (
            .O(N__48937),
            .I(N__48889));
    InMux I__11275 (
            .O(N__48936),
            .I(N__48872));
    InMux I__11274 (
            .O(N__48935),
            .I(N__48872));
    InMux I__11273 (
            .O(N__48934),
            .I(N__48872));
    InMux I__11272 (
            .O(N__48933),
            .I(N__48872));
    InMux I__11271 (
            .O(N__48932),
            .I(N__48872));
    InMux I__11270 (
            .O(N__48931),
            .I(N__48872));
    InMux I__11269 (
            .O(N__48930),
            .I(N__48872));
    InMux I__11268 (
            .O(N__48929),
            .I(N__48872));
    Span4Mux_v I__11267 (
            .O(N__48926),
            .I(N__48867));
    LocalMux I__11266 (
            .O(N__48923),
            .I(N__48867));
    LocalMux I__11265 (
            .O(N__48912),
            .I(N__48864));
    InMux I__11264 (
            .O(N__48911),
            .I(N__48853));
    InMux I__11263 (
            .O(N__48910),
            .I(N__48853));
    InMux I__11262 (
            .O(N__48909),
            .I(N__48853));
    InMux I__11261 (
            .O(N__48908),
            .I(N__48853));
    InMux I__11260 (
            .O(N__48907),
            .I(N__48853));
    LocalMux I__11259 (
            .O(N__48904),
            .I(N__48850));
    InMux I__11258 (
            .O(N__48903),
            .I(N__48845));
    InMux I__11257 (
            .O(N__48902),
            .I(N__48845));
    InMux I__11256 (
            .O(N__48901),
            .I(N__48834));
    InMux I__11255 (
            .O(N__48900),
            .I(N__48834));
    InMux I__11254 (
            .O(N__48899),
            .I(N__48834));
    InMux I__11253 (
            .O(N__48898),
            .I(N__48834));
    InMux I__11252 (
            .O(N__48897),
            .I(N__48834));
    Odrv4 I__11251 (
            .O(N__48894),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    Odrv4 I__11250 (
            .O(N__48889),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    LocalMux I__11249 (
            .O(N__48872),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    Odrv4 I__11248 (
            .O(N__48867),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    Odrv4 I__11247 (
            .O(N__48864),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    LocalMux I__11246 (
            .O(N__48853),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    Odrv4 I__11245 (
            .O(N__48850),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    LocalMux I__11244 (
            .O(N__48845),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    LocalMux I__11243 (
            .O(N__48834),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    IoInMux I__11242 (
            .O(N__48815),
            .I(N__48812));
    LocalMux I__11241 (
            .O(N__48812),
            .I(N__48809));
    Span4Mux_s3_h I__11240 (
            .O(N__48809),
            .I(N__48806));
    Span4Mux_v I__11239 (
            .O(N__48806),
            .I(N__48803));
    Span4Mux_h I__11238 (
            .O(N__48803),
            .I(N__48799));
    InMux I__11237 (
            .O(N__48802),
            .I(N__48796));
    Odrv4 I__11236 (
            .O(N__48799),
            .I(RAM_DATA_cl_5Z0Z_15));
    LocalMux I__11235 (
            .O(N__48796),
            .I(RAM_DATA_cl_5Z0Z_15));
    CascadeMux I__11234 (
            .O(N__48791),
            .I(N__48787));
    InMux I__11233 (
            .O(N__48790),
            .I(N__48784));
    InMux I__11232 (
            .O(N__48787),
            .I(N__48781));
    LocalMux I__11231 (
            .O(N__48784),
            .I(N__48776));
    LocalMux I__11230 (
            .O(N__48781),
            .I(N__48776));
    Odrv4 I__11229 (
            .O(N__48776),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1 ));
    InMux I__11228 (
            .O(N__48773),
            .I(N__48766));
    InMux I__11227 (
            .O(N__48772),
            .I(N__48766));
    InMux I__11226 (
            .O(N__48771),
            .I(N__48763));
    LocalMux I__11225 (
            .O(N__48766),
            .I(N__48760));
    LocalMux I__11224 (
            .O(N__48763),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0 ));
    Odrv4 I__11223 (
            .O(N__48760),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0 ));
    InMux I__11222 (
            .O(N__48755),
            .I(N__48745));
    InMux I__11221 (
            .O(N__48754),
            .I(N__48745));
    InMux I__11220 (
            .O(N__48753),
            .I(N__48745));
    InMux I__11219 (
            .O(N__48752),
            .I(N__48742));
    LocalMux I__11218 (
            .O(N__48745),
            .I(N__48739));
    LocalMux I__11217 (
            .O(N__48742),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1 ));
    Odrv4 I__11216 (
            .O(N__48739),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1 ));
    InMux I__11215 (
            .O(N__48734),
            .I(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0 ));
    InMux I__11214 (
            .O(N__48731),
            .I(N__48722));
    InMux I__11213 (
            .O(N__48730),
            .I(N__48722));
    InMux I__11212 (
            .O(N__48729),
            .I(N__48722));
    LocalMux I__11211 (
            .O(N__48722),
            .I(N__48719));
    Span4Mux_v I__11210 (
            .O(N__48719),
            .I(N__48714));
    InMux I__11209 (
            .O(N__48718),
            .I(N__48708));
    InMux I__11208 (
            .O(N__48717),
            .I(N__48708));
    Span4Mux_h I__11207 (
            .O(N__48714),
            .I(N__48705));
    InMux I__11206 (
            .O(N__48713),
            .I(N__48702));
    LocalMux I__11205 (
            .O(N__48708),
            .I(N__48699));
    Odrv4 I__11204 (
            .O(N__48705),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2 ));
    LocalMux I__11203 (
            .O(N__48702),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2 ));
    Odrv4 I__11202 (
            .O(N__48699),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2 ));
    InMux I__11201 (
            .O(N__48692),
            .I(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1 ));
    CascadeMux I__11200 (
            .O(N__48689),
            .I(N__48686));
    InMux I__11199 (
            .O(N__48686),
            .I(N__48682));
    InMux I__11198 (
            .O(N__48685),
            .I(N__48679));
    LocalMux I__11197 (
            .O(N__48682),
            .I(N__48676));
    LocalMux I__11196 (
            .O(N__48679),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3 ));
    Odrv4 I__11195 (
            .O(N__48676),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3 ));
    InMux I__11194 (
            .O(N__48671),
            .I(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2 ));
    InMux I__11193 (
            .O(N__48668),
            .I(N__48662));
    InMux I__11192 (
            .O(N__48667),
            .I(N__48659));
    InMux I__11191 (
            .O(N__48666),
            .I(N__48656));
    InMux I__11190 (
            .O(N__48665),
            .I(N__48653));
    LocalMux I__11189 (
            .O(N__48662),
            .I(N__48650));
    LocalMux I__11188 (
            .O(N__48659),
            .I(sCounterDACZ0Z_3));
    LocalMux I__11187 (
            .O(N__48656),
            .I(sCounterDACZ0Z_3));
    LocalMux I__11186 (
            .O(N__48653),
            .I(sCounterDACZ0Z_3));
    Odrv4 I__11185 (
            .O(N__48650),
            .I(sCounterDACZ0Z_3));
    InMux I__11184 (
            .O(N__48641),
            .I(un2_scounterdac_cry_2));
    InMux I__11183 (
            .O(N__48638),
            .I(N__48633));
    InMux I__11182 (
            .O(N__48637),
            .I(N__48628));
    InMux I__11181 (
            .O(N__48636),
            .I(N__48628));
    LocalMux I__11180 (
            .O(N__48633),
            .I(sCounterDACZ0Z_4));
    LocalMux I__11179 (
            .O(N__48628),
            .I(sCounterDACZ0Z_4));
    InMux I__11178 (
            .O(N__48623),
            .I(un2_scounterdac_cry_3));
    CascadeMux I__11177 (
            .O(N__48620),
            .I(N__48615));
    CascadeMux I__11176 (
            .O(N__48619),
            .I(N__48612));
    InMux I__11175 (
            .O(N__48618),
            .I(N__48608));
    InMux I__11174 (
            .O(N__48615),
            .I(N__48601));
    InMux I__11173 (
            .O(N__48612),
            .I(N__48601));
    InMux I__11172 (
            .O(N__48611),
            .I(N__48601));
    LocalMux I__11171 (
            .O(N__48608),
            .I(sCounterDACZ0Z_5));
    LocalMux I__11170 (
            .O(N__48601),
            .I(sCounterDACZ0Z_5));
    InMux I__11169 (
            .O(N__48596),
            .I(un2_scounterdac_cry_4));
    InMux I__11168 (
            .O(N__48593),
            .I(N__48588));
    InMux I__11167 (
            .O(N__48592),
            .I(N__48583));
    InMux I__11166 (
            .O(N__48591),
            .I(N__48583));
    LocalMux I__11165 (
            .O(N__48588),
            .I(sCounterDACZ0Z_6));
    LocalMux I__11164 (
            .O(N__48583),
            .I(sCounterDACZ0Z_6));
    InMux I__11163 (
            .O(N__48578),
            .I(N__48575));
    LocalMux I__11162 (
            .O(N__48575),
            .I(un2_scounterdac_cry_5_THRU_CO));
    InMux I__11161 (
            .O(N__48572),
            .I(un2_scounterdac_cry_5));
    InMux I__11160 (
            .O(N__48569),
            .I(N__48565));
    InMux I__11159 (
            .O(N__48568),
            .I(N__48562));
    LocalMux I__11158 (
            .O(N__48565),
            .I(sCounterDACZ0Z_7));
    LocalMux I__11157 (
            .O(N__48562),
            .I(sCounterDACZ0Z_7));
    InMux I__11156 (
            .O(N__48557),
            .I(un2_scounterdac_cry_6));
    InMux I__11155 (
            .O(N__48554),
            .I(N__48550));
    InMux I__11154 (
            .O(N__48553),
            .I(N__48547));
    LocalMux I__11153 (
            .O(N__48550),
            .I(N__48544));
    LocalMux I__11152 (
            .O(N__48547),
            .I(N_30_mux));
    Odrv4 I__11151 (
            .O(N__48544),
            .I(N_30_mux));
    InMux I__11150 (
            .O(N__48539),
            .I(N__48536));
    LocalMux I__11149 (
            .O(N__48536),
            .I(N__48530));
    InMux I__11148 (
            .O(N__48535),
            .I(N__48527));
    InMux I__11147 (
            .O(N__48534),
            .I(N__48522));
    InMux I__11146 (
            .O(N__48533),
            .I(N__48522));
    Odrv12 I__11145 (
            .O(N__48530),
            .I(sCounterDACZ0Z_8));
    LocalMux I__11144 (
            .O(N__48527),
            .I(sCounterDACZ0Z_8));
    LocalMux I__11143 (
            .O(N__48522),
            .I(sCounterDACZ0Z_8));
    InMux I__11142 (
            .O(N__48515),
            .I(un2_scounterdac_cry_7));
    InMux I__11141 (
            .O(N__48512),
            .I(bfn_20_11_0_));
    CascadeMux I__11140 (
            .O(N__48509),
            .I(N__48506));
    InMux I__11139 (
            .O(N__48506),
            .I(N__48502));
    InMux I__11138 (
            .O(N__48505),
            .I(N__48499));
    LocalMux I__11137 (
            .O(N__48502),
            .I(N__48496));
    LocalMux I__11136 (
            .O(N__48499),
            .I(sCounterDACZ0Z_9));
    Odrv4 I__11135 (
            .O(N__48496),
            .I(sCounterDACZ0Z_9));
    ClkMux I__11134 (
            .O(N__48491),
            .I(N__48347));
    ClkMux I__11133 (
            .O(N__48490),
            .I(N__48347));
    ClkMux I__11132 (
            .O(N__48489),
            .I(N__48347));
    ClkMux I__11131 (
            .O(N__48488),
            .I(N__48347));
    ClkMux I__11130 (
            .O(N__48487),
            .I(N__48347));
    ClkMux I__11129 (
            .O(N__48486),
            .I(N__48347));
    ClkMux I__11128 (
            .O(N__48485),
            .I(N__48347));
    ClkMux I__11127 (
            .O(N__48484),
            .I(N__48347));
    ClkMux I__11126 (
            .O(N__48483),
            .I(N__48347));
    ClkMux I__11125 (
            .O(N__48482),
            .I(N__48347));
    ClkMux I__11124 (
            .O(N__48481),
            .I(N__48347));
    ClkMux I__11123 (
            .O(N__48480),
            .I(N__48347));
    ClkMux I__11122 (
            .O(N__48479),
            .I(N__48347));
    ClkMux I__11121 (
            .O(N__48478),
            .I(N__48347));
    ClkMux I__11120 (
            .O(N__48477),
            .I(N__48347));
    ClkMux I__11119 (
            .O(N__48476),
            .I(N__48347));
    ClkMux I__11118 (
            .O(N__48475),
            .I(N__48347));
    ClkMux I__11117 (
            .O(N__48474),
            .I(N__48347));
    ClkMux I__11116 (
            .O(N__48473),
            .I(N__48347));
    ClkMux I__11115 (
            .O(N__48472),
            .I(N__48347));
    ClkMux I__11114 (
            .O(N__48471),
            .I(N__48347));
    ClkMux I__11113 (
            .O(N__48470),
            .I(N__48347));
    ClkMux I__11112 (
            .O(N__48469),
            .I(N__48347));
    ClkMux I__11111 (
            .O(N__48468),
            .I(N__48347));
    ClkMux I__11110 (
            .O(N__48467),
            .I(N__48347));
    ClkMux I__11109 (
            .O(N__48466),
            .I(N__48347));
    ClkMux I__11108 (
            .O(N__48465),
            .I(N__48347));
    ClkMux I__11107 (
            .O(N__48464),
            .I(N__48347));
    ClkMux I__11106 (
            .O(N__48463),
            .I(N__48347));
    ClkMux I__11105 (
            .O(N__48462),
            .I(N__48347));
    ClkMux I__11104 (
            .O(N__48461),
            .I(N__48347));
    ClkMux I__11103 (
            .O(N__48460),
            .I(N__48347));
    ClkMux I__11102 (
            .O(N__48459),
            .I(N__48347));
    ClkMux I__11101 (
            .O(N__48458),
            .I(N__48347));
    ClkMux I__11100 (
            .O(N__48457),
            .I(N__48347));
    ClkMux I__11099 (
            .O(N__48456),
            .I(N__48347));
    ClkMux I__11098 (
            .O(N__48455),
            .I(N__48347));
    ClkMux I__11097 (
            .O(N__48454),
            .I(N__48347));
    ClkMux I__11096 (
            .O(N__48453),
            .I(N__48347));
    ClkMux I__11095 (
            .O(N__48452),
            .I(N__48347));
    ClkMux I__11094 (
            .O(N__48451),
            .I(N__48347));
    ClkMux I__11093 (
            .O(N__48450),
            .I(N__48347));
    ClkMux I__11092 (
            .O(N__48449),
            .I(N__48347));
    ClkMux I__11091 (
            .O(N__48448),
            .I(N__48347));
    ClkMux I__11090 (
            .O(N__48447),
            .I(N__48347));
    ClkMux I__11089 (
            .O(N__48446),
            .I(N__48347));
    ClkMux I__11088 (
            .O(N__48445),
            .I(N__48347));
    ClkMux I__11087 (
            .O(N__48444),
            .I(N__48347));
    GlobalMux I__11086 (
            .O(N__48347),
            .I(N__48344));
    gio2CtrlBuf I__11085 (
            .O(N__48344),
            .I(pll_clk64_0_g));
    InMux I__11084 (
            .O(N__48341),
            .I(N__48338));
    LocalMux I__11083 (
            .O(N__48338),
            .I(N__48335));
    Span12Mux_h I__11082 (
            .O(N__48335),
            .I(N__48332));
    Odrv12 I__11081 (
            .O(N__48332),
            .I(\spi_slave_inst.un23_i_ssn_3 ));
    InMux I__11080 (
            .O(N__48329),
            .I(N__48325));
    InMux I__11079 (
            .O(N__48328),
            .I(N__48321));
    LocalMux I__11078 (
            .O(N__48325),
            .I(N__48318));
    InMux I__11077 (
            .O(N__48324),
            .I(N__48315));
    LocalMux I__11076 (
            .O(N__48321),
            .I(N__48310));
    Span12Mux_h I__11075 (
            .O(N__48318),
            .I(N__48310));
    LocalMux I__11074 (
            .O(N__48315),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4 ));
    Odrv12 I__11073 (
            .O(N__48310),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4 ));
    InMux I__11072 (
            .O(N__48305),
            .I(N__48300));
    InMux I__11071 (
            .O(N__48304),
            .I(N__48297));
    InMux I__11070 (
            .O(N__48303),
            .I(N__48294));
    LocalMux I__11069 (
            .O(N__48300),
            .I(N__48289));
    LocalMux I__11068 (
            .O(N__48297),
            .I(N__48289));
    LocalMux I__11067 (
            .O(N__48294),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3 ));
    Odrv12 I__11066 (
            .O(N__48289),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3 ));
    InMux I__11065 (
            .O(N__48284),
            .I(N__48281));
    LocalMux I__11064 (
            .O(N__48281),
            .I(N__48278));
    Span12Mux_v I__11063 (
            .O(N__48278),
            .I(N__48275));
    Span12Mux_h I__11062 (
            .O(N__48275),
            .I(N__48272));
    Span12Mux_v I__11061 (
            .O(N__48272),
            .I(N__48269));
    Odrv12 I__11060 (
            .O(N__48269),
            .I(\spi_slave_inst.rx_done_pos_sclk_iZ0 ));
    ClkMux I__11059 (
            .O(N__48266),
            .I(N__48242));
    ClkMux I__11058 (
            .O(N__48265),
            .I(N__48242));
    ClkMux I__11057 (
            .O(N__48264),
            .I(N__48242));
    ClkMux I__11056 (
            .O(N__48263),
            .I(N__48242));
    ClkMux I__11055 (
            .O(N__48262),
            .I(N__48242));
    ClkMux I__11054 (
            .O(N__48261),
            .I(N__48242));
    ClkMux I__11053 (
            .O(N__48260),
            .I(N__48242));
    ClkMux I__11052 (
            .O(N__48259),
            .I(N__48242));
    GlobalMux I__11051 (
            .O(N__48242),
            .I(N__48239));
    gio2CtrlBuf I__11050 (
            .O(N__48239),
            .I(spi_sclk_g));
    CEMux I__11049 (
            .O(N__48236),
            .I(N__48233));
    LocalMux I__11048 (
            .O(N__48233),
            .I(N__48228));
    CEMux I__11047 (
            .O(N__48232),
            .I(N__48225));
    CEMux I__11046 (
            .O(N__48231),
            .I(N__48222));
    Span4Mux_h I__11045 (
            .O(N__48228),
            .I(N__48219));
    LocalMux I__11044 (
            .O(N__48225),
            .I(N__48216));
    LocalMux I__11043 (
            .O(N__48222),
            .I(N__48213));
    Span4Mux_v I__11042 (
            .O(N__48219),
            .I(N__48210));
    Span4Mux_v I__11041 (
            .O(N__48216),
            .I(N__48207));
    Span12Mux_h I__11040 (
            .O(N__48213),
            .I(N__48204));
    Span4Mux_v I__11039 (
            .O(N__48210),
            .I(N__48201));
    Span4Mux_h I__11038 (
            .O(N__48207),
            .I(N__48198));
    Odrv12 I__11037 (
            .O(N__48204),
            .I(\spi_slave_inst.spi_cs_iZ0 ));
    Odrv4 I__11036 (
            .O(N__48201),
            .I(\spi_slave_inst.spi_cs_iZ0 ));
    Odrv4 I__11035 (
            .O(N__48198),
            .I(\spi_slave_inst.spi_cs_iZ0 ));
    CascadeMux I__11034 (
            .O(N__48191),
            .I(N_23_mux_cascade_));
    CascadeMux I__11033 (
            .O(N__48188),
            .I(N_25_mux_cascade_));
    InMux I__11032 (
            .O(N__48185),
            .I(N__48182));
    LocalMux I__11031 (
            .O(N__48182),
            .I(m15_1));
    IoInMux I__11030 (
            .O(N__48179),
            .I(N__48176));
    LocalMux I__11029 (
            .O(N__48176),
            .I(N__48173));
    IoSpan4Mux I__11028 (
            .O(N__48173),
            .I(N__48170));
    Span4Mux_s0_h I__11027 (
            .O(N__48170),
            .I(N__48167));
    Span4Mux_h I__11026 (
            .O(N__48167),
            .I(N__48164));
    Odrv4 I__11025 (
            .O(N__48164),
            .I(op_eq_scounterdac10));
    InMux I__11024 (
            .O(N__48161),
            .I(N__48158));
    LocalMux I__11023 (
            .O(N__48158),
            .I(m8_2));
    InMux I__11022 (
            .O(N__48155),
            .I(N__48152));
    LocalMux I__11021 (
            .O(N__48152),
            .I(N_23_mux));
    CascadeMux I__11020 (
            .O(N__48149),
            .I(N_30_mux_cascade_));
    InMux I__11019 (
            .O(N__48146),
            .I(N__48143));
    LocalMux I__11018 (
            .O(N__48143),
            .I(N_25_mux));
    InMux I__11017 (
            .O(N__48140),
            .I(N__48137));
    LocalMux I__11016 (
            .O(N__48137),
            .I(N__48134));
    Odrv12 I__11015 (
            .O(N__48134),
            .I(N_32_mux));
    InMux I__11014 (
            .O(N__48131),
            .I(N__48119));
    InMux I__11013 (
            .O(N__48130),
            .I(N__48119));
    InMux I__11012 (
            .O(N__48129),
            .I(N__48119));
    InMux I__11011 (
            .O(N__48128),
            .I(N__48116));
    InMux I__11010 (
            .O(N__48127),
            .I(N__48113));
    InMux I__11009 (
            .O(N__48126),
            .I(N__48110));
    LocalMux I__11008 (
            .O(N__48119),
            .I(N__48103));
    LocalMux I__11007 (
            .O(N__48116),
            .I(N__48103));
    LocalMux I__11006 (
            .O(N__48113),
            .I(N__48103));
    LocalMux I__11005 (
            .O(N__48110),
            .I(sCounterDACZ0Z_0));
    Odrv12 I__11004 (
            .O(N__48103),
            .I(sCounterDACZ0Z_0));
    CascadeMux I__11003 (
            .O(N__48098),
            .I(N__48094));
    CascadeMux I__11002 (
            .O(N__48097),
            .I(N__48091));
    InMux I__11001 (
            .O(N__48094),
            .I(N__48086));
    InMux I__11000 (
            .O(N__48091),
            .I(N__48079));
    InMux I__10999 (
            .O(N__48090),
            .I(N__48079));
    InMux I__10998 (
            .O(N__48089),
            .I(N__48079));
    LocalMux I__10997 (
            .O(N__48086),
            .I(sCounterDACZ0Z_1));
    LocalMux I__10996 (
            .O(N__48079),
            .I(sCounterDACZ0Z_1));
    InMux I__10995 (
            .O(N__48074),
            .I(N__48070));
    InMux I__10994 (
            .O(N__48073),
            .I(N__48067));
    LocalMux I__10993 (
            .O(N__48070),
            .I(sCounterDACZ0Z_2));
    LocalMux I__10992 (
            .O(N__48067),
            .I(sCounterDACZ0Z_2));
    InMux I__10991 (
            .O(N__48062),
            .I(un2_scounterdac_cry_1));
    CascadeMux I__10990 (
            .O(N__48059),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_ ));
    InMux I__10989 (
            .O(N__48056),
            .I(N__48053));
    LocalMux I__10988 (
            .O(N__48053),
            .I(N__48048));
    InMux I__10987 (
            .O(N__48052),
            .I(N__48045));
    InMux I__10986 (
            .O(N__48051),
            .I(N__48042));
    Span4Mux_v I__10985 (
            .O(N__48048),
            .I(N__48038));
    LocalMux I__10984 (
            .O(N__48045),
            .I(N__48033));
    LocalMux I__10983 (
            .O(N__48042),
            .I(N__48033));
    InMux I__10982 (
            .O(N__48041),
            .I(N__48029));
    Span4Mux_v I__10981 (
            .O(N__48038),
            .I(N__48024));
    Span4Mux_v I__10980 (
            .O(N__48033),
            .I(N__48024));
    InMux I__10979 (
            .O(N__48032),
            .I(N__48021));
    LocalMux I__10978 (
            .O(N__48029),
            .I(N__48018));
    Span4Mux_h I__10977 (
            .O(N__48024),
            .I(N__48015));
    LocalMux I__10976 (
            .O(N__48021),
            .I(N__48012));
    Span4Mux_h I__10975 (
            .O(N__48018),
            .I(N__48008));
    Span4Mux_h I__10974 (
            .O(N__48015),
            .I(N__48001));
    Span4Mux_v I__10973 (
            .O(N__48012),
            .I(N__48001));
    InMux I__10972 (
            .O(N__48011),
            .I(N__47998));
    Span4Mux_h I__10971 (
            .O(N__48008),
            .I(N__47995));
    InMux I__10970 (
            .O(N__48007),
            .I(N__47992));
    InMux I__10969 (
            .O(N__48006),
            .I(N__47989));
    Span4Mux_h I__10968 (
            .O(N__48001),
            .I(N__47984));
    LocalMux I__10967 (
            .O(N__47998),
            .I(N__47984));
    Sp12to4 I__10966 (
            .O(N__47995),
            .I(N__47977));
    LocalMux I__10965 (
            .O(N__47992),
            .I(N__47977));
    LocalMux I__10964 (
            .O(N__47989),
            .I(N__47977));
    Span4Mux_h I__10963 (
            .O(N__47984),
            .I(N__47974));
    Span12Mux_v I__10962 (
            .O(N__47977),
            .I(N__47971));
    Span4Mux_v I__10961 (
            .O(N__47974),
            .I(N__47968));
    Span12Mux_h I__10960 (
            .O(N__47971),
            .I(N__47965));
    Sp12to4 I__10959 (
            .O(N__47968),
            .I(N__47962));
    Odrv12 I__10958 (
            .O(N__47965),
            .I(spi_select_c));
    Odrv12 I__10957 (
            .O(N__47962),
            .I(spi_select_c));
    InMux I__10956 (
            .O(N__47957),
            .I(N__47951));
    InMux I__10955 (
            .O(N__47956),
            .I(N__47951));
    LocalMux I__10954 (
            .O(N__47951),
            .I(N__47948));
    Span4Mux_h I__10953 (
            .O(N__47948),
            .I(N__47944));
    InMux I__10952 (
            .O(N__47947),
            .I(N__47941));
    Span4Mux_h I__10951 (
            .O(N__47944),
            .I(N__47936));
    LocalMux I__10950 (
            .O(N__47941),
            .I(N__47936));
    Span4Mux_v I__10949 (
            .O(N__47936),
            .I(N__47933));
    Span4Mux_h I__10948 (
            .O(N__47933),
            .I(N__47930));
    Span4Mux_v I__10947 (
            .O(N__47930),
            .I(N__47925));
    InMux I__10946 (
            .O(N__47929),
            .I(N__47922));
    InMux I__10945 (
            .O(N__47928),
            .I(N__47919));
    Sp12to4 I__10944 (
            .O(N__47925),
            .I(N__47912));
    LocalMux I__10943 (
            .O(N__47922),
            .I(N__47912));
    LocalMux I__10942 (
            .O(N__47919),
            .I(N__47912));
    Span12Mux_v I__10941 (
            .O(N__47912),
            .I(N__47909));
    Odrv12 I__10940 (
            .O(N__47909),
            .I(spi_cs_ft_c));
    CascadeMux I__10939 (
            .O(N__47906),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_ ));
    InMux I__10938 (
            .O(N__47903),
            .I(N__47900));
    LocalMux I__10937 (
            .O(N__47900),
            .I(N__47897));
    Span4Mux_v I__10936 (
            .O(N__47897),
            .I(N__47894));
    Span4Mux_h I__10935 (
            .O(N__47894),
            .I(N__47889));
    InMux I__10934 (
            .O(N__47893),
            .I(N__47882));
    InMux I__10933 (
            .O(N__47892),
            .I(N__47882));
    Span4Mux_h I__10932 (
            .O(N__47889),
            .I(N__47879));
    InMux I__10931 (
            .O(N__47888),
            .I(N__47876));
    InMux I__10930 (
            .O(N__47887),
            .I(N__47873));
    LocalMux I__10929 (
            .O(N__47882),
            .I(N__47870));
    Span4Mux_v I__10928 (
            .O(N__47879),
            .I(N__47867));
    LocalMux I__10927 (
            .O(N__47876),
            .I(N__47864));
    LocalMux I__10926 (
            .O(N__47873),
            .I(N__47861));
    Span12Mux_v I__10925 (
            .O(N__47870),
            .I(N__47858));
    Sp12to4 I__10924 (
            .O(N__47867),
            .I(N__47855));
    Span4Mux_h I__10923 (
            .O(N__47864),
            .I(N__47852));
    Span4Mux_h I__10922 (
            .O(N__47861),
            .I(N__47849));
    Span12Mux_v I__10921 (
            .O(N__47858),
            .I(N__47846));
    Span12Mux_s6_h I__10920 (
            .O(N__47855),
            .I(N__47839));
    Sp12to4 I__10919 (
            .O(N__47852),
            .I(N__47839));
    Sp12to4 I__10918 (
            .O(N__47849),
            .I(N__47839));
    Span12Mux_h I__10917 (
            .O(N__47846),
            .I(N__47834));
    Span12Mux_v I__10916 (
            .O(N__47839),
            .I(N__47834));
    Odrv12 I__10915 (
            .O(N__47834),
            .I(spi_cs_rpi_c));
    InMux I__10914 (
            .O(N__47831),
            .I(N__47828));
    LocalMux I__10913 (
            .O(N__47828),
            .I(N__47825));
    Span4Mux_v I__10912 (
            .O(N__47825),
            .I(N__47822));
    Span4Mux_v I__10911 (
            .O(N__47822),
            .I(N__47819));
    Odrv4 I__10910 (
            .O(N__47819),
            .I(\spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1 ));
    InMux I__10909 (
            .O(N__47816),
            .I(N__47813));
    LocalMux I__10908 (
            .O(N__47813),
            .I(N__47810));
    Span4Mux_v I__10907 (
            .O(N__47810),
            .I(N__47807));
    Span4Mux_v I__10906 (
            .O(N__47807),
            .I(N__47804));
    Odrv4 I__10905 (
            .O(N__47804),
            .I(\spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3 ));
    CascadeMux I__10904 (
            .O(N__47801),
            .I(\spi_slave_inst.N_1393_cascade_ ));
    IoInMux I__10903 (
            .O(N__47798),
            .I(N__47795));
    LocalMux I__10902 (
            .O(N__47795),
            .I(N__47792));
    IoSpan4Mux I__10901 (
            .O(N__47792),
            .I(N__47789));
    Span4Mux_s2_h I__10900 (
            .O(N__47789),
            .I(N__47786));
    Span4Mux_v I__10899 (
            .O(N__47786),
            .I(N__47783));
    Sp12to4 I__10898 (
            .O(N__47783),
            .I(N__47779));
    InMux I__10897 (
            .O(N__47782),
            .I(N__47776));
    Span12Mux_h I__10896 (
            .O(N__47779),
            .I(N__47773));
    LocalMux I__10895 (
            .O(N__47776),
            .I(N__47770));
    Odrv12 I__10894 (
            .O(N__47773),
            .I(spi_miso));
    Odrv12 I__10893 (
            .O(N__47770),
            .I(spi_miso));
    InMux I__10892 (
            .O(N__47765),
            .I(N__47762));
    LocalMux I__10891 (
            .O(N__47762),
            .I(N__47759));
    Span4Mux_v I__10890 (
            .O(N__47759),
            .I(N__47756));
    Odrv4 I__10889 (
            .O(N__47756),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_0 ));
    InMux I__10888 (
            .O(N__47753),
            .I(N__47750));
    LocalMux I__10887 (
            .O(N__47750),
            .I(N__47747));
    Span4Mux_v I__10886 (
            .O(N__47747),
            .I(N__47744));
    Odrv4 I__10885 (
            .O(N__47744),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_4 ));
    CascadeMux I__10884 (
            .O(N__47741),
            .I(\spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0_cascade_ ));
    InMux I__10883 (
            .O(N__47738),
            .I(N__47735));
    LocalMux I__10882 (
            .O(N__47735),
            .I(N__47732));
    Span4Mux_v I__10881 (
            .O(N__47732),
            .I(N__47729));
    Span4Mux_v I__10880 (
            .O(N__47729),
            .I(N__47726));
    Odrv4 I__10879 (
            .O(N__47726),
            .I(\spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2 ));
    InMux I__10878 (
            .O(N__47723),
            .I(N__47720));
    LocalMux I__10877 (
            .O(N__47720),
            .I(\spi_slave_inst.N_1396 ));
    InMux I__10876 (
            .O(N__47717),
            .I(N__47714));
    LocalMux I__10875 (
            .O(N__47714),
            .I(N__47711));
    Span12Mux_h I__10874 (
            .O(N__47711),
            .I(N__47708));
    Span12Mux_h I__10873 (
            .O(N__47708),
            .I(N__47705));
    Odrv12 I__10872 (
            .O(N__47705),
            .I(ADC7_c));
    IoInMux I__10871 (
            .O(N__47702),
            .I(N__47699));
    LocalMux I__10870 (
            .O(N__47699),
            .I(N__47696));
    IoSpan4Mux I__10869 (
            .O(N__47696),
            .I(N__47693));
    Span4Mux_s2_h I__10868 (
            .O(N__47693),
            .I(N__47690));
    Sp12to4 I__10867 (
            .O(N__47690),
            .I(N__47687));
    Span12Mux_s9_h I__10866 (
            .O(N__47687),
            .I(N__47684));
    Span12Mux_v I__10865 (
            .O(N__47684),
            .I(N__47681));
    Odrv12 I__10864 (
            .O(N__47681),
            .I(RAM_DATA_1Z0Z_8));
    InMux I__10863 (
            .O(N__47678),
            .I(N__47675));
    LocalMux I__10862 (
            .O(N__47675),
            .I(N__47672));
    Span4Mux_v I__10861 (
            .O(N__47672),
            .I(N__47669));
    Sp12to4 I__10860 (
            .O(N__47669),
            .I(N__47666));
    Span12Mux_h I__10859 (
            .O(N__47666),
            .I(N__47663));
    Span12Mux_h I__10858 (
            .O(N__47663),
            .I(N__47660));
    Odrv12 I__10857 (
            .O(N__47660),
            .I(ADC8_c));
    IoInMux I__10856 (
            .O(N__47657),
            .I(N__47654));
    LocalMux I__10855 (
            .O(N__47654),
            .I(N__47651));
    IoSpan4Mux I__10854 (
            .O(N__47651),
            .I(N__47648));
    IoSpan4Mux I__10853 (
            .O(N__47648),
            .I(N__47645));
    Sp12to4 I__10852 (
            .O(N__47645),
            .I(N__47642));
    Span12Mux_s9_h I__10851 (
            .O(N__47642),
            .I(N__47639));
    Odrv12 I__10850 (
            .O(N__47639),
            .I(RAM_DATA_1Z0Z_9));
    InMux I__10849 (
            .O(N__47636),
            .I(N__47633));
    LocalMux I__10848 (
            .O(N__47633),
            .I(N__47630));
    Span12Mux_h I__10847 (
            .O(N__47630),
            .I(N__47627));
    Span12Mux_h I__10846 (
            .O(N__47627),
            .I(N__47624));
    Span12Mux_v I__10845 (
            .O(N__47624),
            .I(N__47621));
    Odrv12 I__10844 (
            .O(N__47621),
            .I(top_tour2_c));
    IoInMux I__10843 (
            .O(N__47618),
            .I(N__47615));
    LocalMux I__10842 (
            .O(N__47615),
            .I(N__47612));
    IoSpan4Mux I__10841 (
            .O(N__47612),
            .I(N__47609));
    Sp12to4 I__10840 (
            .O(N__47609),
            .I(N__47606));
    Span12Mux_s9_h I__10839 (
            .O(N__47606),
            .I(N__47603));
    Odrv12 I__10838 (
            .O(N__47603),
            .I(RAM_DATA_1Z0Z_12));
    IoInMux I__10837 (
            .O(N__47600),
            .I(N__47597));
    LocalMux I__10836 (
            .O(N__47597),
            .I(N__47594));
    Span4Mux_s0_v I__10835 (
            .O(N__47594),
            .I(N__47591));
    Span4Mux_v I__10834 (
            .O(N__47591),
            .I(N__47588));
    Span4Mux_v I__10833 (
            .O(N__47588),
            .I(N__47585));
    Odrv4 I__10832 (
            .O(N__47585),
            .I(spi_miso_ft_c));
    InMux I__10831 (
            .O(N__47582),
            .I(N__47579));
    LocalMux I__10830 (
            .O(N__47579),
            .I(N__47576));
    Span4Mux_h I__10829 (
            .O(N__47576),
            .I(N__47573));
    Span4Mux_h I__10828 (
            .O(N__47573),
            .I(N__47570));
    Odrv4 I__10827 (
            .O(N__47570),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_8 ));
    InMux I__10826 (
            .O(N__47567),
            .I(N__47564));
    LocalMux I__10825 (
            .O(N__47564),
            .I(N__47561));
    Span12Mux_h I__10824 (
            .O(N__47561),
            .I(N__47558));
    Odrv12 I__10823 (
            .O(N__47558),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8 ));
    InMux I__10822 (
            .O(N__47555),
            .I(N__47549));
    InMux I__10821 (
            .O(N__47554),
            .I(N__47549));
    LocalMux I__10820 (
            .O(N__47549),
            .I(N__47546));
    Span4Mux_v I__10819 (
            .O(N__47546),
            .I(N__47542));
    CascadeMux I__10818 (
            .O(N__47545),
            .I(N__47539));
    Sp12to4 I__10817 (
            .O(N__47542),
            .I(N__47536));
    InMux I__10816 (
            .O(N__47539),
            .I(N__47533));
    Span12Mux_h I__10815 (
            .O(N__47536),
            .I(N__47530));
    LocalMux I__10814 (
            .O(N__47533),
            .I(sDAC_spi_startZ0));
    Odrv12 I__10813 (
            .O(N__47530),
            .I(sDAC_spi_startZ0));
    InMux I__10812 (
            .O(N__47525),
            .I(N__47522));
    LocalMux I__10811 (
            .O(N__47522),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_5 ));
    InMux I__10810 (
            .O(N__47519),
            .I(N__47516));
    LocalMux I__10809 (
            .O(N__47516),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_5 ));
    InMux I__10808 (
            .O(N__47513),
            .I(N__47508));
    InMux I__10807 (
            .O(N__47512),
            .I(N__47503));
    InMux I__10806 (
            .O(N__47511),
            .I(N__47493));
    LocalMux I__10805 (
            .O(N__47508),
            .I(N__47489));
    InMux I__10804 (
            .O(N__47507),
            .I(N__47486));
    InMux I__10803 (
            .O(N__47506),
            .I(N__47477));
    LocalMux I__10802 (
            .O(N__47503),
            .I(N__47474));
    InMux I__10801 (
            .O(N__47502),
            .I(N__47471));
    InMux I__10800 (
            .O(N__47501),
            .I(N__47468));
    InMux I__10799 (
            .O(N__47500),
            .I(N__47465));
    InMux I__10798 (
            .O(N__47499),
            .I(N__47462));
    InMux I__10797 (
            .O(N__47498),
            .I(N__47454));
    InMux I__10796 (
            .O(N__47497),
            .I(N__47451));
    InMux I__10795 (
            .O(N__47496),
            .I(N__47448));
    LocalMux I__10794 (
            .O(N__47493),
            .I(N__47443));
    InMux I__10793 (
            .O(N__47492),
            .I(N__47440));
    Span4Mux_v I__10792 (
            .O(N__47489),
            .I(N__47432));
    LocalMux I__10791 (
            .O(N__47486),
            .I(N__47432));
    InMux I__10790 (
            .O(N__47485),
            .I(N__47429));
    InMux I__10789 (
            .O(N__47484),
            .I(N__47426));
    InMux I__10788 (
            .O(N__47483),
            .I(N__47423));
    InMux I__10787 (
            .O(N__47482),
            .I(N__47420));
    InMux I__10786 (
            .O(N__47481),
            .I(N__47417));
    InMux I__10785 (
            .O(N__47480),
            .I(N__47414));
    LocalMux I__10784 (
            .O(N__47477),
            .I(N__47410));
    Span4Mux_v I__10783 (
            .O(N__47474),
            .I(N__47399));
    LocalMux I__10782 (
            .O(N__47471),
            .I(N__47399));
    LocalMux I__10781 (
            .O(N__47468),
            .I(N__47399));
    LocalMux I__10780 (
            .O(N__47465),
            .I(N__47399));
    LocalMux I__10779 (
            .O(N__47462),
            .I(N__47399));
    InMux I__10778 (
            .O(N__47461),
            .I(N__47396));
    InMux I__10777 (
            .O(N__47460),
            .I(N__47390));
    InMux I__10776 (
            .O(N__47459),
            .I(N__47387));
    InMux I__10775 (
            .O(N__47458),
            .I(N__47384));
    InMux I__10774 (
            .O(N__47457),
            .I(N__47381));
    LocalMux I__10773 (
            .O(N__47454),
            .I(N__47374));
    LocalMux I__10772 (
            .O(N__47451),
            .I(N__47374));
    LocalMux I__10771 (
            .O(N__47448),
            .I(N__47371));
    InMux I__10770 (
            .O(N__47447),
            .I(N__47368));
    InMux I__10769 (
            .O(N__47446),
            .I(N__47365));
    Span4Mux_v I__10768 (
            .O(N__47443),
            .I(N__47358));
    LocalMux I__10767 (
            .O(N__47440),
            .I(N__47358));
    InMux I__10766 (
            .O(N__47439),
            .I(N__47355));
    InMux I__10765 (
            .O(N__47438),
            .I(N__47352));
    InMux I__10764 (
            .O(N__47437),
            .I(N__47349));
    Span4Mux_v I__10763 (
            .O(N__47432),
            .I(N__47330));
    LocalMux I__10762 (
            .O(N__47429),
            .I(N__47330));
    LocalMux I__10761 (
            .O(N__47426),
            .I(N__47330));
    LocalMux I__10760 (
            .O(N__47423),
            .I(N__47330));
    LocalMux I__10759 (
            .O(N__47420),
            .I(N__47330));
    LocalMux I__10758 (
            .O(N__47417),
            .I(N__47330));
    LocalMux I__10757 (
            .O(N__47414),
            .I(N__47325));
    InMux I__10756 (
            .O(N__47413),
            .I(N__47322));
    Span4Mux_h I__10755 (
            .O(N__47410),
            .I(N__47315));
    Span4Mux_v I__10754 (
            .O(N__47399),
            .I(N__47315));
    LocalMux I__10753 (
            .O(N__47396),
            .I(N__47315));
    InMux I__10752 (
            .O(N__47395),
            .I(N__47312));
    InMux I__10751 (
            .O(N__47394),
            .I(N__47309));
    InMux I__10750 (
            .O(N__47393),
            .I(N__47306));
    LocalMux I__10749 (
            .O(N__47390),
            .I(N__47301));
    LocalMux I__10748 (
            .O(N__47387),
            .I(N__47301));
    LocalMux I__10747 (
            .O(N__47384),
            .I(N__47298));
    LocalMux I__10746 (
            .O(N__47381),
            .I(N__47295));
    InMux I__10745 (
            .O(N__47380),
            .I(N__47292));
    InMux I__10744 (
            .O(N__47379),
            .I(N__47289));
    Span4Mux_h I__10743 (
            .O(N__47374),
            .I(N__47282));
    Span4Mux_v I__10742 (
            .O(N__47371),
            .I(N__47282));
    LocalMux I__10741 (
            .O(N__47368),
            .I(N__47282));
    LocalMux I__10740 (
            .O(N__47365),
            .I(N__47279));
    InMux I__10739 (
            .O(N__47364),
            .I(N__47276));
    InMux I__10738 (
            .O(N__47363),
            .I(N__47272));
    Span4Mux_v I__10737 (
            .O(N__47358),
            .I(N__47267));
    LocalMux I__10736 (
            .O(N__47355),
            .I(N__47267));
    LocalMux I__10735 (
            .O(N__47352),
            .I(N__47264));
    LocalMux I__10734 (
            .O(N__47349),
            .I(N__47261));
    InMux I__10733 (
            .O(N__47348),
            .I(N__47258));
    InMux I__10732 (
            .O(N__47347),
            .I(N__47255));
    InMux I__10731 (
            .O(N__47346),
            .I(N__47252));
    InMux I__10730 (
            .O(N__47345),
            .I(N__47248));
    InMux I__10729 (
            .O(N__47344),
            .I(N__47241));
    InMux I__10728 (
            .O(N__47343),
            .I(N__47238));
    Span4Mux_v I__10727 (
            .O(N__47330),
            .I(N__47235));
    InMux I__10726 (
            .O(N__47329),
            .I(N__47232));
    InMux I__10725 (
            .O(N__47328),
            .I(N__47229));
    Span4Mux_v I__10724 (
            .O(N__47325),
            .I(N__47224));
    LocalMux I__10723 (
            .O(N__47322),
            .I(N__47224));
    Span4Mux_v I__10722 (
            .O(N__47315),
            .I(N__47215));
    LocalMux I__10721 (
            .O(N__47312),
            .I(N__47215));
    LocalMux I__10720 (
            .O(N__47309),
            .I(N__47215));
    LocalMux I__10719 (
            .O(N__47306),
            .I(N__47215));
    Span4Mux_v I__10718 (
            .O(N__47301),
            .I(N__47210));
    Span4Mux_v I__10717 (
            .O(N__47298),
            .I(N__47210));
    Span4Mux_v I__10716 (
            .O(N__47295),
            .I(N__47203));
    LocalMux I__10715 (
            .O(N__47292),
            .I(N__47203));
    LocalMux I__10714 (
            .O(N__47289),
            .I(N__47203));
    Span4Mux_v I__10713 (
            .O(N__47282),
            .I(N__47195));
    Span4Mux_h I__10712 (
            .O(N__47279),
            .I(N__47195));
    LocalMux I__10711 (
            .O(N__47276),
            .I(N__47195));
    InMux I__10710 (
            .O(N__47275),
            .I(N__47192));
    LocalMux I__10709 (
            .O(N__47272),
            .I(N__47189));
    Span4Mux_v I__10708 (
            .O(N__47267),
            .I(N__47178));
    Span4Mux_v I__10707 (
            .O(N__47264),
            .I(N__47178));
    Span4Mux_h I__10706 (
            .O(N__47261),
            .I(N__47178));
    LocalMux I__10705 (
            .O(N__47258),
            .I(N__47178));
    LocalMux I__10704 (
            .O(N__47255),
            .I(N__47178));
    LocalMux I__10703 (
            .O(N__47252),
            .I(N__47175));
    InMux I__10702 (
            .O(N__47251),
            .I(N__47171));
    LocalMux I__10701 (
            .O(N__47248),
            .I(N__47166));
    InMux I__10700 (
            .O(N__47247),
            .I(N__47163));
    InMux I__10699 (
            .O(N__47246),
            .I(N__47160));
    InMux I__10698 (
            .O(N__47245),
            .I(N__47157));
    InMux I__10697 (
            .O(N__47244),
            .I(N__47154));
    LocalMux I__10696 (
            .O(N__47241),
            .I(N__47149));
    LocalMux I__10695 (
            .O(N__47238),
            .I(N__47149));
    Sp12to4 I__10694 (
            .O(N__47235),
            .I(N__47144));
    LocalMux I__10693 (
            .O(N__47232),
            .I(N__47144));
    LocalMux I__10692 (
            .O(N__47229),
            .I(N__47141));
    Span4Mux_v I__10691 (
            .O(N__47224),
            .I(N__47138));
    Span4Mux_v I__10690 (
            .O(N__47215),
            .I(N__47135));
    Span4Mux_h I__10689 (
            .O(N__47210),
            .I(N__47130));
    Span4Mux_v I__10688 (
            .O(N__47203),
            .I(N__47130));
    InMux I__10687 (
            .O(N__47202),
            .I(N__47127));
    Span4Mux_h I__10686 (
            .O(N__47195),
            .I(N__47122));
    LocalMux I__10685 (
            .O(N__47192),
            .I(N__47122));
    Span4Mux_v I__10684 (
            .O(N__47189),
            .I(N__47115));
    Span4Mux_h I__10683 (
            .O(N__47178),
            .I(N__47110));
    Span4Mux_v I__10682 (
            .O(N__47175),
            .I(N__47110));
    InMux I__10681 (
            .O(N__47174),
            .I(N__47107));
    LocalMux I__10680 (
            .O(N__47171),
            .I(N__47104));
    InMux I__10679 (
            .O(N__47170),
            .I(N__47101));
    InMux I__10678 (
            .O(N__47169),
            .I(N__47098));
    Span4Mux_h I__10677 (
            .O(N__47166),
            .I(N__47087));
    LocalMux I__10676 (
            .O(N__47163),
            .I(N__47087));
    LocalMux I__10675 (
            .O(N__47160),
            .I(N__47087));
    LocalMux I__10674 (
            .O(N__47157),
            .I(N__47087));
    LocalMux I__10673 (
            .O(N__47154),
            .I(N__47087));
    Span12Mux_v I__10672 (
            .O(N__47149),
            .I(N__47080));
    Span12Mux_h I__10671 (
            .O(N__47144),
            .I(N__47080));
    Span12Mux_s10_v I__10670 (
            .O(N__47141),
            .I(N__47080));
    Span4Mux_v I__10669 (
            .O(N__47138),
            .I(N__47075));
    Span4Mux_v I__10668 (
            .O(N__47135),
            .I(N__47075));
    Span4Mux_v I__10667 (
            .O(N__47130),
            .I(N__47070));
    LocalMux I__10666 (
            .O(N__47127),
            .I(N__47070));
    Span4Mux_h I__10665 (
            .O(N__47122),
            .I(N__47067));
    InMux I__10664 (
            .O(N__47121),
            .I(N__47064));
    InMux I__10663 (
            .O(N__47120),
            .I(N__47061));
    InMux I__10662 (
            .O(N__47119),
            .I(N__47058));
    InMux I__10661 (
            .O(N__47118),
            .I(N__47055));
    Span4Mux_v I__10660 (
            .O(N__47115),
            .I(N__47048));
    Span4Mux_h I__10659 (
            .O(N__47110),
            .I(N__47048));
    LocalMux I__10658 (
            .O(N__47107),
            .I(N__47048));
    Span4Mux_v I__10657 (
            .O(N__47104),
            .I(N__47039));
    LocalMux I__10656 (
            .O(N__47101),
            .I(N__47039));
    LocalMux I__10655 (
            .O(N__47098),
            .I(N__47039));
    Span4Mux_v I__10654 (
            .O(N__47087),
            .I(N__47039));
    Odrv12 I__10653 (
            .O(N__47080),
            .I(spi_data_mosi_2));
    Odrv4 I__10652 (
            .O(N__47075),
            .I(spi_data_mosi_2));
    Odrv4 I__10651 (
            .O(N__47070),
            .I(spi_data_mosi_2));
    Odrv4 I__10650 (
            .O(N__47067),
            .I(spi_data_mosi_2));
    LocalMux I__10649 (
            .O(N__47064),
            .I(spi_data_mosi_2));
    LocalMux I__10648 (
            .O(N__47061),
            .I(spi_data_mosi_2));
    LocalMux I__10647 (
            .O(N__47058),
            .I(spi_data_mosi_2));
    LocalMux I__10646 (
            .O(N__47055),
            .I(spi_data_mosi_2));
    Odrv4 I__10645 (
            .O(N__47048),
            .I(spi_data_mosi_2));
    Odrv4 I__10644 (
            .O(N__47039),
            .I(spi_data_mosi_2));
    InMux I__10643 (
            .O(N__47018),
            .I(N__47014));
    InMux I__10642 (
            .O(N__47017),
            .I(N__47011));
    LocalMux I__10641 (
            .O(N__47014),
            .I(sCounterADCZ0Z_2));
    LocalMux I__10640 (
            .O(N__47011),
            .I(sCounterADCZ0Z_2));
    InMux I__10639 (
            .O(N__47006),
            .I(N__47003));
    LocalMux I__10638 (
            .O(N__47003),
            .I(sEEADC_freqZ0Z_2));
    InMux I__10637 (
            .O(N__47000),
            .I(N__46996));
    InMux I__10636 (
            .O(N__46999),
            .I(N__46993));
    LocalMux I__10635 (
            .O(N__46996),
            .I(sCounterADCZ0Z_3));
    LocalMux I__10634 (
            .O(N__46993),
            .I(sCounterADCZ0Z_3));
    InMux I__10633 (
            .O(N__46988),
            .I(N__46985));
    LocalMux I__10632 (
            .O(N__46985),
            .I(N__46982));
    Span12Mux_v I__10631 (
            .O(N__46982),
            .I(N__46979));
    Span12Mux_h I__10630 (
            .O(N__46979),
            .I(N__46976));
    Odrv12 I__10629 (
            .O(N__46976),
            .I(un11_sacqtime_NE_3));
    CascadeMux I__10628 (
            .O(N__46973),
            .I(un11_sacqtime_NE_0_0_cascade_));
    CascadeMux I__10627 (
            .O(N__46970),
            .I(N__46967));
    InMux I__10626 (
            .O(N__46967),
            .I(N__46964));
    LocalMux I__10625 (
            .O(N__46964),
            .I(N__46953));
    InMux I__10624 (
            .O(N__46963),
            .I(N__46944));
    InMux I__10623 (
            .O(N__46962),
            .I(N__46944));
    InMux I__10622 (
            .O(N__46961),
            .I(N__46944));
    InMux I__10621 (
            .O(N__46960),
            .I(N__46944));
    InMux I__10620 (
            .O(N__46959),
            .I(N__46935));
    InMux I__10619 (
            .O(N__46958),
            .I(N__46935));
    InMux I__10618 (
            .O(N__46957),
            .I(N__46935));
    InMux I__10617 (
            .O(N__46956),
            .I(N__46935));
    Span4Mux_h I__10616 (
            .O(N__46953),
            .I(N__46932));
    LocalMux I__10615 (
            .O(N__46944),
            .I(un11_sacqtime_NE_0));
    LocalMux I__10614 (
            .O(N__46935),
            .I(un11_sacqtime_NE_0));
    Odrv4 I__10613 (
            .O(N__46932),
            .I(un11_sacqtime_NE_0));
    InMux I__10612 (
            .O(N__46925),
            .I(N__46916));
    InMux I__10611 (
            .O(N__46924),
            .I(N__46910));
    InMux I__10610 (
            .O(N__46923),
            .I(N__46902));
    InMux I__10609 (
            .O(N__46922),
            .I(N__46898));
    InMux I__10608 (
            .O(N__46921),
            .I(N__46895));
    InMux I__10607 (
            .O(N__46920),
            .I(N__46892));
    InMux I__10606 (
            .O(N__46919),
            .I(N__46888));
    LocalMux I__10605 (
            .O(N__46916),
            .I(N__46885));
    InMux I__10604 (
            .O(N__46915),
            .I(N__46882));
    InMux I__10603 (
            .O(N__46914),
            .I(N__46879));
    InMux I__10602 (
            .O(N__46913),
            .I(N__46876));
    LocalMux I__10601 (
            .O(N__46910),
            .I(N__46873));
    InMux I__10600 (
            .O(N__46909),
            .I(N__46870));
    InMux I__10599 (
            .O(N__46908),
            .I(N__46867));
    InMux I__10598 (
            .O(N__46907),
            .I(N__46863));
    InMux I__10597 (
            .O(N__46906),
            .I(N__46860));
    InMux I__10596 (
            .O(N__46905),
            .I(N__46848));
    LocalMux I__10595 (
            .O(N__46902),
            .I(N__46844));
    InMux I__10594 (
            .O(N__46901),
            .I(N__46841));
    LocalMux I__10593 (
            .O(N__46898),
            .I(N__46833));
    LocalMux I__10592 (
            .O(N__46895),
            .I(N__46833));
    LocalMux I__10591 (
            .O(N__46892),
            .I(N__46833));
    InMux I__10590 (
            .O(N__46891),
            .I(N__46830));
    LocalMux I__10589 (
            .O(N__46888),
            .I(N__46826));
    Span4Mux_v I__10588 (
            .O(N__46885),
            .I(N__46817));
    LocalMux I__10587 (
            .O(N__46882),
            .I(N__46817));
    LocalMux I__10586 (
            .O(N__46879),
            .I(N__46817));
    LocalMux I__10585 (
            .O(N__46876),
            .I(N__46817));
    Span4Mux_h I__10584 (
            .O(N__46873),
            .I(N__46810));
    LocalMux I__10583 (
            .O(N__46870),
            .I(N__46810));
    LocalMux I__10582 (
            .O(N__46867),
            .I(N__46810));
    InMux I__10581 (
            .O(N__46866),
            .I(N__46807));
    LocalMux I__10580 (
            .O(N__46863),
            .I(N__46804));
    LocalMux I__10579 (
            .O(N__46860),
            .I(N__46801));
    InMux I__10578 (
            .O(N__46859),
            .I(N__46798));
    InMux I__10577 (
            .O(N__46858),
            .I(N__46795));
    InMux I__10576 (
            .O(N__46857),
            .I(N__46790));
    InMux I__10575 (
            .O(N__46856),
            .I(N__46786));
    InMux I__10574 (
            .O(N__46855),
            .I(N__46783));
    InMux I__10573 (
            .O(N__46854),
            .I(N__46780));
    InMux I__10572 (
            .O(N__46853),
            .I(N__46776));
    InMux I__10571 (
            .O(N__46852),
            .I(N__46771));
    InMux I__10570 (
            .O(N__46851),
            .I(N__46766));
    LocalMux I__10569 (
            .O(N__46848),
            .I(N__46759));
    InMux I__10568 (
            .O(N__46847),
            .I(N__46756));
    Span4Mux_v I__10567 (
            .O(N__46844),
            .I(N__46753));
    LocalMux I__10566 (
            .O(N__46841),
            .I(N__46747));
    InMux I__10565 (
            .O(N__46840),
            .I(N__46743));
    Span4Mux_h I__10564 (
            .O(N__46833),
            .I(N__46738));
    LocalMux I__10563 (
            .O(N__46830),
            .I(N__46738));
    InMux I__10562 (
            .O(N__46829),
            .I(N__46735));
    Span4Mux_h I__10561 (
            .O(N__46826),
            .I(N__46726));
    Span4Mux_h I__10560 (
            .O(N__46817),
            .I(N__46726));
    Span4Mux_v I__10559 (
            .O(N__46810),
            .I(N__46726));
    LocalMux I__10558 (
            .O(N__46807),
            .I(N__46726));
    Span4Mux_v I__10557 (
            .O(N__46804),
            .I(N__46719));
    Span4Mux_h I__10556 (
            .O(N__46801),
            .I(N__46719));
    LocalMux I__10555 (
            .O(N__46798),
            .I(N__46719));
    LocalMux I__10554 (
            .O(N__46795),
            .I(N__46716));
    InMux I__10553 (
            .O(N__46794),
            .I(N__46713));
    InMux I__10552 (
            .O(N__46793),
            .I(N__46710));
    LocalMux I__10551 (
            .O(N__46790),
            .I(N__46704));
    InMux I__10550 (
            .O(N__46789),
            .I(N__46701));
    LocalMux I__10549 (
            .O(N__46786),
            .I(N__46696));
    LocalMux I__10548 (
            .O(N__46783),
            .I(N__46696));
    LocalMux I__10547 (
            .O(N__46780),
            .I(N__46693));
    InMux I__10546 (
            .O(N__46779),
            .I(N__46690));
    LocalMux I__10545 (
            .O(N__46776),
            .I(N__46686));
    InMux I__10544 (
            .O(N__46775),
            .I(N__46683));
    InMux I__10543 (
            .O(N__46774),
            .I(N__46680));
    LocalMux I__10542 (
            .O(N__46771),
            .I(N__46677));
    InMux I__10541 (
            .O(N__46770),
            .I(N__46674));
    InMux I__10540 (
            .O(N__46769),
            .I(N__46671));
    LocalMux I__10539 (
            .O(N__46766),
            .I(N__46668));
    InMux I__10538 (
            .O(N__46765),
            .I(N__46665));
    InMux I__10537 (
            .O(N__46764),
            .I(N__46662));
    InMux I__10536 (
            .O(N__46763),
            .I(N__46659));
    InMux I__10535 (
            .O(N__46762),
            .I(N__46656));
    Span4Mux_h I__10534 (
            .O(N__46759),
            .I(N__46651));
    LocalMux I__10533 (
            .O(N__46756),
            .I(N__46651));
    Span4Mux_v I__10532 (
            .O(N__46753),
            .I(N__46647));
    InMux I__10531 (
            .O(N__46752),
            .I(N__46644));
    InMux I__10530 (
            .O(N__46751),
            .I(N__46641));
    InMux I__10529 (
            .O(N__46750),
            .I(N__46638));
    Span4Mux_v I__10528 (
            .O(N__46747),
            .I(N__46635));
    InMux I__10527 (
            .O(N__46746),
            .I(N__46632));
    LocalMux I__10526 (
            .O(N__46743),
            .I(N__46629));
    Span4Mux_h I__10525 (
            .O(N__46738),
            .I(N__46624));
    LocalMux I__10524 (
            .O(N__46735),
            .I(N__46624));
    Span4Mux_v I__10523 (
            .O(N__46726),
            .I(N__46621));
    Span4Mux_v I__10522 (
            .O(N__46719),
            .I(N__46614));
    Span4Mux_h I__10521 (
            .O(N__46716),
            .I(N__46614));
    LocalMux I__10520 (
            .O(N__46713),
            .I(N__46614));
    LocalMux I__10519 (
            .O(N__46710),
            .I(N__46611));
    InMux I__10518 (
            .O(N__46709),
            .I(N__46608));
    InMux I__10517 (
            .O(N__46708),
            .I(N__46605));
    InMux I__10516 (
            .O(N__46707),
            .I(N__46600));
    Span4Mux_v I__10515 (
            .O(N__46704),
            .I(N__46593));
    LocalMux I__10514 (
            .O(N__46701),
            .I(N__46593));
    Span4Mux_h I__10513 (
            .O(N__46696),
            .I(N__46586));
    Span4Mux_v I__10512 (
            .O(N__46693),
            .I(N__46586));
    LocalMux I__10511 (
            .O(N__46690),
            .I(N__46586));
    InMux I__10510 (
            .O(N__46689),
            .I(N__46583));
    Span4Mux_h I__10509 (
            .O(N__46686),
            .I(N__46572));
    LocalMux I__10508 (
            .O(N__46683),
            .I(N__46572));
    LocalMux I__10507 (
            .O(N__46680),
            .I(N__46572));
    Span4Mux_h I__10506 (
            .O(N__46677),
            .I(N__46572));
    LocalMux I__10505 (
            .O(N__46674),
            .I(N__46572));
    LocalMux I__10504 (
            .O(N__46671),
            .I(N__46569));
    Span4Mux_h I__10503 (
            .O(N__46668),
            .I(N__46566));
    LocalMux I__10502 (
            .O(N__46665),
            .I(N__46557));
    LocalMux I__10501 (
            .O(N__46662),
            .I(N__46557));
    LocalMux I__10500 (
            .O(N__46659),
            .I(N__46557));
    LocalMux I__10499 (
            .O(N__46656),
            .I(N__46557));
    Span4Mux_h I__10498 (
            .O(N__46651),
            .I(N__46554));
    InMux I__10497 (
            .O(N__46650),
            .I(N__46551));
    Sp12to4 I__10496 (
            .O(N__46647),
            .I(N__46538));
    LocalMux I__10495 (
            .O(N__46644),
            .I(N__46538));
    LocalMux I__10494 (
            .O(N__46641),
            .I(N__46538));
    LocalMux I__10493 (
            .O(N__46638),
            .I(N__46538));
    Sp12to4 I__10492 (
            .O(N__46635),
            .I(N__46538));
    LocalMux I__10491 (
            .O(N__46632),
            .I(N__46538));
    Span4Mux_h I__10490 (
            .O(N__46629),
            .I(N__46533));
    Span4Mux_h I__10489 (
            .O(N__46624),
            .I(N__46533));
    Span4Mux_v I__10488 (
            .O(N__46621),
            .I(N__46522));
    Span4Mux_h I__10487 (
            .O(N__46614),
            .I(N__46522));
    Span4Mux_v I__10486 (
            .O(N__46611),
            .I(N__46522));
    LocalMux I__10485 (
            .O(N__46608),
            .I(N__46522));
    LocalMux I__10484 (
            .O(N__46605),
            .I(N__46522));
    InMux I__10483 (
            .O(N__46604),
            .I(N__46515));
    InMux I__10482 (
            .O(N__46603),
            .I(N__46512));
    LocalMux I__10481 (
            .O(N__46600),
            .I(N__46509));
    InMux I__10480 (
            .O(N__46599),
            .I(N__46506));
    InMux I__10479 (
            .O(N__46598),
            .I(N__46503));
    Span4Mux_h I__10478 (
            .O(N__46593),
            .I(N__46494));
    Span4Mux_v I__10477 (
            .O(N__46586),
            .I(N__46494));
    LocalMux I__10476 (
            .O(N__46583),
            .I(N__46494));
    Span4Mux_v I__10475 (
            .O(N__46572),
            .I(N__46494));
    Span4Mux_h I__10474 (
            .O(N__46569),
            .I(N__46491));
    Sp12to4 I__10473 (
            .O(N__46566),
            .I(N__46478));
    Span12Mux_h I__10472 (
            .O(N__46557),
            .I(N__46478));
    Sp12to4 I__10471 (
            .O(N__46554),
            .I(N__46478));
    LocalMux I__10470 (
            .O(N__46551),
            .I(N__46478));
    Span12Mux_h I__10469 (
            .O(N__46538),
            .I(N__46478));
    Sp12to4 I__10468 (
            .O(N__46533),
            .I(N__46478));
    Span4Mux_h I__10467 (
            .O(N__46522),
            .I(N__46475));
    InMux I__10466 (
            .O(N__46521),
            .I(N__46472));
    InMux I__10465 (
            .O(N__46520),
            .I(N__46469));
    InMux I__10464 (
            .O(N__46519),
            .I(N__46466));
    InMux I__10463 (
            .O(N__46518),
            .I(N__46463));
    LocalMux I__10462 (
            .O(N__46515),
            .I(N__46458));
    LocalMux I__10461 (
            .O(N__46512),
            .I(N__46458));
    Span4Mux_v I__10460 (
            .O(N__46509),
            .I(N__46449));
    LocalMux I__10459 (
            .O(N__46506),
            .I(N__46449));
    LocalMux I__10458 (
            .O(N__46503),
            .I(N__46449));
    Span4Mux_h I__10457 (
            .O(N__46494),
            .I(N__46449));
    Odrv4 I__10456 (
            .O(N__46491),
            .I(spi_data_mosi_3));
    Odrv12 I__10455 (
            .O(N__46478),
            .I(spi_data_mosi_3));
    Odrv4 I__10454 (
            .O(N__46475),
            .I(spi_data_mosi_3));
    LocalMux I__10453 (
            .O(N__46472),
            .I(spi_data_mosi_3));
    LocalMux I__10452 (
            .O(N__46469),
            .I(spi_data_mosi_3));
    LocalMux I__10451 (
            .O(N__46466),
            .I(spi_data_mosi_3));
    LocalMux I__10450 (
            .O(N__46463),
            .I(spi_data_mosi_3));
    Odrv4 I__10449 (
            .O(N__46458),
            .I(spi_data_mosi_3));
    Odrv4 I__10448 (
            .O(N__46449),
            .I(spi_data_mosi_3));
    CascadeMux I__10447 (
            .O(N__46430),
            .I(N__46427));
    InMux I__10446 (
            .O(N__46427),
            .I(N__46424));
    LocalMux I__10445 (
            .O(N__46424),
            .I(sEEADC_freqZ0Z_3));
    InMux I__10444 (
            .O(N__46421),
            .I(N__46417));
    InMux I__10443 (
            .O(N__46420),
            .I(N__46414));
    LocalMux I__10442 (
            .O(N__46417),
            .I(sCounterADCZ0Z_1));
    LocalMux I__10441 (
            .O(N__46414),
            .I(sCounterADCZ0Z_1));
    InMux I__10440 (
            .O(N__46409),
            .I(N__46405));
    InMux I__10439 (
            .O(N__46408),
            .I(N__46402));
    LocalMux I__10438 (
            .O(N__46405),
            .I(sCounterADCZ0Z_0));
    LocalMux I__10437 (
            .O(N__46402),
            .I(sCounterADCZ0Z_0));
    InMux I__10436 (
            .O(N__46397),
            .I(N__46394));
    LocalMux I__10435 (
            .O(N__46394),
            .I(un11_sacqtime_NE_1));
    InMux I__10434 (
            .O(N__46391),
            .I(N__46376));
    InMux I__10433 (
            .O(N__46390),
            .I(N__46371));
    InMux I__10432 (
            .O(N__46389),
            .I(N__46368));
    InMux I__10431 (
            .O(N__46388),
            .I(N__46365));
    InMux I__10430 (
            .O(N__46387),
            .I(N__46362));
    InMux I__10429 (
            .O(N__46386),
            .I(N__46359));
    InMux I__10428 (
            .O(N__46385),
            .I(N__46356));
    InMux I__10427 (
            .O(N__46384),
            .I(N__46353));
    InMux I__10426 (
            .O(N__46383),
            .I(N__46349));
    InMux I__10425 (
            .O(N__46382),
            .I(N__46346));
    InMux I__10424 (
            .O(N__46381),
            .I(N__46339));
    InMux I__10423 (
            .O(N__46380),
            .I(N__46335));
    InMux I__10422 (
            .O(N__46379),
            .I(N__46332));
    LocalMux I__10421 (
            .O(N__46376),
            .I(N__46328));
    InMux I__10420 (
            .O(N__46375),
            .I(N__46325));
    InMux I__10419 (
            .O(N__46374),
            .I(N__46318));
    LocalMux I__10418 (
            .O(N__46371),
            .I(N__46309));
    LocalMux I__10417 (
            .O(N__46368),
            .I(N__46309));
    LocalMux I__10416 (
            .O(N__46365),
            .I(N__46300));
    LocalMux I__10415 (
            .O(N__46362),
            .I(N__46300));
    LocalMux I__10414 (
            .O(N__46359),
            .I(N__46300));
    LocalMux I__10413 (
            .O(N__46356),
            .I(N__46300));
    LocalMux I__10412 (
            .O(N__46353),
            .I(N__46297));
    InMux I__10411 (
            .O(N__46352),
            .I(N__46294));
    LocalMux I__10410 (
            .O(N__46349),
            .I(N__46288));
    LocalMux I__10409 (
            .O(N__46346),
            .I(N__46288));
    InMux I__10408 (
            .O(N__46345),
            .I(N__46285));
    InMux I__10407 (
            .O(N__46344),
            .I(N__46282));
    InMux I__10406 (
            .O(N__46343),
            .I(N__46276));
    InMux I__10405 (
            .O(N__46342),
            .I(N__46273));
    LocalMux I__10404 (
            .O(N__46339),
            .I(N__46270));
    InMux I__10403 (
            .O(N__46338),
            .I(N__46267));
    LocalMux I__10402 (
            .O(N__46335),
            .I(N__46262));
    LocalMux I__10401 (
            .O(N__46332),
            .I(N__46262));
    InMux I__10400 (
            .O(N__46331),
            .I(N__46259));
    Span4Mux_v I__10399 (
            .O(N__46328),
            .I(N__46254));
    LocalMux I__10398 (
            .O(N__46325),
            .I(N__46254));
    InMux I__10397 (
            .O(N__46324),
            .I(N__46251));
    InMux I__10396 (
            .O(N__46323),
            .I(N__46248));
    InMux I__10395 (
            .O(N__46322),
            .I(N__46245));
    InMux I__10394 (
            .O(N__46321),
            .I(N__46242));
    LocalMux I__10393 (
            .O(N__46318),
            .I(N__46239));
    InMux I__10392 (
            .O(N__46317),
            .I(N__46236));
    InMux I__10391 (
            .O(N__46316),
            .I(N__46230));
    InMux I__10390 (
            .O(N__46315),
            .I(N__46227));
    InMux I__10389 (
            .O(N__46314),
            .I(N__46224));
    Span4Mux_h I__10388 (
            .O(N__46309),
            .I(N__46215));
    Span4Mux_v I__10387 (
            .O(N__46300),
            .I(N__46215));
    Span4Mux_h I__10386 (
            .O(N__46297),
            .I(N__46215));
    LocalMux I__10385 (
            .O(N__46294),
            .I(N__46215));
    InMux I__10384 (
            .O(N__46293),
            .I(N__46212));
    Span4Mux_v I__10383 (
            .O(N__46288),
            .I(N__46202));
    LocalMux I__10382 (
            .O(N__46285),
            .I(N__46202));
    LocalMux I__10381 (
            .O(N__46282),
            .I(N__46202));
    InMux I__10380 (
            .O(N__46281),
            .I(N__46199));
    InMux I__10379 (
            .O(N__46280),
            .I(N__46196));
    InMux I__10378 (
            .O(N__46279),
            .I(N__46193));
    LocalMux I__10377 (
            .O(N__46276),
            .I(N__46184));
    LocalMux I__10376 (
            .O(N__46273),
            .I(N__46184));
    Span4Mux_h I__10375 (
            .O(N__46270),
            .I(N__46184));
    LocalMux I__10374 (
            .O(N__46267),
            .I(N__46184));
    Span4Mux_v I__10373 (
            .O(N__46262),
            .I(N__46179));
    LocalMux I__10372 (
            .O(N__46259),
            .I(N__46179));
    Span4Mux_h I__10371 (
            .O(N__46254),
            .I(N__46174));
    LocalMux I__10370 (
            .O(N__46251),
            .I(N__46174));
    LocalMux I__10369 (
            .O(N__46248),
            .I(N__46167));
    LocalMux I__10368 (
            .O(N__46245),
            .I(N__46167));
    LocalMux I__10367 (
            .O(N__46242),
            .I(N__46167));
    Span4Mux_h I__10366 (
            .O(N__46239),
            .I(N__46162));
    LocalMux I__10365 (
            .O(N__46236),
            .I(N__46162));
    InMux I__10364 (
            .O(N__46235),
            .I(N__46159));
    InMux I__10363 (
            .O(N__46234),
            .I(N__46156));
    InMux I__10362 (
            .O(N__46233),
            .I(N__46153));
    LocalMux I__10361 (
            .O(N__46230),
            .I(N__46150));
    LocalMux I__10360 (
            .O(N__46227),
            .I(N__46136));
    LocalMux I__10359 (
            .O(N__46224),
            .I(N__46136));
    Span4Mux_v I__10358 (
            .O(N__46215),
            .I(N__46131));
    LocalMux I__10357 (
            .O(N__46212),
            .I(N__46131));
    CascadeMux I__10356 (
            .O(N__46211),
            .I(N__46127));
    InMux I__10355 (
            .O(N__46210),
            .I(N__46124));
    InMux I__10354 (
            .O(N__46209),
            .I(N__46121));
    Span4Mux_h I__10353 (
            .O(N__46202),
            .I(N__46118));
    LocalMux I__10352 (
            .O(N__46199),
            .I(N__46115));
    LocalMux I__10351 (
            .O(N__46196),
            .I(N__46106));
    LocalMux I__10350 (
            .O(N__46193),
            .I(N__46106));
    Span4Mux_h I__10349 (
            .O(N__46184),
            .I(N__46106));
    Span4Mux_h I__10348 (
            .O(N__46179),
            .I(N__46106));
    Span4Mux_v I__10347 (
            .O(N__46174),
            .I(N__46101));
    Span4Mux_v I__10346 (
            .O(N__46167),
            .I(N__46101));
    Span4Mux_v I__10345 (
            .O(N__46162),
            .I(N__46098));
    LocalMux I__10344 (
            .O(N__46159),
            .I(N__46093));
    LocalMux I__10343 (
            .O(N__46156),
            .I(N__46093));
    LocalMux I__10342 (
            .O(N__46153),
            .I(N__46090));
    Span4Mux_v I__10341 (
            .O(N__46150),
            .I(N__46087));
    InMux I__10340 (
            .O(N__46149),
            .I(N__46084));
    InMux I__10339 (
            .O(N__46148),
            .I(N__46081));
    InMux I__10338 (
            .O(N__46147),
            .I(N__46078));
    InMux I__10337 (
            .O(N__46146),
            .I(N__46075));
    InMux I__10336 (
            .O(N__46145),
            .I(N__46072));
    InMux I__10335 (
            .O(N__46144),
            .I(N__46069));
    InMux I__10334 (
            .O(N__46143),
            .I(N__46066));
    InMux I__10333 (
            .O(N__46142),
            .I(N__46063));
    InMux I__10332 (
            .O(N__46141),
            .I(N__46060));
    Span4Mux_v I__10331 (
            .O(N__46136),
            .I(N__46055));
    Span4Mux_v I__10330 (
            .O(N__46131),
            .I(N__46055));
    InMux I__10329 (
            .O(N__46130),
            .I(N__46047));
    InMux I__10328 (
            .O(N__46127),
            .I(N__46044));
    LocalMux I__10327 (
            .O(N__46124),
            .I(N__46039));
    LocalMux I__10326 (
            .O(N__46121),
            .I(N__46034));
    Span4Mux_h I__10325 (
            .O(N__46118),
            .I(N__46034));
    Span4Mux_h I__10324 (
            .O(N__46115),
            .I(N__46029));
    Span4Mux_v I__10323 (
            .O(N__46106),
            .I(N__46029));
    Span4Mux_h I__10322 (
            .O(N__46101),
            .I(N__46022));
    Span4Mux_h I__10321 (
            .O(N__46098),
            .I(N__46022));
    Span4Mux_v I__10320 (
            .O(N__46093),
            .I(N__46022));
    Span4Mux_v I__10319 (
            .O(N__46090),
            .I(N__46019));
    Sp12to4 I__10318 (
            .O(N__46087),
            .I(N__46016));
    LocalMux I__10317 (
            .O(N__46084),
            .I(N__46010));
    LocalMux I__10316 (
            .O(N__46081),
            .I(N__46010));
    LocalMux I__10315 (
            .O(N__46078),
            .I(N__46005));
    LocalMux I__10314 (
            .O(N__46075),
            .I(N__46005));
    LocalMux I__10313 (
            .O(N__46072),
            .I(N__46002));
    LocalMux I__10312 (
            .O(N__46069),
            .I(N__45999));
    LocalMux I__10311 (
            .O(N__46066),
            .I(N__45990));
    LocalMux I__10310 (
            .O(N__46063),
            .I(N__45990));
    LocalMux I__10309 (
            .O(N__46060),
            .I(N__45990));
    Span4Mux_h I__10308 (
            .O(N__46055),
            .I(N__45990));
    InMux I__10307 (
            .O(N__46054),
            .I(N__45987));
    InMux I__10306 (
            .O(N__46053),
            .I(N__45980));
    InMux I__10305 (
            .O(N__46052),
            .I(N__45980));
    InMux I__10304 (
            .O(N__46051),
            .I(N__45980));
    InMux I__10303 (
            .O(N__46050),
            .I(N__45974));
    LocalMux I__10302 (
            .O(N__46047),
            .I(N__45969));
    LocalMux I__10301 (
            .O(N__46044),
            .I(N__45969));
    InMux I__10300 (
            .O(N__46043),
            .I(N__45966));
    InMux I__10299 (
            .O(N__46042),
            .I(N__45963));
    Span4Mux_h I__10298 (
            .O(N__46039),
            .I(N__45956));
    Span4Mux_h I__10297 (
            .O(N__46034),
            .I(N__45956));
    Span4Mux_v I__10296 (
            .O(N__46029),
            .I(N__45956));
    Sp12to4 I__10295 (
            .O(N__46022),
            .I(N__45953));
    Sp12to4 I__10294 (
            .O(N__46019),
            .I(N__45948));
    Span12Mux_v I__10293 (
            .O(N__46016),
            .I(N__45948));
    InMux I__10292 (
            .O(N__46015),
            .I(N__45945));
    Span4Mux_v I__10291 (
            .O(N__46010),
            .I(N__45942));
    Span4Mux_v I__10290 (
            .O(N__46005),
            .I(N__45935));
    Span4Mux_h I__10289 (
            .O(N__46002),
            .I(N__45935));
    Span4Mux_v I__10288 (
            .O(N__45999),
            .I(N__45935));
    Span4Mux_v I__10287 (
            .O(N__45990),
            .I(N__45932));
    LocalMux I__10286 (
            .O(N__45987),
            .I(N__45927));
    LocalMux I__10285 (
            .O(N__45980),
            .I(N__45927));
    InMux I__10284 (
            .O(N__45979),
            .I(N__45924));
    InMux I__10283 (
            .O(N__45978),
            .I(N__45921));
    InMux I__10282 (
            .O(N__45977),
            .I(N__45918));
    LocalMux I__10281 (
            .O(N__45974),
            .I(N__45911));
    Span4Mux_v I__10280 (
            .O(N__45969),
            .I(N__45911));
    LocalMux I__10279 (
            .O(N__45966),
            .I(N__45911));
    LocalMux I__10278 (
            .O(N__45963),
            .I(N__45908));
    Span4Mux_v I__10277 (
            .O(N__45956),
            .I(N__45905));
    Span12Mux_h I__10276 (
            .O(N__45953),
            .I(N__45900));
    Span12Mux_h I__10275 (
            .O(N__45948),
            .I(N__45900));
    LocalMux I__10274 (
            .O(N__45945),
            .I(N__45889));
    Span4Mux_v I__10273 (
            .O(N__45942),
            .I(N__45889));
    Span4Mux_h I__10272 (
            .O(N__45935),
            .I(N__45889));
    Span4Mux_h I__10271 (
            .O(N__45932),
            .I(N__45889));
    Span4Mux_h I__10270 (
            .O(N__45927),
            .I(N__45889));
    LocalMux I__10269 (
            .O(N__45924),
            .I(spi_data_mosi_0));
    LocalMux I__10268 (
            .O(N__45921),
            .I(spi_data_mosi_0));
    LocalMux I__10267 (
            .O(N__45918),
            .I(spi_data_mosi_0));
    Odrv4 I__10266 (
            .O(N__45911),
            .I(spi_data_mosi_0));
    Odrv4 I__10265 (
            .O(N__45908),
            .I(spi_data_mosi_0));
    Odrv4 I__10264 (
            .O(N__45905),
            .I(spi_data_mosi_0));
    Odrv12 I__10263 (
            .O(N__45900),
            .I(spi_data_mosi_0));
    Odrv4 I__10262 (
            .O(N__45889),
            .I(spi_data_mosi_0));
    InMux I__10261 (
            .O(N__45872),
            .I(N__45869));
    LocalMux I__10260 (
            .O(N__45869),
            .I(sEEADC_freqZ0Z_0));
    CascadeMux I__10259 (
            .O(N__45866),
            .I(N__45863));
    InMux I__10258 (
            .O(N__45863),
            .I(N__45860));
    LocalMux I__10257 (
            .O(N__45860),
            .I(sEEADC_freqZ0Z_1));
    InMux I__10256 (
            .O(N__45857),
            .I(N__45853));
    InMux I__10255 (
            .O(N__45856),
            .I(N__45850));
    LocalMux I__10254 (
            .O(N__45853),
            .I(sCounterADCZ0Z_7));
    LocalMux I__10253 (
            .O(N__45850),
            .I(sCounterADCZ0Z_7));
    CascadeMux I__10252 (
            .O(N__45845),
            .I(N__45841));
    InMux I__10251 (
            .O(N__45844),
            .I(N__45838));
    InMux I__10250 (
            .O(N__45841),
            .I(N__45835));
    LocalMux I__10249 (
            .O(N__45838),
            .I(sCounterADCZ0Z_6));
    LocalMux I__10248 (
            .O(N__45835),
            .I(sCounterADCZ0Z_6));
    InMux I__10247 (
            .O(N__45830),
            .I(N__45827));
    LocalMux I__10246 (
            .O(N__45827),
            .I(un11_sacqtime_NE_2));
    InMux I__10245 (
            .O(N__45824),
            .I(N__45821));
    LocalMux I__10244 (
            .O(N__45821),
            .I(N__45818));
    Odrv4 I__10243 (
            .O(N__45818),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_4 ));
    InMux I__10242 (
            .O(N__45815),
            .I(N__45812));
    LocalMux I__10241 (
            .O(N__45812),
            .I(N__45809));
    Odrv4 I__10240 (
            .O(N__45809),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_0 ));
    InMux I__10239 (
            .O(N__45806),
            .I(N__45803));
    LocalMux I__10238 (
            .O(N__45803),
            .I(N__45800));
    Odrv4 I__10237 (
            .O(N__45800),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_2 ));
    InMux I__10236 (
            .O(N__45797),
            .I(N__45794));
    LocalMux I__10235 (
            .O(N__45794),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_2 ));
    InMux I__10234 (
            .O(N__45791),
            .I(N__45788));
    LocalMux I__10233 (
            .O(N__45788),
            .I(N__45785));
    Odrv4 I__10232 (
            .O(N__45785),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_1 ));
    InMux I__10231 (
            .O(N__45782),
            .I(N__45779));
    LocalMux I__10230 (
            .O(N__45779),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_1 ));
    InMux I__10229 (
            .O(N__45776),
            .I(N__45773));
    LocalMux I__10228 (
            .O(N__45773),
            .I(N__45768));
    InMux I__10227 (
            .O(N__45772),
            .I(N__45765));
    InMux I__10226 (
            .O(N__45771),
            .I(N__45762));
    Span12Mux_h I__10225 (
            .O(N__45768),
            .I(N__45757));
    LocalMux I__10224 (
            .O(N__45765),
            .I(N__45757));
    LocalMux I__10223 (
            .O(N__45762),
            .I(button_debounce_counterZ0Z_1));
    Odrv12 I__10222 (
            .O(N__45757),
            .I(button_debounce_counterZ0Z_1));
    InMux I__10221 (
            .O(N__45752),
            .I(N__45748));
    CascadeMux I__10220 (
            .O(N__45751),
            .I(N__45745));
    LocalMux I__10219 (
            .O(N__45748),
            .I(N__45740));
    InMux I__10218 (
            .O(N__45745),
            .I(N__45737));
    InMux I__10217 (
            .O(N__45744),
            .I(N__45732));
    InMux I__10216 (
            .O(N__45743),
            .I(N__45732));
    Span12Mux_h I__10215 (
            .O(N__45740),
            .I(N__45727));
    LocalMux I__10214 (
            .O(N__45737),
            .I(N__45727));
    LocalMux I__10213 (
            .O(N__45732),
            .I(button_debounce_counterZ0Z_0));
    Odrv12 I__10212 (
            .O(N__45727),
            .I(button_debounce_counterZ0Z_0));
    InMux I__10211 (
            .O(N__45722),
            .I(N__45719));
    LocalMux I__10210 (
            .O(N__45719),
            .I(N__45711));
    SRMux I__10209 (
            .O(N__45718),
            .I(N__45698));
    SRMux I__10208 (
            .O(N__45717),
            .I(N__45698));
    SRMux I__10207 (
            .O(N__45716),
            .I(N__45698));
    SRMux I__10206 (
            .O(N__45715),
            .I(N__45698));
    SRMux I__10205 (
            .O(N__45714),
            .I(N__45698));
    Glb2LocalMux I__10204 (
            .O(N__45711),
            .I(N__45698));
    GlobalMux I__10203 (
            .O(N__45698),
            .I(N__45695));
    gio2CtrlBuf I__10202 (
            .O(N__45695),
            .I(N_3154_g));
    InMux I__10201 (
            .O(N__45692),
            .I(N__45689));
    LocalMux I__10200 (
            .O(N__45689),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_3 ));
    InMux I__10199 (
            .O(N__45686),
            .I(N__45683));
    LocalMux I__10198 (
            .O(N__45683),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_3 ));
    InMux I__10197 (
            .O(N__45680),
            .I(N__45677));
    LocalMux I__10196 (
            .O(N__45677),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_6 ));
    InMux I__10195 (
            .O(N__45674),
            .I(N__45671));
    LocalMux I__10194 (
            .O(N__45671),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_6 ));
    InMux I__10193 (
            .O(N__45668),
            .I(N__45665));
    LocalMux I__10192 (
            .O(N__45665),
            .I(N__45662));
    Span4Mux_v I__10191 (
            .O(N__45662),
            .I(N__45659));
    Span4Mux_h I__10190 (
            .O(N__45659),
            .I(N__45656));
    Odrv4 I__10189 (
            .O(N__45656),
            .I(sDAC_mem_13Z0Z_0));
    InMux I__10188 (
            .O(N__45653),
            .I(N__45650));
    LocalMux I__10187 (
            .O(N__45650),
            .I(N__45647));
    Span4Mux_v I__10186 (
            .O(N__45647),
            .I(N__45644));
    Span4Mux_h I__10185 (
            .O(N__45644),
            .I(N__45641));
    Odrv4 I__10184 (
            .O(N__45641),
            .I(sDAC_mem_13Z0Z_1));
    InMux I__10183 (
            .O(N__45638),
            .I(N__45635));
    LocalMux I__10182 (
            .O(N__45635),
            .I(N__45632));
    Span4Mux_h I__10181 (
            .O(N__45632),
            .I(N__45629));
    Span4Mux_h I__10180 (
            .O(N__45629),
            .I(N__45626));
    Odrv4 I__10179 (
            .O(N__45626),
            .I(sDAC_mem_13Z0Z_2));
    InMux I__10178 (
            .O(N__45623),
            .I(N__45620));
    LocalMux I__10177 (
            .O(N__45620),
            .I(N__45617));
    Span12Mux_h I__10176 (
            .O(N__45617),
            .I(N__45614));
    Odrv12 I__10175 (
            .O(N__45614),
            .I(sDAC_mem_13Z0Z_3));
    InMux I__10174 (
            .O(N__45611),
            .I(N__45608));
    LocalMux I__10173 (
            .O(N__45608),
            .I(N__45597));
    InMux I__10172 (
            .O(N__45607),
            .I(N__45594));
    InMux I__10171 (
            .O(N__45606),
            .I(N__45589));
    InMux I__10170 (
            .O(N__45605),
            .I(N__45586));
    InMux I__10169 (
            .O(N__45604),
            .I(N__45582));
    InMux I__10168 (
            .O(N__45603),
            .I(N__45571));
    InMux I__10167 (
            .O(N__45602),
            .I(N__45564));
    InMux I__10166 (
            .O(N__45601),
            .I(N__45555));
    InMux I__10165 (
            .O(N__45600),
            .I(N__45551));
    Span4Mux_v I__10164 (
            .O(N__45597),
            .I(N__45546));
    LocalMux I__10163 (
            .O(N__45594),
            .I(N__45546));
    InMux I__10162 (
            .O(N__45593),
            .I(N__45543));
    InMux I__10161 (
            .O(N__45592),
            .I(N__45540));
    LocalMux I__10160 (
            .O(N__45589),
            .I(N__45535));
    LocalMux I__10159 (
            .O(N__45586),
            .I(N__45535));
    InMux I__10158 (
            .O(N__45585),
            .I(N__45532));
    LocalMux I__10157 (
            .O(N__45582),
            .I(N__45525));
    InMux I__10156 (
            .O(N__45581),
            .I(N__45522));
    InMux I__10155 (
            .O(N__45580),
            .I(N__45519));
    InMux I__10154 (
            .O(N__45579),
            .I(N__45516));
    InMux I__10153 (
            .O(N__45578),
            .I(N__45513));
    InMux I__10152 (
            .O(N__45577),
            .I(N__45510));
    InMux I__10151 (
            .O(N__45576),
            .I(N__45503));
    InMux I__10150 (
            .O(N__45575),
            .I(N__45500));
    InMux I__10149 (
            .O(N__45574),
            .I(N__45497));
    LocalMux I__10148 (
            .O(N__45571),
            .I(N__45494));
    InMux I__10147 (
            .O(N__45570),
            .I(N__45491));
    InMux I__10146 (
            .O(N__45569),
            .I(N__45488));
    InMux I__10145 (
            .O(N__45568),
            .I(N__45485));
    InMux I__10144 (
            .O(N__45567),
            .I(N__45482));
    LocalMux I__10143 (
            .O(N__45564),
            .I(N__45478));
    InMux I__10142 (
            .O(N__45563),
            .I(N__45475));
    InMux I__10141 (
            .O(N__45562),
            .I(N__45472));
    InMux I__10140 (
            .O(N__45561),
            .I(N__45469));
    InMux I__10139 (
            .O(N__45560),
            .I(N__45466));
    InMux I__10138 (
            .O(N__45559),
            .I(N__45463));
    InMux I__10137 (
            .O(N__45558),
            .I(N__45460));
    LocalMux I__10136 (
            .O(N__45555),
            .I(N__45457));
    InMux I__10135 (
            .O(N__45554),
            .I(N__45454));
    LocalMux I__10134 (
            .O(N__45551),
            .I(N__45451));
    Span4Mux_v I__10133 (
            .O(N__45546),
            .I(N__45444));
    LocalMux I__10132 (
            .O(N__45543),
            .I(N__45444));
    LocalMux I__10131 (
            .O(N__45540),
            .I(N__45444));
    Span4Mux_v I__10130 (
            .O(N__45535),
            .I(N__45439));
    LocalMux I__10129 (
            .O(N__45532),
            .I(N__45439));
    InMux I__10128 (
            .O(N__45531),
            .I(N__45436));
    InMux I__10127 (
            .O(N__45530),
            .I(N__45433));
    InMux I__10126 (
            .O(N__45529),
            .I(N__45430));
    InMux I__10125 (
            .O(N__45528),
            .I(N__45427));
    Span4Mux_v I__10124 (
            .O(N__45525),
            .I(N__45414));
    LocalMux I__10123 (
            .O(N__45522),
            .I(N__45414));
    LocalMux I__10122 (
            .O(N__45519),
            .I(N__45414));
    LocalMux I__10121 (
            .O(N__45516),
            .I(N__45414));
    LocalMux I__10120 (
            .O(N__45513),
            .I(N__45414));
    LocalMux I__10119 (
            .O(N__45510),
            .I(N__45414));
    InMux I__10118 (
            .O(N__45509),
            .I(N__45407));
    InMux I__10117 (
            .O(N__45508),
            .I(N__45404));
    InMux I__10116 (
            .O(N__45507),
            .I(N__45401));
    InMux I__10115 (
            .O(N__45506),
            .I(N__45398));
    LocalMux I__10114 (
            .O(N__45503),
            .I(N__45394));
    LocalMux I__10113 (
            .O(N__45500),
            .I(N__45389));
    LocalMux I__10112 (
            .O(N__45497),
            .I(N__45389));
    Span4Mux_v I__10111 (
            .O(N__45494),
            .I(N__45384));
    LocalMux I__10110 (
            .O(N__45491),
            .I(N__45375));
    LocalMux I__10109 (
            .O(N__45488),
            .I(N__45375));
    LocalMux I__10108 (
            .O(N__45485),
            .I(N__45375));
    LocalMux I__10107 (
            .O(N__45482),
            .I(N__45375));
    CascadeMux I__10106 (
            .O(N__45481),
            .I(N__45369));
    Span4Mux_v I__10105 (
            .O(N__45478),
            .I(N__45360));
    LocalMux I__10104 (
            .O(N__45475),
            .I(N__45360));
    LocalMux I__10103 (
            .O(N__45472),
            .I(N__45360));
    LocalMux I__10102 (
            .O(N__45469),
            .I(N__45360));
    LocalMux I__10101 (
            .O(N__45466),
            .I(N__45354));
    LocalMux I__10100 (
            .O(N__45463),
            .I(N__45354));
    LocalMux I__10099 (
            .O(N__45460),
            .I(N__45351));
    Span4Mux_v I__10098 (
            .O(N__45457),
            .I(N__45343));
    LocalMux I__10097 (
            .O(N__45454),
            .I(N__45343));
    Span4Mux_v I__10096 (
            .O(N__45451),
            .I(N__45338));
    Span4Mux_v I__10095 (
            .O(N__45444),
            .I(N__45338));
    Span4Mux_v I__10094 (
            .O(N__45439),
            .I(N__45333));
    LocalMux I__10093 (
            .O(N__45436),
            .I(N__45333));
    LocalMux I__10092 (
            .O(N__45433),
            .I(N__45326));
    LocalMux I__10091 (
            .O(N__45430),
            .I(N__45326));
    LocalMux I__10090 (
            .O(N__45427),
            .I(N__45326));
    Span4Mux_v I__10089 (
            .O(N__45414),
            .I(N__45323));
    InMux I__10088 (
            .O(N__45413),
            .I(N__45320));
    InMux I__10087 (
            .O(N__45412),
            .I(N__45317));
    InMux I__10086 (
            .O(N__45411),
            .I(N__45314));
    InMux I__10085 (
            .O(N__45410),
            .I(N__45311));
    LocalMux I__10084 (
            .O(N__45407),
            .I(N__45308));
    LocalMux I__10083 (
            .O(N__45404),
            .I(N__45301));
    LocalMux I__10082 (
            .O(N__45401),
            .I(N__45301));
    LocalMux I__10081 (
            .O(N__45398),
            .I(N__45301));
    InMux I__10080 (
            .O(N__45397),
            .I(N__45298));
    Span4Mux_v I__10079 (
            .O(N__45394),
            .I(N__45291));
    Span4Mux_v I__10078 (
            .O(N__45389),
            .I(N__45291));
    InMux I__10077 (
            .O(N__45388),
            .I(N__45288));
    InMux I__10076 (
            .O(N__45387),
            .I(N__45285));
    Span4Mux_h I__10075 (
            .O(N__45384),
            .I(N__45280));
    Span4Mux_v I__10074 (
            .O(N__45375),
            .I(N__45280));
    InMux I__10073 (
            .O(N__45374),
            .I(N__45277));
    InMux I__10072 (
            .O(N__45373),
            .I(N__45274));
    InMux I__10071 (
            .O(N__45372),
            .I(N__45271));
    InMux I__10070 (
            .O(N__45369),
            .I(N__45268));
    Sp12to4 I__10069 (
            .O(N__45360),
            .I(N__45265));
    InMux I__10068 (
            .O(N__45359),
            .I(N__45262));
    Span4Mux_v I__10067 (
            .O(N__45354),
            .I(N__45257));
    Span4Mux_v I__10066 (
            .O(N__45351),
            .I(N__45257));
    InMux I__10065 (
            .O(N__45350),
            .I(N__45254));
    InMux I__10064 (
            .O(N__45349),
            .I(N__45251));
    InMux I__10063 (
            .O(N__45348),
            .I(N__45248));
    Span4Mux_v I__10062 (
            .O(N__45343),
            .I(N__45245));
    Span4Mux_h I__10061 (
            .O(N__45338),
            .I(N__45238));
    Span4Mux_v I__10060 (
            .O(N__45333),
            .I(N__45238));
    Span4Mux_v I__10059 (
            .O(N__45326),
            .I(N__45238));
    Span4Mux_v I__10058 (
            .O(N__45323),
            .I(N__45227));
    LocalMux I__10057 (
            .O(N__45320),
            .I(N__45227));
    LocalMux I__10056 (
            .O(N__45317),
            .I(N__45227));
    LocalMux I__10055 (
            .O(N__45314),
            .I(N__45227));
    LocalMux I__10054 (
            .O(N__45311),
            .I(N__45227));
    Span4Mux_v I__10053 (
            .O(N__45308),
            .I(N__45221));
    Span4Mux_v I__10052 (
            .O(N__45301),
            .I(N__45218));
    LocalMux I__10051 (
            .O(N__45298),
            .I(N__45215));
    InMux I__10050 (
            .O(N__45297),
            .I(N__45212));
    InMux I__10049 (
            .O(N__45296),
            .I(N__45209));
    Span4Mux_v I__10048 (
            .O(N__45291),
            .I(N__45202));
    LocalMux I__10047 (
            .O(N__45288),
            .I(N__45202));
    LocalMux I__10046 (
            .O(N__45285),
            .I(N__45202));
    Span4Mux_v I__10045 (
            .O(N__45280),
            .I(N__45191));
    LocalMux I__10044 (
            .O(N__45277),
            .I(N__45191));
    LocalMux I__10043 (
            .O(N__45274),
            .I(N__45191));
    LocalMux I__10042 (
            .O(N__45271),
            .I(N__45191));
    LocalMux I__10041 (
            .O(N__45268),
            .I(N__45191));
    Span12Mux_v I__10040 (
            .O(N__45265),
            .I(N__45178));
    LocalMux I__10039 (
            .O(N__45262),
            .I(N__45178));
    Sp12to4 I__10038 (
            .O(N__45257),
            .I(N__45178));
    LocalMux I__10037 (
            .O(N__45254),
            .I(N__45178));
    LocalMux I__10036 (
            .O(N__45251),
            .I(N__45178));
    LocalMux I__10035 (
            .O(N__45248),
            .I(N__45178));
    Span4Mux_v I__10034 (
            .O(N__45245),
            .I(N__45171));
    Span4Mux_h I__10033 (
            .O(N__45238),
            .I(N__45171));
    Span4Mux_v I__10032 (
            .O(N__45227),
            .I(N__45171));
    InMux I__10031 (
            .O(N__45226),
            .I(N__45168));
    InMux I__10030 (
            .O(N__45225),
            .I(N__45165));
    InMux I__10029 (
            .O(N__45224),
            .I(N__45162));
    Span4Mux_h I__10028 (
            .O(N__45221),
            .I(N__45147));
    Span4Mux_h I__10027 (
            .O(N__45218),
            .I(N__45147));
    Span4Mux_v I__10026 (
            .O(N__45215),
            .I(N__45147));
    LocalMux I__10025 (
            .O(N__45212),
            .I(N__45147));
    LocalMux I__10024 (
            .O(N__45209),
            .I(N__45147));
    Span4Mux_v I__10023 (
            .O(N__45202),
            .I(N__45147));
    Span4Mux_v I__10022 (
            .O(N__45191),
            .I(N__45147));
    Odrv12 I__10021 (
            .O(N__45178),
            .I(spi_data_mosi_4));
    Odrv4 I__10020 (
            .O(N__45171),
            .I(spi_data_mosi_4));
    LocalMux I__10019 (
            .O(N__45168),
            .I(spi_data_mosi_4));
    LocalMux I__10018 (
            .O(N__45165),
            .I(spi_data_mosi_4));
    LocalMux I__10017 (
            .O(N__45162),
            .I(spi_data_mosi_4));
    Odrv4 I__10016 (
            .O(N__45147),
            .I(spi_data_mosi_4));
    InMux I__10015 (
            .O(N__45134),
            .I(N__45131));
    LocalMux I__10014 (
            .O(N__45131),
            .I(N__45128));
    Span4Mux_v I__10013 (
            .O(N__45128),
            .I(N__45125));
    Span4Mux_h I__10012 (
            .O(N__45125),
            .I(N__45122));
    Odrv4 I__10011 (
            .O(N__45122),
            .I(sDAC_mem_13Z0Z_4));
    InMux I__10010 (
            .O(N__45119),
            .I(N__45111));
    InMux I__10009 (
            .O(N__45118),
            .I(N__45108));
    InMux I__10008 (
            .O(N__45117),
            .I(N__45097));
    InMux I__10007 (
            .O(N__45116),
            .I(N__45091));
    InMux I__10006 (
            .O(N__45115),
            .I(N__45086));
    InMux I__10005 (
            .O(N__45114),
            .I(N__45082));
    LocalMux I__10004 (
            .O(N__45111),
            .I(N__45072));
    LocalMux I__10003 (
            .O(N__45108),
            .I(N__45072));
    InMux I__10002 (
            .O(N__45107),
            .I(N__45069));
    InMux I__10001 (
            .O(N__45106),
            .I(N__45061));
    InMux I__10000 (
            .O(N__45105),
            .I(N__45058));
    InMux I__9999 (
            .O(N__45104),
            .I(N__45050));
    InMux I__9998 (
            .O(N__45103),
            .I(N__45047));
    InMux I__9997 (
            .O(N__45102),
            .I(N__45044));
    InMux I__9996 (
            .O(N__45101),
            .I(N__45041));
    InMux I__9995 (
            .O(N__45100),
            .I(N__45038));
    LocalMux I__9994 (
            .O(N__45097),
            .I(N__45034));
    InMux I__9993 (
            .O(N__45096),
            .I(N__45031));
    InMux I__9992 (
            .O(N__45095),
            .I(N__45028));
    InMux I__9991 (
            .O(N__45094),
            .I(N__45025));
    LocalMux I__9990 (
            .O(N__45091),
            .I(N__45022));
    InMux I__9989 (
            .O(N__45090),
            .I(N__45019));
    InMux I__9988 (
            .O(N__45089),
            .I(N__45016));
    LocalMux I__9987 (
            .O(N__45086),
            .I(N__45013));
    InMux I__9986 (
            .O(N__45085),
            .I(N__45010));
    LocalMux I__9985 (
            .O(N__45082),
            .I(N__45006));
    InMux I__9984 (
            .O(N__45081),
            .I(N__45002));
    InMux I__9983 (
            .O(N__45080),
            .I(N__44997));
    InMux I__9982 (
            .O(N__45079),
            .I(N__44994));
    InMux I__9981 (
            .O(N__45078),
            .I(N__44991));
    InMux I__9980 (
            .O(N__45077),
            .I(N__44988));
    Span4Mux_h I__9979 (
            .O(N__45072),
            .I(N__44983));
    LocalMux I__9978 (
            .O(N__45069),
            .I(N__44983));
    InMux I__9977 (
            .O(N__45068),
            .I(N__44977));
    InMux I__9976 (
            .O(N__45067),
            .I(N__44974));
    InMux I__9975 (
            .O(N__45066),
            .I(N__44971));
    InMux I__9974 (
            .O(N__45065),
            .I(N__44968));
    InMux I__9973 (
            .O(N__45064),
            .I(N__44965));
    LocalMux I__9972 (
            .O(N__45061),
            .I(N__44962));
    LocalMux I__9971 (
            .O(N__45058),
            .I(N__44959));
    InMux I__9970 (
            .O(N__45057),
            .I(N__44956));
    InMux I__9969 (
            .O(N__45056),
            .I(N__44953));
    InMux I__9968 (
            .O(N__45055),
            .I(N__44948));
    InMux I__9967 (
            .O(N__45054),
            .I(N__44945));
    InMux I__9966 (
            .O(N__45053),
            .I(N__44942));
    LocalMux I__9965 (
            .O(N__45050),
            .I(N__44939));
    LocalMux I__9964 (
            .O(N__45047),
            .I(N__44930));
    LocalMux I__9963 (
            .O(N__45044),
            .I(N__44930));
    LocalMux I__9962 (
            .O(N__45041),
            .I(N__44930));
    LocalMux I__9961 (
            .O(N__45038),
            .I(N__44930));
    InMux I__9960 (
            .O(N__45037),
            .I(N__44925));
    Span4Mux_v I__9959 (
            .O(N__45034),
            .I(N__44920));
    LocalMux I__9958 (
            .O(N__45031),
            .I(N__44915));
    LocalMux I__9957 (
            .O(N__45028),
            .I(N__44915));
    LocalMux I__9956 (
            .O(N__45025),
            .I(N__44908));
    Span4Mux_v I__9955 (
            .O(N__45022),
            .I(N__44908));
    LocalMux I__9954 (
            .O(N__45019),
            .I(N__44908));
    LocalMux I__9953 (
            .O(N__45016),
            .I(N__44905));
    Span4Mux_h I__9952 (
            .O(N__45013),
            .I(N__44902));
    LocalMux I__9951 (
            .O(N__45010),
            .I(N__44899));
    InMux I__9950 (
            .O(N__45009),
            .I(N__44896));
    Span4Mux_h I__9949 (
            .O(N__45006),
            .I(N__44893));
    InMux I__9948 (
            .O(N__45005),
            .I(N__44890));
    LocalMux I__9947 (
            .O(N__45002),
            .I(N__44887));
    InMux I__9946 (
            .O(N__45001),
            .I(N__44884));
    InMux I__9945 (
            .O(N__45000),
            .I(N__44881));
    LocalMux I__9944 (
            .O(N__44997),
            .I(N__44876));
    LocalMux I__9943 (
            .O(N__44994),
            .I(N__44876));
    LocalMux I__9942 (
            .O(N__44991),
            .I(N__44871));
    LocalMux I__9941 (
            .O(N__44988),
            .I(N__44871));
    Span4Mux_v I__9940 (
            .O(N__44983),
            .I(N__44868));
    InMux I__9939 (
            .O(N__44982),
            .I(N__44864));
    InMux I__9938 (
            .O(N__44981),
            .I(N__44861));
    InMux I__9937 (
            .O(N__44980),
            .I(N__44858));
    LocalMux I__9936 (
            .O(N__44977),
            .I(N__44853));
    LocalMux I__9935 (
            .O(N__44974),
            .I(N__44853));
    LocalMux I__9934 (
            .O(N__44971),
            .I(N__44842));
    LocalMux I__9933 (
            .O(N__44968),
            .I(N__44842));
    LocalMux I__9932 (
            .O(N__44965),
            .I(N__44842));
    Span4Mux_h I__9931 (
            .O(N__44962),
            .I(N__44842));
    Span4Mux_v I__9930 (
            .O(N__44959),
            .I(N__44842));
    LocalMux I__9929 (
            .O(N__44956),
            .I(N__44835));
    LocalMux I__9928 (
            .O(N__44953),
            .I(N__44835));
    InMux I__9927 (
            .O(N__44952),
            .I(N__44830));
    InMux I__9926 (
            .O(N__44951),
            .I(N__44827));
    LocalMux I__9925 (
            .O(N__44948),
            .I(N__44820));
    LocalMux I__9924 (
            .O(N__44945),
            .I(N__44820));
    LocalMux I__9923 (
            .O(N__44942),
            .I(N__44820));
    Span4Mux_v I__9922 (
            .O(N__44939),
            .I(N__44815));
    Span4Mux_v I__9921 (
            .O(N__44930),
            .I(N__44815));
    InMux I__9920 (
            .O(N__44929),
            .I(N__44812));
    InMux I__9919 (
            .O(N__44928),
            .I(N__44809));
    LocalMux I__9918 (
            .O(N__44925),
            .I(N__44806));
    InMux I__9917 (
            .O(N__44924),
            .I(N__44803));
    InMux I__9916 (
            .O(N__44923),
            .I(N__44800));
    Span4Mux_h I__9915 (
            .O(N__44920),
            .I(N__44793));
    Span4Mux_v I__9914 (
            .O(N__44915),
            .I(N__44793));
    Span4Mux_v I__9913 (
            .O(N__44908),
            .I(N__44793));
    Span4Mux_v I__9912 (
            .O(N__44905),
            .I(N__44788));
    Span4Mux_h I__9911 (
            .O(N__44902),
            .I(N__44788));
    Span4Mux_v I__9910 (
            .O(N__44899),
            .I(N__44781));
    LocalMux I__9909 (
            .O(N__44896),
            .I(N__44781));
    Span4Mux_h I__9908 (
            .O(N__44893),
            .I(N__44781));
    LocalMux I__9907 (
            .O(N__44890),
            .I(N__44774));
    Span4Mux_h I__9906 (
            .O(N__44887),
            .I(N__44774));
    LocalMux I__9905 (
            .O(N__44884),
            .I(N__44774));
    LocalMux I__9904 (
            .O(N__44881),
            .I(N__44771));
    Span4Mux_v I__9903 (
            .O(N__44876),
            .I(N__44764));
    Span4Mux_v I__9902 (
            .O(N__44871),
            .I(N__44764));
    Span4Mux_h I__9901 (
            .O(N__44868),
            .I(N__44764));
    InMux I__9900 (
            .O(N__44867),
            .I(N__44760));
    LocalMux I__9899 (
            .O(N__44864),
            .I(N__44753));
    LocalMux I__9898 (
            .O(N__44861),
            .I(N__44753));
    LocalMux I__9897 (
            .O(N__44858),
            .I(N__44753));
    Span4Mux_v I__9896 (
            .O(N__44853),
            .I(N__44748));
    Span4Mux_v I__9895 (
            .O(N__44842),
            .I(N__44748));
    InMux I__9894 (
            .O(N__44841),
            .I(N__44745));
    InMux I__9893 (
            .O(N__44840),
            .I(N__44742));
    Span4Mux_v I__9892 (
            .O(N__44835),
            .I(N__44739));
    InMux I__9891 (
            .O(N__44834),
            .I(N__44734));
    InMux I__9890 (
            .O(N__44833),
            .I(N__44734));
    LocalMux I__9889 (
            .O(N__44830),
            .I(N__44727));
    LocalMux I__9888 (
            .O(N__44827),
            .I(N__44720));
    Span4Mux_v I__9887 (
            .O(N__44820),
            .I(N__44720));
    Span4Mux_h I__9886 (
            .O(N__44815),
            .I(N__44720));
    LocalMux I__9885 (
            .O(N__44812),
            .I(N__44707));
    LocalMux I__9884 (
            .O(N__44809),
            .I(N__44707));
    Span4Mux_h I__9883 (
            .O(N__44806),
            .I(N__44707));
    LocalMux I__9882 (
            .O(N__44803),
            .I(N__44707));
    LocalMux I__9881 (
            .O(N__44800),
            .I(N__44707));
    Span4Mux_v I__9880 (
            .O(N__44793),
            .I(N__44707));
    Span4Mux_h I__9879 (
            .O(N__44788),
            .I(N__44702));
    Span4Mux_v I__9878 (
            .O(N__44781),
            .I(N__44702));
    Span4Mux_v I__9877 (
            .O(N__44774),
            .I(N__44699));
    Span4Mux_h I__9876 (
            .O(N__44771),
            .I(N__44694));
    Span4Mux_h I__9875 (
            .O(N__44764),
            .I(N__44694));
    InMux I__9874 (
            .O(N__44763),
            .I(N__44691));
    LocalMux I__9873 (
            .O(N__44760),
            .I(N__44684));
    Span4Mux_v I__9872 (
            .O(N__44753),
            .I(N__44684));
    Span4Mux_h I__9871 (
            .O(N__44748),
            .I(N__44684));
    LocalMux I__9870 (
            .O(N__44745),
            .I(N__44675));
    LocalMux I__9869 (
            .O(N__44742),
            .I(N__44675));
    Span4Mux_v I__9868 (
            .O(N__44739),
            .I(N__44675));
    LocalMux I__9867 (
            .O(N__44734),
            .I(N__44675));
    InMux I__9866 (
            .O(N__44733),
            .I(N__44672));
    InMux I__9865 (
            .O(N__44732),
            .I(N__44669));
    InMux I__9864 (
            .O(N__44731),
            .I(N__44666));
    InMux I__9863 (
            .O(N__44730),
            .I(N__44663));
    Span4Mux_v I__9862 (
            .O(N__44727),
            .I(N__44656));
    Span4Mux_h I__9861 (
            .O(N__44720),
            .I(N__44656));
    Span4Mux_v I__9860 (
            .O(N__44707),
            .I(N__44656));
    Span4Mux_v I__9859 (
            .O(N__44702),
            .I(N__44653));
    Span4Mux_h I__9858 (
            .O(N__44699),
            .I(N__44648));
    Span4Mux_v I__9857 (
            .O(N__44694),
            .I(N__44648));
    LocalMux I__9856 (
            .O(N__44691),
            .I(N__44641));
    Span4Mux_h I__9855 (
            .O(N__44684),
            .I(N__44641));
    Span4Mux_v I__9854 (
            .O(N__44675),
            .I(N__44641));
    LocalMux I__9853 (
            .O(N__44672),
            .I(spi_data_mosi_5));
    LocalMux I__9852 (
            .O(N__44669),
            .I(spi_data_mosi_5));
    LocalMux I__9851 (
            .O(N__44666),
            .I(spi_data_mosi_5));
    LocalMux I__9850 (
            .O(N__44663),
            .I(spi_data_mosi_5));
    Odrv4 I__9849 (
            .O(N__44656),
            .I(spi_data_mosi_5));
    Odrv4 I__9848 (
            .O(N__44653),
            .I(spi_data_mosi_5));
    Odrv4 I__9847 (
            .O(N__44648),
            .I(spi_data_mosi_5));
    Odrv4 I__9846 (
            .O(N__44641),
            .I(spi_data_mosi_5));
    InMux I__9845 (
            .O(N__44624),
            .I(N__44621));
    LocalMux I__9844 (
            .O(N__44621),
            .I(N__44618));
    Span4Mux_v I__9843 (
            .O(N__44618),
            .I(N__44615));
    Span4Mux_h I__9842 (
            .O(N__44615),
            .I(N__44612));
    Odrv4 I__9841 (
            .O(N__44612),
            .I(sDAC_mem_13Z0Z_5));
    InMux I__9840 (
            .O(N__44609),
            .I(N__44606));
    LocalMux I__9839 (
            .O(N__44606),
            .I(N__44603));
    Span4Mux_h I__9838 (
            .O(N__44603),
            .I(N__44600));
    Odrv4 I__9837 (
            .O(N__44600),
            .I(sDAC_mem_13Z0Z_6));
    InMux I__9836 (
            .O(N__44597),
            .I(N__44594));
    LocalMux I__9835 (
            .O(N__44594),
            .I(N__44591));
    Span4Mux_v I__9834 (
            .O(N__44591),
            .I(N__44588));
    Odrv4 I__9833 (
            .O(N__44588),
            .I(sDAC_mem_13Z0Z_7));
    CEMux I__9832 (
            .O(N__44585),
            .I(N__44582));
    LocalMux I__9831 (
            .O(N__44582),
            .I(N__44579));
    Span4Mux_h I__9830 (
            .O(N__44579),
            .I(N__44576));
    Span4Mux_h I__9829 (
            .O(N__44576),
            .I(N__44573));
    Odrv4 I__9828 (
            .O(N__44573),
            .I(sDAC_mem_13_1_sqmuxa));
    InMux I__9827 (
            .O(N__44570),
            .I(N__44567));
    LocalMux I__9826 (
            .O(N__44567),
            .I(N__44564));
    Span4Mux_v I__9825 (
            .O(N__44564),
            .I(N__44561));
    Span4Mux_h I__9824 (
            .O(N__44561),
            .I(N__44558));
    Span4Mux_v I__9823 (
            .O(N__44558),
            .I(N__44554));
    InMux I__9822 (
            .O(N__44557),
            .I(N__44551));
    Span4Mux_h I__9821 (
            .O(N__44554),
            .I(N__44548));
    LocalMux I__9820 (
            .O(N__44551),
            .I(\spi_slave_inst.tx_ready_iZ0 ));
    Odrv4 I__9819 (
            .O(N__44548),
            .I(\spi_slave_inst.tx_ready_iZ0 ));
    InMux I__9818 (
            .O(N__44543),
            .I(N__44540));
    LocalMux I__9817 (
            .O(N__44540),
            .I(N__44537));
    Span4Mux_v I__9816 (
            .O(N__44537),
            .I(N__44534));
    Odrv4 I__9815 (
            .O(N__44534),
            .I(sDAC_mem_33Z0Z_7));
    CEMux I__9814 (
            .O(N__44531),
            .I(N__44528));
    LocalMux I__9813 (
            .O(N__44528),
            .I(N__44525));
    Odrv4 I__9812 (
            .O(N__44525),
            .I(sDAC_mem_33_1_sqmuxa));
    InMux I__9811 (
            .O(N__44522),
            .I(N__44519));
    LocalMux I__9810 (
            .O(N__44519),
            .I(N__44516));
    Odrv4 I__9809 (
            .O(N__44516),
            .I(sDAC_mem_5Z0Z_0));
    InMux I__9808 (
            .O(N__44513),
            .I(N__44510));
    LocalMux I__9807 (
            .O(N__44510),
            .I(N__44507));
    Odrv4 I__9806 (
            .O(N__44507),
            .I(sDAC_mem_5Z0Z_1));
    InMux I__9805 (
            .O(N__44504),
            .I(N__44501));
    LocalMux I__9804 (
            .O(N__44501),
            .I(N__44498));
    Odrv4 I__9803 (
            .O(N__44498),
            .I(sDAC_mem_5Z0Z_2));
    InMux I__9802 (
            .O(N__44495),
            .I(N__44492));
    LocalMux I__9801 (
            .O(N__44492),
            .I(N__44489));
    Span4Mux_h I__9800 (
            .O(N__44489),
            .I(N__44486));
    Odrv4 I__9799 (
            .O(N__44486),
            .I(sDAC_mem_5Z0Z_3));
    InMux I__9798 (
            .O(N__44483),
            .I(N__44480));
    LocalMux I__9797 (
            .O(N__44480),
            .I(N__44477));
    Span4Mux_h I__9796 (
            .O(N__44477),
            .I(N__44474));
    Odrv4 I__9795 (
            .O(N__44474),
            .I(sDAC_mem_5Z0Z_4));
    InMux I__9794 (
            .O(N__44471),
            .I(N__44468));
    LocalMux I__9793 (
            .O(N__44468),
            .I(N__44465));
    Span4Mux_h I__9792 (
            .O(N__44465),
            .I(N__44462));
    Odrv4 I__9791 (
            .O(N__44462),
            .I(sDAC_mem_5Z0Z_5));
    InMux I__9790 (
            .O(N__44459),
            .I(N__44456));
    LocalMux I__9789 (
            .O(N__44456),
            .I(N__44453));
    Span4Mux_v I__9788 (
            .O(N__44453),
            .I(N__44450));
    Odrv4 I__9787 (
            .O(N__44450),
            .I(sDAC_mem_5Z0Z_6));
    InMux I__9786 (
            .O(N__44447),
            .I(N__44444));
    LocalMux I__9785 (
            .O(N__44444),
            .I(N__44441));
    Span4Mux_h I__9784 (
            .O(N__44441),
            .I(N__44438));
    Odrv4 I__9783 (
            .O(N__44438),
            .I(sDAC_mem_5Z0Z_7));
    CEMux I__9782 (
            .O(N__44435),
            .I(N__44432));
    LocalMux I__9781 (
            .O(N__44432),
            .I(N__44429));
    Span12Mux_s10_h I__9780 (
            .O(N__44429),
            .I(N__44426));
    Odrv12 I__9779 (
            .O(N__44426),
            .I(sDAC_mem_5_1_sqmuxa));
    InMux I__9778 (
            .O(N__44423),
            .I(N__44420));
    LocalMux I__9777 (
            .O(N__44420),
            .I(N__44417));
    Odrv4 I__9776 (
            .O(N__44417),
            .I(sDAC_mem_1Z0Z_6));
    InMux I__9775 (
            .O(N__44414),
            .I(N__44411));
    LocalMux I__9774 (
            .O(N__44411),
            .I(N__44408));
    Span12Mux_v I__9773 (
            .O(N__44408),
            .I(N__44405));
    Odrv12 I__9772 (
            .O(N__44405),
            .I(sDAC_mem_1Z0Z_7));
    CEMux I__9771 (
            .O(N__44402),
            .I(N__44399));
    LocalMux I__9770 (
            .O(N__44399),
            .I(N__44396));
    Span4Mux_v I__9769 (
            .O(N__44396),
            .I(N__44393));
    Odrv4 I__9768 (
            .O(N__44393),
            .I(sDAC_mem_1_1_sqmuxa));
    InMux I__9767 (
            .O(N__44390),
            .I(N__44387));
    LocalMux I__9766 (
            .O(N__44387),
            .I(N__44384));
    Span4Mux_h I__9765 (
            .O(N__44384),
            .I(N__44381));
    Odrv4 I__9764 (
            .O(N__44381),
            .I(sDAC_mem_33Z0Z_0));
    InMux I__9763 (
            .O(N__44378),
            .I(N__44375));
    LocalMux I__9762 (
            .O(N__44375),
            .I(N__44372));
    Odrv4 I__9761 (
            .O(N__44372),
            .I(sDAC_mem_33Z0Z_1));
    InMux I__9760 (
            .O(N__44369),
            .I(N__44366));
    LocalMux I__9759 (
            .O(N__44366),
            .I(N__44363));
    Odrv4 I__9758 (
            .O(N__44363),
            .I(sDAC_mem_33Z0Z_2));
    InMux I__9757 (
            .O(N__44360),
            .I(N__44357));
    LocalMux I__9756 (
            .O(N__44357),
            .I(N__44354));
    Span4Mux_h I__9755 (
            .O(N__44354),
            .I(N__44351));
    Odrv4 I__9754 (
            .O(N__44351),
            .I(sDAC_mem_33Z0Z_3));
    InMux I__9753 (
            .O(N__44348),
            .I(N__44345));
    LocalMux I__9752 (
            .O(N__44345),
            .I(N__44342));
    Span4Mux_h I__9751 (
            .O(N__44342),
            .I(N__44339));
    Odrv4 I__9750 (
            .O(N__44339),
            .I(sDAC_mem_33Z0Z_4));
    InMux I__9749 (
            .O(N__44336),
            .I(N__44333));
    LocalMux I__9748 (
            .O(N__44333),
            .I(N__44330));
    Span4Mux_h I__9747 (
            .O(N__44330),
            .I(N__44327));
    Odrv4 I__9746 (
            .O(N__44327),
            .I(sDAC_mem_33Z0Z_5));
    InMux I__9745 (
            .O(N__44324),
            .I(N__44321));
    LocalMux I__9744 (
            .O(N__44321),
            .I(N__44318));
    Span4Mux_h I__9743 (
            .O(N__44318),
            .I(N__44315));
    Odrv4 I__9742 (
            .O(N__44315),
            .I(sDAC_mem_33Z0Z_6));
    InMux I__9741 (
            .O(N__44312),
            .I(N__44309));
    LocalMux I__9740 (
            .O(N__44309),
            .I(N__44306));
    Span4Mux_h I__9739 (
            .O(N__44306),
            .I(N__44303));
    Span4Mux_h I__9738 (
            .O(N__44303),
            .I(N__44300));
    Odrv4 I__9737 (
            .O(N__44300),
            .I(sDAC_mem_7Z0Z_4));
    InMux I__9736 (
            .O(N__44297),
            .I(N__44294));
    LocalMux I__9735 (
            .O(N__44294),
            .I(N__44291));
    Span4Mux_v I__9734 (
            .O(N__44291),
            .I(N__44288));
    Odrv4 I__9733 (
            .O(N__44288),
            .I(sDAC_mem_7Z0Z_6));
    CEMux I__9732 (
            .O(N__44285),
            .I(N__44282));
    LocalMux I__9731 (
            .O(N__44282),
            .I(N__44279));
    Span4Mux_h I__9730 (
            .O(N__44279),
            .I(N__44275));
    CEMux I__9729 (
            .O(N__44278),
            .I(N__44272));
    Span4Mux_h I__9728 (
            .O(N__44275),
            .I(N__44267));
    LocalMux I__9727 (
            .O(N__44272),
            .I(N__44267));
    Span4Mux_v I__9726 (
            .O(N__44267),
            .I(N__44264));
    Odrv4 I__9725 (
            .O(N__44264),
            .I(sDAC_mem_7_1_sqmuxa));
    InMux I__9724 (
            .O(N__44261),
            .I(N__44258));
    LocalMux I__9723 (
            .O(N__44258),
            .I(N__44255));
    Span4Mux_h I__9722 (
            .O(N__44255),
            .I(N__44252));
    Span4Mux_v I__9721 (
            .O(N__44252),
            .I(N__44249));
    Odrv4 I__9720 (
            .O(N__44249),
            .I(sDAC_mem_3Z0Z_7));
    CEMux I__9719 (
            .O(N__44246),
            .I(N__44240));
    CEMux I__9718 (
            .O(N__44245),
            .I(N__44234));
    CEMux I__9717 (
            .O(N__44244),
            .I(N__44231));
    CEMux I__9716 (
            .O(N__44243),
            .I(N__44228));
    LocalMux I__9715 (
            .O(N__44240),
            .I(N__44225));
    CEMux I__9714 (
            .O(N__44239),
            .I(N__44221));
    CEMux I__9713 (
            .O(N__44238),
            .I(N__44218));
    CEMux I__9712 (
            .O(N__44237),
            .I(N__44215));
    LocalMux I__9711 (
            .O(N__44234),
            .I(N__44212));
    LocalMux I__9710 (
            .O(N__44231),
            .I(N__44209));
    LocalMux I__9709 (
            .O(N__44228),
            .I(N__44206));
    Span4Mux_h I__9708 (
            .O(N__44225),
            .I(N__44203));
    CEMux I__9707 (
            .O(N__44224),
            .I(N__44200));
    LocalMux I__9706 (
            .O(N__44221),
            .I(N__44197));
    LocalMux I__9705 (
            .O(N__44218),
            .I(N__44194));
    LocalMux I__9704 (
            .O(N__44215),
            .I(N__44191));
    Span4Mux_v I__9703 (
            .O(N__44212),
            .I(N__44184));
    Span4Mux_v I__9702 (
            .O(N__44209),
            .I(N__44184));
    Span4Mux_v I__9701 (
            .O(N__44206),
            .I(N__44184));
    Span4Mux_h I__9700 (
            .O(N__44203),
            .I(N__44181));
    LocalMux I__9699 (
            .O(N__44200),
            .I(N__44178));
    Span4Mux_v I__9698 (
            .O(N__44197),
            .I(N__44175));
    Span4Mux_v I__9697 (
            .O(N__44194),
            .I(N__44170));
    Span4Mux_h I__9696 (
            .O(N__44191),
            .I(N__44170));
    Span4Mux_h I__9695 (
            .O(N__44184),
            .I(N__44167));
    Span4Mux_h I__9694 (
            .O(N__44181),
            .I(N__44164));
    Span4Mux_v I__9693 (
            .O(N__44178),
            .I(N__44161));
    Sp12to4 I__9692 (
            .O(N__44175),
            .I(N__44158));
    Span4Mux_h I__9691 (
            .O(N__44170),
            .I(N__44155));
    Span4Mux_h I__9690 (
            .O(N__44167),
            .I(N__44152));
    Span4Mux_h I__9689 (
            .O(N__44164),
            .I(N__44149));
    Sp12to4 I__9688 (
            .O(N__44161),
            .I(N__44144));
    Span12Mux_h I__9687 (
            .O(N__44158),
            .I(N__44144));
    Odrv4 I__9686 (
            .O(N__44155),
            .I(sDAC_mem_3_1_sqmuxa));
    Odrv4 I__9685 (
            .O(N__44152),
            .I(sDAC_mem_3_1_sqmuxa));
    Odrv4 I__9684 (
            .O(N__44149),
            .I(sDAC_mem_3_1_sqmuxa));
    Odrv12 I__9683 (
            .O(N__44144),
            .I(sDAC_mem_3_1_sqmuxa));
    InMux I__9682 (
            .O(N__44135),
            .I(N__44132));
    LocalMux I__9681 (
            .O(N__44132),
            .I(N__44129));
    Span4Mux_h I__9680 (
            .O(N__44129),
            .I(N__44126));
    Odrv4 I__9679 (
            .O(N__44126),
            .I(sDAC_mem_1Z0Z_0));
    InMux I__9678 (
            .O(N__44123),
            .I(N__44120));
    LocalMux I__9677 (
            .O(N__44120),
            .I(N__44117));
    Span4Mux_v I__9676 (
            .O(N__44117),
            .I(N__44114));
    Odrv4 I__9675 (
            .O(N__44114),
            .I(sDAC_mem_1Z0Z_1));
    InMux I__9674 (
            .O(N__44111),
            .I(N__44108));
    LocalMux I__9673 (
            .O(N__44108),
            .I(N__44105));
    Odrv4 I__9672 (
            .O(N__44105),
            .I(sDAC_mem_1Z0Z_2));
    InMux I__9671 (
            .O(N__44102),
            .I(N__44099));
    LocalMux I__9670 (
            .O(N__44099),
            .I(N__44096));
    Odrv4 I__9669 (
            .O(N__44096),
            .I(sDAC_mem_1Z0Z_3));
    InMux I__9668 (
            .O(N__44093),
            .I(N__44090));
    LocalMux I__9667 (
            .O(N__44090),
            .I(N__44087));
    Odrv4 I__9666 (
            .O(N__44087),
            .I(sDAC_mem_1Z0Z_4));
    InMux I__9665 (
            .O(N__44084),
            .I(N__44081));
    LocalMux I__9664 (
            .O(N__44081),
            .I(N__44078));
    Odrv4 I__9663 (
            .O(N__44078),
            .I(sDAC_mem_1Z0Z_5));
    IoInMux I__9662 (
            .O(N__44075),
            .I(N__44072));
    LocalMux I__9661 (
            .O(N__44072),
            .I(N__44069));
    IoSpan4Mux I__9660 (
            .O(N__44069),
            .I(N__44066));
    Span4Mux_s3_h I__9659 (
            .O(N__44066),
            .I(N__44063));
    Span4Mux_v I__9658 (
            .O(N__44063),
            .I(N__44060));
    Span4Mux_v I__9657 (
            .O(N__44060),
            .I(N__44057));
    Sp12to4 I__9656 (
            .O(N__44057),
            .I(N__44053));
    InMux I__9655 (
            .O(N__44056),
            .I(N__44050));
    Odrv12 I__9654 (
            .O(N__44053),
            .I(RAM_DATA_cl_10Z0Z_15));
    LocalMux I__9653 (
            .O(N__44050),
            .I(RAM_DATA_cl_10Z0Z_15));
    IoInMux I__9652 (
            .O(N__44045),
            .I(N__44042));
    LocalMux I__9651 (
            .O(N__44042),
            .I(N__44039));
    Span4Mux_s0_v I__9650 (
            .O(N__44039),
            .I(N__44036));
    Span4Mux_v I__9649 (
            .O(N__44036),
            .I(N__44033));
    Span4Mux_v I__9648 (
            .O(N__44033),
            .I(N__44029));
    CascadeMux I__9647 (
            .O(N__44032),
            .I(N__44026));
    Sp12to4 I__9646 (
            .O(N__44029),
            .I(N__44023));
    InMux I__9645 (
            .O(N__44026),
            .I(N__44020));
    Odrv12 I__9644 (
            .O(N__44023),
            .I(RAM_DATA_cl_3Z0Z_15));
    LocalMux I__9643 (
            .O(N__44020),
            .I(RAM_DATA_cl_3Z0Z_15));
    IoInMux I__9642 (
            .O(N__44015),
            .I(N__44012));
    LocalMux I__9641 (
            .O(N__44012),
            .I(N__44009));
    IoSpan4Mux I__9640 (
            .O(N__44009),
            .I(N__44006));
    Span4Mux_s0_v I__9639 (
            .O(N__44006),
            .I(N__44003));
    Span4Mux_v I__9638 (
            .O(N__44003),
            .I(N__44000));
    Span4Mux_v I__9637 (
            .O(N__44000),
            .I(N__43996));
    InMux I__9636 (
            .O(N__43999),
            .I(N__43993));
    Odrv4 I__9635 (
            .O(N__43996),
            .I(RAM_DATA_cl_4Z0Z_15));
    LocalMux I__9634 (
            .O(N__43993),
            .I(RAM_DATA_cl_4Z0Z_15));
    IoInMux I__9633 (
            .O(N__43988),
            .I(N__43985));
    LocalMux I__9632 (
            .O(N__43985),
            .I(N__43982));
    Span4Mux_s3_h I__9631 (
            .O(N__43982),
            .I(N__43979));
    Span4Mux_v I__9630 (
            .O(N__43979),
            .I(N__43976));
    Span4Mux_v I__9629 (
            .O(N__43976),
            .I(N__43972));
    CascadeMux I__9628 (
            .O(N__43975),
            .I(N__43969));
    Span4Mux_h I__9627 (
            .O(N__43972),
            .I(N__43966));
    InMux I__9626 (
            .O(N__43969),
            .I(N__43963));
    Odrv4 I__9625 (
            .O(N__43966),
            .I(RAM_DATA_cl_2Z0Z_15));
    LocalMux I__9624 (
            .O(N__43963),
            .I(RAM_DATA_cl_2Z0Z_15));
    CEMux I__9623 (
            .O(N__43958),
            .I(N__43922));
    CEMux I__9622 (
            .O(N__43957),
            .I(N__43922));
    CEMux I__9621 (
            .O(N__43956),
            .I(N__43922));
    CEMux I__9620 (
            .O(N__43955),
            .I(N__43922));
    CEMux I__9619 (
            .O(N__43954),
            .I(N__43922));
    CEMux I__9618 (
            .O(N__43953),
            .I(N__43922));
    CEMux I__9617 (
            .O(N__43952),
            .I(N__43922));
    CEMux I__9616 (
            .O(N__43951),
            .I(N__43922));
    CEMux I__9615 (
            .O(N__43950),
            .I(N__43922));
    CEMux I__9614 (
            .O(N__43949),
            .I(N__43922));
    CEMux I__9613 (
            .O(N__43948),
            .I(N__43922));
    CEMux I__9612 (
            .O(N__43947),
            .I(N__43922));
    GlobalMux I__9611 (
            .O(N__43922),
            .I(N__43919));
    gio2CtrlBuf I__9610 (
            .O(N__43919),
            .I(op_eq_scounterdac10_g));
    InMux I__9609 (
            .O(N__43916),
            .I(N__43913));
    LocalMux I__9608 (
            .O(N__43913),
            .I(N__43910));
    Odrv4 I__9607 (
            .O(N__43910),
            .I(sDAC_dataZ0Z_2));
    CEMux I__9606 (
            .O(N__43907),
            .I(N__43904));
    LocalMux I__9605 (
            .O(N__43904),
            .I(N__43898));
    CEMux I__9604 (
            .O(N__43903),
            .I(N__43895));
    CEMux I__9603 (
            .O(N__43902),
            .I(N__43892));
    CEMux I__9602 (
            .O(N__43901),
            .I(N__43889));
    Span4Mux_h I__9601 (
            .O(N__43898),
            .I(N__43883));
    LocalMux I__9600 (
            .O(N__43895),
            .I(N__43883));
    LocalMux I__9599 (
            .O(N__43892),
            .I(N__43880));
    LocalMux I__9598 (
            .O(N__43889),
            .I(N__43877));
    CascadeMux I__9597 (
            .O(N__43888),
            .I(N__43874));
    Span4Mux_h I__9596 (
            .O(N__43883),
            .I(N__43871));
    Span4Mux_h I__9595 (
            .O(N__43880),
            .I(N__43868));
    Span4Mux_h I__9594 (
            .O(N__43877),
            .I(N__43865));
    InMux I__9593 (
            .O(N__43874),
            .I(N__43862));
    Odrv4 I__9592 (
            .O(N__43871),
            .I(\spi_master_inst.spi_data_path_u1.tx_ready_iZ0 ));
    Odrv4 I__9591 (
            .O(N__43868),
            .I(\spi_master_inst.spi_data_path_u1.tx_ready_iZ0 ));
    Odrv4 I__9590 (
            .O(N__43865),
            .I(\spi_master_inst.spi_data_path_u1.tx_ready_iZ0 ));
    LocalMux I__9589 (
            .O(N__43862),
            .I(\spi_master_inst.spi_data_path_u1.tx_ready_iZ0 ));
    InMux I__9588 (
            .O(N__43853),
            .I(N__43850));
    LocalMux I__9587 (
            .O(N__43850),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_2 ));
    InMux I__9586 (
            .O(N__43847),
            .I(N__43844));
    LocalMux I__9585 (
            .O(N__43844),
            .I(N__43841));
    Span12Mux_h I__9584 (
            .O(N__43841),
            .I(N__43838));
    Odrv12 I__9583 (
            .O(N__43838),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2 ));
    InMux I__9582 (
            .O(N__43835),
            .I(N__43832));
    LocalMux I__9581 (
            .O(N__43832),
            .I(N__43829));
    Span4Mux_h I__9580 (
            .O(N__43829),
            .I(N__43826));
    Span4Mux_h I__9579 (
            .O(N__43826),
            .I(N__43823));
    Odrv4 I__9578 (
            .O(N__43823),
            .I(sDAC_mem_7Z0Z_2));
    InMux I__9577 (
            .O(N__43820),
            .I(N__43817));
    LocalMux I__9576 (
            .O(N__43817),
            .I(N__43814));
    Span12Mux_v I__9575 (
            .O(N__43814),
            .I(N__43811));
    Odrv12 I__9574 (
            .O(N__43811),
            .I(sDAC_mem_7Z0Z_3));
    InMux I__9573 (
            .O(N__43808),
            .I(N__43805));
    LocalMux I__9572 (
            .O(N__43805),
            .I(N__43802));
    Span4Mux_h I__9571 (
            .O(N__43802),
            .I(N__43799));
    Span4Mux_v I__9570 (
            .O(N__43799),
            .I(N__43796));
    Span4Mux_v I__9569 (
            .O(N__43796),
            .I(N__43793));
    IoSpan4Mux I__9568 (
            .O(N__43793),
            .I(N__43790));
    Odrv4 I__9567 (
            .O(N__43790),
            .I(RAM_DATA_in_1));
    InMux I__9566 (
            .O(N__43787),
            .I(N__43784));
    LocalMux I__9565 (
            .O(N__43784),
            .I(N__43781));
    Span12Mux_h I__9564 (
            .O(N__43781),
            .I(N__43778));
    Span12Mux_v I__9563 (
            .O(N__43778),
            .I(N__43775));
    Odrv12 I__9562 (
            .O(N__43775),
            .I(RAM_DATA_in_9));
    CascadeMux I__9561 (
            .O(N__43772),
            .I(N__43762));
    CascadeMux I__9560 (
            .O(N__43771),
            .I(N__43759));
    CascadeMux I__9559 (
            .O(N__43770),
            .I(N__43756));
    InMux I__9558 (
            .O(N__43769),
            .I(N__43751));
    InMux I__9557 (
            .O(N__43768),
            .I(N__43751));
    InMux I__9556 (
            .O(N__43767),
            .I(N__43748));
    InMux I__9555 (
            .O(N__43766),
            .I(N__43737));
    InMux I__9554 (
            .O(N__43765),
            .I(N__43737));
    InMux I__9553 (
            .O(N__43762),
            .I(N__43737));
    InMux I__9552 (
            .O(N__43759),
            .I(N__43737));
    InMux I__9551 (
            .O(N__43756),
            .I(N__43737));
    LocalMux I__9550 (
            .O(N__43751),
            .I(N__43732));
    LocalMux I__9549 (
            .O(N__43748),
            .I(N__43729));
    LocalMux I__9548 (
            .O(N__43737),
            .I(N__43726));
    InMux I__9547 (
            .O(N__43736),
            .I(N__43723));
    InMux I__9546 (
            .O(N__43735),
            .I(N__43720));
    Span4Mux_h I__9545 (
            .O(N__43732),
            .I(N__43717));
    Span4Mux_h I__9544 (
            .O(N__43729),
            .I(N__43714));
    Span4Mux_v I__9543 (
            .O(N__43726),
            .I(N__43709));
    LocalMux I__9542 (
            .O(N__43723),
            .I(N__43709));
    LocalMux I__9541 (
            .O(N__43720),
            .I(N_75));
    Odrv4 I__9540 (
            .O(N__43717),
            .I(N_75));
    Odrv4 I__9539 (
            .O(N__43714),
            .I(N_75));
    Odrv4 I__9538 (
            .O(N__43709),
            .I(N_75));
    InMux I__9537 (
            .O(N__43700),
            .I(N__43697));
    LocalMux I__9536 (
            .O(N__43697),
            .I(N__43694));
    Odrv4 I__9535 (
            .O(N__43694),
            .I(spi_data_misoZ0Z_1));
    CEMux I__9534 (
            .O(N__43691),
            .I(N__43688));
    LocalMux I__9533 (
            .O(N__43688),
            .I(N__43683));
    CEMux I__9532 (
            .O(N__43687),
            .I(N__43680));
    CEMux I__9531 (
            .O(N__43686),
            .I(N__43677));
    Span4Mux_v I__9530 (
            .O(N__43683),
            .I(N__43674));
    LocalMux I__9529 (
            .O(N__43680),
            .I(N__43671));
    LocalMux I__9528 (
            .O(N__43677),
            .I(N__43668));
    Odrv4 I__9527 (
            .O(N__43674),
            .I(sSPI_MSB0LSB1_RNIGRPGZ0Z4));
    Odrv4 I__9526 (
            .O(N__43671),
            .I(sSPI_MSB0LSB1_RNIGRPGZ0Z4));
    Odrv12 I__9525 (
            .O(N__43668),
            .I(sSPI_MSB0LSB1_RNIGRPGZ0Z4));
    InMux I__9524 (
            .O(N__43661),
            .I(N__43658));
    LocalMux I__9523 (
            .O(N__43658),
            .I(N__43655));
    Span4Mux_v I__9522 (
            .O(N__43655),
            .I(N__43652));
    Span4Mux_h I__9521 (
            .O(N__43652),
            .I(N__43649));
    Sp12to4 I__9520 (
            .O(N__43649),
            .I(N__43646));
    Span12Mux_h I__9519 (
            .O(N__43646),
            .I(N__43642));
    InMux I__9518 (
            .O(N__43645),
            .I(N__43639));
    Odrv12 I__9517 (
            .O(N__43642),
            .I(sRAM_pointer_writeZ0Z_8));
    LocalMux I__9516 (
            .O(N__43639),
            .I(sRAM_pointer_writeZ0Z_8));
    CascadeMux I__9515 (
            .O(N__43634),
            .I(N__43631));
    InMux I__9514 (
            .O(N__43631),
            .I(N__43628));
    LocalMux I__9513 (
            .O(N__43628),
            .I(N__43625));
    Span4Mux_h I__9512 (
            .O(N__43625),
            .I(N__43622));
    Span4Mux_h I__9511 (
            .O(N__43622),
            .I(N__43618));
    InMux I__9510 (
            .O(N__43621),
            .I(N__43615));
    Odrv4 I__9509 (
            .O(N__43618),
            .I(sRAM_pointer_readZ0Z_8));
    LocalMux I__9508 (
            .O(N__43615),
            .I(sRAM_pointer_readZ0Z_8));
    IoInMux I__9507 (
            .O(N__43610),
            .I(N__43607));
    LocalMux I__9506 (
            .O(N__43607),
            .I(N__43604));
    IoSpan4Mux I__9505 (
            .O(N__43604),
            .I(N__43601));
    Span4Mux_s3_h I__9504 (
            .O(N__43601),
            .I(N__43598));
    Span4Mux_h I__9503 (
            .O(N__43598),
            .I(N__43595));
    Span4Mux_v I__9502 (
            .O(N__43595),
            .I(N__43592));
    Odrv4 I__9501 (
            .O(N__43592),
            .I(RAM_ADD_c_8));
    InMux I__9500 (
            .O(N__43589),
            .I(N__43586));
    LocalMux I__9499 (
            .O(N__43586),
            .I(N__43583));
    Span4Mux_h I__9498 (
            .O(N__43583),
            .I(N__43580));
    Span4Mux_h I__9497 (
            .O(N__43580),
            .I(N__43577));
    Sp12to4 I__9496 (
            .O(N__43577),
            .I(N__43574));
    Span12Mux_v I__9495 (
            .O(N__43574),
            .I(N__43570));
    InMux I__9494 (
            .O(N__43573),
            .I(N__43567));
    Odrv12 I__9493 (
            .O(N__43570),
            .I(sRAM_pointer_writeZ0Z_4));
    LocalMux I__9492 (
            .O(N__43567),
            .I(sRAM_pointer_writeZ0Z_4));
    CascadeMux I__9491 (
            .O(N__43562),
            .I(N__43559));
    InMux I__9490 (
            .O(N__43559),
            .I(N__43556));
    LocalMux I__9489 (
            .O(N__43556),
            .I(N__43553));
    Span4Mux_h I__9488 (
            .O(N__43553),
            .I(N__43550));
    Span4Mux_h I__9487 (
            .O(N__43550),
            .I(N__43546));
    InMux I__9486 (
            .O(N__43549),
            .I(N__43543));
    Odrv4 I__9485 (
            .O(N__43546),
            .I(sRAM_pointer_readZ0Z_4));
    LocalMux I__9484 (
            .O(N__43543),
            .I(sRAM_pointer_readZ0Z_4));
    IoInMux I__9483 (
            .O(N__43538),
            .I(N__43535));
    LocalMux I__9482 (
            .O(N__43535),
            .I(N__43532));
    Span4Mux_s2_v I__9481 (
            .O(N__43532),
            .I(N__43529));
    Span4Mux_h I__9480 (
            .O(N__43529),
            .I(N__43526));
    Span4Mux_v I__9479 (
            .O(N__43526),
            .I(N__43523));
    Odrv4 I__9478 (
            .O(N__43523),
            .I(RAM_ADD_c_4));
    InMux I__9477 (
            .O(N__43520),
            .I(N__43517));
    LocalMux I__9476 (
            .O(N__43517),
            .I(N__43514));
    Span12Mux_v I__9475 (
            .O(N__43514),
            .I(N__43511));
    Span12Mux_h I__9474 (
            .O(N__43511),
            .I(N__43507));
    InMux I__9473 (
            .O(N__43510),
            .I(N__43504));
    Odrv12 I__9472 (
            .O(N__43507),
            .I(sRAM_pointer_writeZ0Z_3));
    LocalMux I__9471 (
            .O(N__43504),
            .I(sRAM_pointer_writeZ0Z_3));
    InMux I__9470 (
            .O(N__43499),
            .I(N__43478));
    InMux I__9469 (
            .O(N__43498),
            .I(N__43478));
    InMux I__9468 (
            .O(N__43497),
            .I(N__43478));
    InMux I__9467 (
            .O(N__43496),
            .I(N__43478));
    InMux I__9466 (
            .O(N__43495),
            .I(N__43469));
    InMux I__9465 (
            .O(N__43494),
            .I(N__43469));
    InMux I__9464 (
            .O(N__43493),
            .I(N__43469));
    InMux I__9463 (
            .O(N__43492),
            .I(N__43469));
    CascadeMux I__9462 (
            .O(N__43491),
            .I(N__43463));
    CascadeMux I__9461 (
            .O(N__43490),
            .I(N__43459));
    CascadeMux I__9460 (
            .O(N__43489),
            .I(N__43455));
    CascadeMux I__9459 (
            .O(N__43488),
            .I(N__43451));
    CascadeMux I__9458 (
            .O(N__43487),
            .I(N__43447));
    LocalMux I__9457 (
            .O(N__43478),
            .I(N__43440));
    LocalMux I__9456 (
            .O(N__43469),
            .I(N__43440));
    InMux I__9455 (
            .O(N__43468),
            .I(N__43433));
    InMux I__9454 (
            .O(N__43467),
            .I(N__43433));
    InMux I__9453 (
            .O(N__43466),
            .I(N__43430));
    InMux I__9452 (
            .O(N__43463),
            .I(N__43413));
    InMux I__9451 (
            .O(N__43462),
            .I(N__43413));
    InMux I__9450 (
            .O(N__43459),
            .I(N__43413));
    InMux I__9449 (
            .O(N__43458),
            .I(N__43413));
    InMux I__9448 (
            .O(N__43455),
            .I(N__43413));
    InMux I__9447 (
            .O(N__43454),
            .I(N__43413));
    InMux I__9446 (
            .O(N__43451),
            .I(N__43413));
    InMux I__9445 (
            .O(N__43450),
            .I(N__43413));
    InMux I__9444 (
            .O(N__43447),
            .I(N__43408));
    InMux I__9443 (
            .O(N__43446),
            .I(N__43408));
    InMux I__9442 (
            .O(N__43445),
            .I(N__43405));
    Span4Mux_h I__9441 (
            .O(N__43440),
            .I(N__43402));
    InMux I__9440 (
            .O(N__43439),
            .I(N__43399));
    InMux I__9439 (
            .O(N__43438),
            .I(N__43396));
    LocalMux I__9438 (
            .O(N__43433),
            .I(N__43385));
    LocalMux I__9437 (
            .O(N__43430),
            .I(N__43385));
    LocalMux I__9436 (
            .O(N__43413),
            .I(N__43385));
    LocalMux I__9435 (
            .O(N__43408),
            .I(N__43385));
    LocalMux I__9434 (
            .O(N__43405),
            .I(N__43385));
    Odrv4 I__9433 (
            .O(N__43402),
            .I(un1_sacqtime_cry_23_THRU_CO));
    LocalMux I__9432 (
            .O(N__43399),
            .I(un1_sacqtime_cry_23_THRU_CO));
    LocalMux I__9431 (
            .O(N__43396),
            .I(un1_sacqtime_cry_23_THRU_CO));
    Odrv12 I__9430 (
            .O(N__43385),
            .I(un1_sacqtime_cry_23_THRU_CO));
    CascadeMux I__9429 (
            .O(N__43376),
            .I(N__43373));
    InMux I__9428 (
            .O(N__43373),
            .I(N__43370));
    LocalMux I__9427 (
            .O(N__43370),
            .I(N__43367));
    Span12Mux_h I__9426 (
            .O(N__43367),
            .I(N__43363));
    InMux I__9425 (
            .O(N__43366),
            .I(N__43360));
    Odrv12 I__9424 (
            .O(N__43363),
            .I(sRAM_pointer_readZ0Z_3));
    LocalMux I__9423 (
            .O(N__43360),
            .I(sRAM_pointer_readZ0Z_3));
    InMux I__9422 (
            .O(N__43355),
            .I(N__43317));
    InMux I__9421 (
            .O(N__43354),
            .I(N__43317));
    InMux I__9420 (
            .O(N__43353),
            .I(N__43317));
    InMux I__9419 (
            .O(N__43352),
            .I(N__43317));
    InMux I__9418 (
            .O(N__43351),
            .I(N__43317));
    InMux I__9417 (
            .O(N__43350),
            .I(N__43317));
    InMux I__9416 (
            .O(N__43349),
            .I(N__43317));
    InMux I__9415 (
            .O(N__43348),
            .I(N__43317));
    InMux I__9414 (
            .O(N__43347),
            .I(N__43308));
    InMux I__9413 (
            .O(N__43346),
            .I(N__43308));
    InMux I__9412 (
            .O(N__43345),
            .I(N__43308));
    InMux I__9411 (
            .O(N__43344),
            .I(N__43291));
    InMux I__9410 (
            .O(N__43343),
            .I(N__43291));
    InMux I__9409 (
            .O(N__43342),
            .I(N__43291));
    InMux I__9408 (
            .O(N__43341),
            .I(N__43291));
    InMux I__9407 (
            .O(N__43340),
            .I(N__43291));
    InMux I__9406 (
            .O(N__43339),
            .I(N__43291));
    InMux I__9405 (
            .O(N__43338),
            .I(N__43291));
    InMux I__9404 (
            .O(N__43337),
            .I(N__43291));
    InMux I__9403 (
            .O(N__43336),
            .I(N__43286));
    InMux I__9402 (
            .O(N__43335),
            .I(N__43286));
    InMux I__9401 (
            .O(N__43334),
            .I(N__43283));
    LocalMux I__9400 (
            .O(N__43317),
            .I(N__43280));
    InMux I__9399 (
            .O(N__43316),
            .I(N__43277));
    InMux I__9398 (
            .O(N__43315),
            .I(N__43274));
    LocalMux I__9397 (
            .O(N__43308),
            .I(N__43265));
    LocalMux I__9396 (
            .O(N__43291),
            .I(N__43265));
    LocalMux I__9395 (
            .O(N__43286),
            .I(N__43265));
    LocalMux I__9394 (
            .O(N__43283),
            .I(N__43265));
    Span4Mux_h I__9393 (
            .O(N__43280),
            .I(N__43262));
    LocalMux I__9392 (
            .O(N__43277),
            .I(N__43255));
    LocalMux I__9391 (
            .O(N__43274),
            .I(N__43255));
    Span4Mux_h I__9390 (
            .O(N__43265),
            .I(N__43255));
    Span4Mux_h I__9389 (
            .O(N__43262),
            .I(N__43252));
    Span4Mux_h I__9388 (
            .O(N__43255),
            .I(N__43249));
    Odrv4 I__9387 (
            .O(N__43252),
            .I(un4_sacqtime_cry_23_THRU_CO));
    Odrv4 I__9386 (
            .O(N__43249),
            .I(un4_sacqtime_cry_23_THRU_CO));
    IoInMux I__9385 (
            .O(N__43244),
            .I(N__43241));
    LocalMux I__9384 (
            .O(N__43241),
            .I(N__43238));
    Span4Mux_s1_v I__9383 (
            .O(N__43238),
            .I(N__43235));
    Span4Mux_v I__9382 (
            .O(N__43235),
            .I(N__43232));
    Span4Mux_v I__9381 (
            .O(N__43232),
            .I(N__43229));
    Odrv4 I__9380 (
            .O(N__43229),
            .I(RAM_ADD_c_3));
    CEMux I__9379 (
            .O(N__43226),
            .I(N__43222));
    CEMux I__9378 (
            .O(N__43225),
            .I(N__43219));
    LocalMux I__9377 (
            .O(N__43222),
            .I(N__43215));
    LocalMux I__9376 (
            .O(N__43219),
            .I(N__43212));
    CEMux I__9375 (
            .O(N__43218),
            .I(N__43209));
    Span4Mux_v I__9374 (
            .O(N__43215),
            .I(N__43206));
    Span4Mux_h I__9373 (
            .O(N__43212),
            .I(N__43203));
    LocalMux I__9372 (
            .O(N__43209),
            .I(N__43200));
    Span4Mux_h I__9371 (
            .O(N__43206),
            .I(N__43193));
    Span4Mux_h I__9370 (
            .O(N__43203),
            .I(N__43193));
    Span4Mux_v I__9369 (
            .O(N__43200),
            .I(N__43193));
    Odrv4 I__9368 (
            .O(N__43193),
            .I(N_67_i));
    IoInMux I__9367 (
            .O(N__43190),
            .I(N__43187));
    LocalMux I__9366 (
            .O(N__43187),
            .I(N__43184));
    Span12Mux_s8_v I__9365 (
            .O(N__43184),
            .I(N__43180));
    InMux I__9364 (
            .O(N__43183),
            .I(N__43177));
    Odrv12 I__9363 (
            .O(N__43180),
            .I(RAM_DATA_cl_13Z0Z_15));
    LocalMux I__9362 (
            .O(N__43177),
            .I(RAM_DATA_cl_13Z0Z_15));
    IoInMux I__9361 (
            .O(N__43172),
            .I(N__43169));
    LocalMux I__9360 (
            .O(N__43169),
            .I(N__43166));
    Span4Mux_s2_v I__9359 (
            .O(N__43166),
            .I(N__43163));
    Span4Mux_h I__9358 (
            .O(N__43163),
            .I(N__43160));
    Span4Mux_h I__9357 (
            .O(N__43160),
            .I(N__43156));
    CascadeMux I__9356 (
            .O(N__43159),
            .I(N__43153));
    Span4Mux_v I__9355 (
            .O(N__43156),
            .I(N__43150));
    InMux I__9354 (
            .O(N__43153),
            .I(N__43147));
    Odrv4 I__9353 (
            .O(N__43150),
            .I(RAM_DATA_cl_14Z0Z_15));
    LocalMux I__9352 (
            .O(N__43147),
            .I(RAM_DATA_cl_14Z0Z_15));
    IoInMux I__9351 (
            .O(N__43142),
            .I(N__43139));
    LocalMux I__9350 (
            .O(N__43139),
            .I(N__43136));
    Span4Mux_s3_h I__9349 (
            .O(N__43136),
            .I(N__43133));
    Span4Mux_v I__9348 (
            .O(N__43133),
            .I(N__43130));
    Span4Mux_v I__9347 (
            .O(N__43130),
            .I(N__43127));
    Span4Mux_h I__9346 (
            .O(N__43127),
            .I(N__43123));
    InMux I__9345 (
            .O(N__43126),
            .I(N__43120));
    Odrv4 I__9344 (
            .O(N__43123),
            .I(RAM_DATA_cl_15Z0Z_15));
    LocalMux I__9343 (
            .O(N__43120),
            .I(RAM_DATA_cl_15Z0Z_15));
    IoInMux I__9342 (
            .O(N__43115),
            .I(N__43112));
    LocalMux I__9341 (
            .O(N__43112),
            .I(N__43109));
    IoSpan4Mux I__9340 (
            .O(N__43109),
            .I(N__43106));
    Span4Mux_s2_h I__9339 (
            .O(N__43106),
            .I(N__43103));
    Sp12to4 I__9338 (
            .O(N__43103),
            .I(N__43100));
    Span12Mux_s10_h I__9337 (
            .O(N__43100),
            .I(N__43096));
    CascadeMux I__9336 (
            .O(N__43099),
            .I(N__43093));
    Span12Mux_v I__9335 (
            .O(N__43096),
            .I(N__43090));
    InMux I__9334 (
            .O(N__43093),
            .I(N__43087));
    Odrv12 I__9333 (
            .O(N__43090),
            .I(RAM_DATA_cl_1Z0Z_15));
    LocalMux I__9332 (
            .O(N__43087),
            .I(RAM_DATA_cl_1Z0Z_15));
    InMux I__9331 (
            .O(N__43082),
            .I(sCounterADC_cry_2));
    InMux I__9330 (
            .O(N__43079),
            .I(N__43076));
    LocalMux I__9329 (
            .O(N__43076),
            .I(N__43073));
    Span4Mux_v I__9328 (
            .O(N__43073),
            .I(N__43070));
    Span4Mux_h I__9327 (
            .O(N__43070),
            .I(N__43066));
    InMux I__9326 (
            .O(N__43069),
            .I(N__43063));
    Span4Mux_h I__9325 (
            .O(N__43066),
            .I(N__43060));
    LocalMux I__9324 (
            .O(N__43063),
            .I(sCounterADCZ0Z_4));
    Odrv4 I__9323 (
            .O(N__43060),
            .I(sCounterADCZ0Z_4));
    InMux I__9322 (
            .O(N__43055),
            .I(sCounterADC_cry_3));
    InMux I__9321 (
            .O(N__43052),
            .I(N__43049));
    LocalMux I__9320 (
            .O(N__43049),
            .I(N__43046));
    Span4Mux_v I__9319 (
            .O(N__43046),
            .I(N__43043));
    Span4Mux_h I__9318 (
            .O(N__43043),
            .I(N__43039));
    InMux I__9317 (
            .O(N__43042),
            .I(N__43036));
    Span4Mux_h I__9316 (
            .O(N__43039),
            .I(N__43033));
    LocalMux I__9315 (
            .O(N__43036),
            .I(sCounterADCZ0Z_5));
    Odrv4 I__9314 (
            .O(N__43033),
            .I(sCounterADCZ0Z_5));
    InMux I__9313 (
            .O(N__43028),
            .I(sCounterADC_cry_4));
    InMux I__9312 (
            .O(N__43025),
            .I(sCounterADC_cry_5));
    InMux I__9311 (
            .O(N__43022),
            .I(sCounterADC_cry_6));
    InMux I__9310 (
            .O(N__43019),
            .I(N__43016));
    LocalMux I__9309 (
            .O(N__43016),
            .I(N__43013));
    Span4Mux_v I__9308 (
            .O(N__43013),
            .I(N__43010));
    Sp12to4 I__9307 (
            .O(N__43010),
            .I(N__43007));
    Span12Mux_h I__9306 (
            .O(N__43007),
            .I(N__43004));
    Odrv12 I__9305 (
            .O(N__43004),
            .I(RAM_DATA_in_5));
    InMux I__9304 (
            .O(N__43001),
            .I(N__42998));
    LocalMux I__9303 (
            .O(N__42998),
            .I(N__42995));
    Span12Mux_v I__9302 (
            .O(N__42995),
            .I(N__42992));
    Odrv12 I__9301 (
            .O(N__42992),
            .I(RAM_DATA_in_13));
    InMux I__9300 (
            .O(N__42989),
            .I(N__42986));
    LocalMux I__9299 (
            .O(N__42986),
            .I(N__42983));
    Odrv4 I__9298 (
            .O(N__42983),
            .I(spi_data_misoZ0Z_5));
    InMux I__9297 (
            .O(N__42980),
            .I(N__42977));
    LocalMux I__9296 (
            .O(N__42977),
            .I(N__42974));
    Span12Mux_v I__9295 (
            .O(N__42974),
            .I(N__42971));
    Odrv12 I__9294 (
            .O(N__42971),
            .I(RAM_DATA_in_15));
    CascadeMux I__9293 (
            .O(N__42968),
            .I(N__42965));
    InMux I__9292 (
            .O(N__42965),
            .I(N__42962));
    LocalMux I__9291 (
            .O(N__42962),
            .I(N__42959));
    Span4Mux_v I__9290 (
            .O(N__42959),
            .I(N__42956));
    Span4Mux_v I__9289 (
            .O(N__42956),
            .I(N__42953));
    Span4Mux_h I__9288 (
            .O(N__42953),
            .I(N__42950));
    Span4Mux_h I__9287 (
            .O(N__42950),
            .I(N__42947));
    Odrv4 I__9286 (
            .O(N__42947),
            .I(RAM_DATA_in_7));
    InMux I__9285 (
            .O(N__42944),
            .I(N__42941));
    LocalMux I__9284 (
            .O(N__42941),
            .I(N__42938));
    Odrv4 I__9283 (
            .O(N__42938),
            .I(spi_data_misoZ0Z_7));
    InMux I__9282 (
            .O(N__42935),
            .I(N__42932));
    LocalMux I__9281 (
            .O(N__42932),
            .I(N__42929));
    Span4Mux_v I__9280 (
            .O(N__42929),
            .I(N__42926));
    Sp12to4 I__9279 (
            .O(N__42926),
            .I(N__42923));
    Span12Mux_h I__9278 (
            .O(N__42923),
            .I(N__42920));
    Odrv12 I__9277 (
            .O(N__42920),
            .I(RAM_DATA_in_3));
    CascadeMux I__9276 (
            .O(N__42917),
            .I(N__42914));
    InMux I__9275 (
            .O(N__42914),
            .I(N__42911));
    LocalMux I__9274 (
            .O(N__42911),
            .I(N__42908));
    Span4Mux_h I__9273 (
            .O(N__42908),
            .I(N__42905));
    Sp12to4 I__9272 (
            .O(N__42905),
            .I(N__42902));
    Span12Mux_v I__9271 (
            .O(N__42902),
            .I(N__42899));
    Odrv12 I__9270 (
            .O(N__42899),
            .I(RAM_DATA_in_11));
    InMux I__9269 (
            .O(N__42896),
            .I(N__42893));
    LocalMux I__9268 (
            .O(N__42893),
            .I(N__42890));
    Odrv4 I__9267 (
            .O(N__42890),
            .I(spi_data_misoZ0Z_3));
    InMux I__9266 (
            .O(N__42887),
            .I(N__42884));
    LocalMux I__9265 (
            .O(N__42884),
            .I(N__42881));
    Span12Mux_v I__9264 (
            .O(N__42881),
            .I(N__42878));
    Span12Mux_v I__9263 (
            .O(N__42878),
            .I(N__42875));
    Odrv12 I__9262 (
            .O(N__42875),
            .I(RAM_DATA_in_10));
    InMux I__9261 (
            .O(N__42872),
            .I(N__42869));
    LocalMux I__9260 (
            .O(N__42869),
            .I(N__42866));
    Span4Mux_v I__9259 (
            .O(N__42866),
            .I(N__42863));
    Sp12to4 I__9258 (
            .O(N__42863),
            .I(N__42860));
    Span12Mux_h I__9257 (
            .O(N__42860),
            .I(N__42857));
    Odrv12 I__9256 (
            .O(N__42857),
            .I(RAM_DATA_in_2));
    InMux I__9255 (
            .O(N__42854),
            .I(N__42851));
    LocalMux I__9254 (
            .O(N__42851),
            .I(N__42848));
    Odrv4 I__9253 (
            .O(N__42848),
            .I(spi_data_misoZ0Z_2));
    InMux I__9252 (
            .O(N__42845),
            .I(N__42842));
    LocalMux I__9251 (
            .O(N__42842),
            .I(N__42839));
    Odrv4 I__9250 (
            .O(N__42839),
            .I(spi_data_misoZ0Z_4));
    InMux I__9249 (
            .O(N__42836),
            .I(N__42833));
    LocalMux I__9248 (
            .O(N__42833),
            .I(spi_data_misoZ0Z_6));
    CEMux I__9247 (
            .O(N__42830),
            .I(N__42827));
    LocalMux I__9246 (
            .O(N__42827),
            .I(N__42824));
    Span4Mux_v I__9245 (
            .O(N__42824),
            .I(N__42821));
    Span4Mux_v I__9244 (
            .O(N__42821),
            .I(N__42818));
    Sp12to4 I__9243 (
            .O(N__42818),
            .I(N__42815));
    Odrv12 I__9242 (
            .O(N__42815),
            .I(\spi_slave_inst.un4_i_wr ));
    InMux I__9241 (
            .O(N__42812),
            .I(bfn_18_15_0_));
    InMux I__9240 (
            .O(N__42809),
            .I(sCounterADC_cry_0));
    InMux I__9239 (
            .O(N__42806),
            .I(sCounterADC_cry_1));
    InMux I__9238 (
            .O(N__42803),
            .I(N__42800));
    LocalMux I__9237 (
            .O(N__42800),
            .I(N__42797));
    Span4Mux_h I__9236 (
            .O(N__42797),
            .I(N__42794));
    Odrv4 I__9235 (
            .O(N__42794),
            .I(sDAC_mem_25Z0Z_7));
    CascadeMux I__9234 (
            .O(N__42791),
            .I(N__42788));
    InMux I__9233 (
            .O(N__42788),
            .I(N__42784));
    InMux I__9232 (
            .O(N__42787),
            .I(N__42781));
    LocalMux I__9231 (
            .O(N__42784),
            .I(N__42776));
    LocalMux I__9230 (
            .O(N__42781),
            .I(N__42776));
    Odrv12 I__9229 (
            .O(N__42776),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa ));
    InMux I__9228 (
            .O(N__42773),
            .I(N__42769));
    CascadeMux I__9227 (
            .O(N__42772),
            .I(N__42765));
    LocalMux I__9226 (
            .O(N__42769),
            .I(N__42762));
    InMux I__9225 (
            .O(N__42768),
            .I(N__42759));
    InMux I__9224 (
            .O(N__42765),
            .I(N__42756));
    Span12Mux_h I__9223 (
            .O(N__42762),
            .I(N__42753));
    LocalMux I__9222 (
            .O(N__42759),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0 ));
    LocalMux I__9221 (
            .O(N__42756),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0 ));
    Odrv12 I__9220 (
            .O(N__42753),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0 ));
    InMux I__9219 (
            .O(N__42746),
            .I(N__42743));
    LocalMux I__9218 (
            .O(N__42743),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO ));
    CascadeMux I__9217 (
            .O(N__42740),
            .I(N__42737));
    InMux I__9216 (
            .O(N__42737),
            .I(N__42733));
    CascadeMux I__9215 (
            .O(N__42736),
            .I(N__42730));
    LocalMux I__9214 (
            .O(N__42733),
            .I(N__42726));
    InMux I__9213 (
            .O(N__42730),
            .I(N__42723));
    InMux I__9212 (
            .O(N__42729),
            .I(N__42720));
    Span12Mux_h I__9211 (
            .O(N__42726),
            .I(N__42717));
    LocalMux I__9210 (
            .O(N__42723),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1 ));
    LocalMux I__9209 (
            .O(N__42720),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1 ));
    Odrv12 I__9208 (
            .O(N__42717),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1 ));
    CascadeMux I__9207 (
            .O(N__42710),
            .I(N__42707));
    InMux I__9206 (
            .O(N__42707),
            .I(N__42702));
    InMux I__9205 (
            .O(N__42706),
            .I(N__42697));
    InMux I__9204 (
            .O(N__42705),
            .I(N__42697));
    LocalMux I__9203 (
            .O(N__42702),
            .I(N__42692));
    LocalMux I__9202 (
            .O(N__42697),
            .I(N__42692));
    Odrv12 I__9201 (
            .O(N__42692),
            .I(\spi_slave_inst.un23_i_ssn ));
    InMux I__9200 (
            .O(N__42689),
            .I(N__42686));
    LocalMux I__9199 (
            .O(N__42686),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO ));
    InMux I__9198 (
            .O(N__42683),
            .I(N__42680));
    LocalMux I__9197 (
            .O(N__42680),
            .I(N__42675));
    InMux I__9196 (
            .O(N__42679),
            .I(N__42672));
    InMux I__9195 (
            .O(N__42678),
            .I(N__42669));
    Span12Mux_h I__9194 (
            .O(N__42675),
            .I(N__42666));
    LocalMux I__9193 (
            .O(N__42672),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2 ));
    LocalMux I__9192 (
            .O(N__42669),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2 ));
    Odrv12 I__9191 (
            .O(N__42666),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2 ));
    InMux I__9190 (
            .O(N__42659),
            .I(N__42656));
    LocalMux I__9189 (
            .O(N__42656),
            .I(N__42653));
    Odrv4 I__9188 (
            .O(N__42653),
            .I(spi_data_misoZ0Z_0));
    CascadeMux I__9187 (
            .O(N__42650),
            .I(N__42647));
    InMux I__9186 (
            .O(N__42647),
            .I(N__42644));
    LocalMux I__9185 (
            .O(N__42644),
            .I(sDAC_mem_4Z0Z_1));
    CEMux I__9184 (
            .O(N__42641),
            .I(N__42637));
    CEMux I__9183 (
            .O(N__42640),
            .I(N__42633));
    LocalMux I__9182 (
            .O(N__42637),
            .I(N__42630));
    CEMux I__9181 (
            .O(N__42636),
            .I(N__42627));
    LocalMux I__9180 (
            .O(N__42633),
            .I(N__42619));
    Span4Mux_h I__9179 (
            .O(N__42630),
            .I(N__42619));
    LocalMux I__9178 (
            .O(N__42627),
            .I(N__42619));
    CEMux I__9177 (
            .O(N__42626),
            .I(N__42616));
    Span4Mux_v I__9176 (
            .O(N__42619),
            .I(N__42613));
    LocalMux I__9175 (
            .O(N__42616),
            .I(N__42610));
    Span4Mux_h I__9174 (
            .O(N__42613),
            .I(N__42607));
    Span12Mux_h I__9173 (
            .O(N__42610),
            .I(N__42604));
    Sp12to4 I__9172 (
            .O(N__42607),
            .I(N__42601));
    Odrv12 I__9171 (
            .O(N__42604),
            .I(sDAC_mem_4_1_sqmuxa));
    Odrv12 I__9170 (
            .O(N__42601),
            .I(sDAC_mem_4_1_sqmuxa));
    CascadeMux I__9169 (
            .O(N__42596),
            .I(N__42592));
    CascadeMux I__9168 (
            .O(N__42595),
            .I(N__42589));
    InMux I__9167 (
            .O(N__42592),
            .I(N__42581));
    InMux I__9166 (
            .O(N__42589),
            .I(N__42581));
    InMux I__9165 (
            .O(N__42588),
            .I(N__42581));
    LocalMux I__9164 (
            .O(N__42581),
            .I(N__42577));
    CascadeMux I__9163 (
            .O(N__42580),
            .I(N__42571));
    Span4Mux_v I__9162 (
            .O(N__42577),
            .I(N__42563));
    InMux I__9161 (
            .O(N__42576),
            .I(N__42560));
    CascadeMux I__9160 (
            .O(N__42575),
            .I(N__42553));
    CascadeMux I__9159 (
            .O(N__42574),
            .I(N__42546));
    InMux I__9158 (
            .O(N__42571),
            .I(N__42538));
    InMux I__9157 (
            .O(N__42570),
            .I(N__42538));
    InMux I__9156 (
            .O(N__42569),
            .I(N__42538));
    InMux I__9155 (
            .O(N__42568),
            .I(N__42533));
    InMux I__9154 (
            .O(N__42567),
            .I(N__42533));
    InMux I__9153 (
            .O(N__42566),
            .I(N__42530));
    Span4Mux_h I__9152 (
            .O(N__42563),
            .I(N__42516));
    LocalMux I__9151 (
            .O(N__42560),
            .I(N__42516));
    InMux I__9150 (
            .O(N__42559),
            .I(N__42507));
    InMux I__9149 (
            .O(N__42558),
            .I(N__42500));
    InMux I__9148 (
            .O(N__42557),
            .I(N__42500));
    InMux I__9147 (
            .O(N__42556),
            .I(N__42500));
    InMux I__9146 (
            .O(N__42553),
            .I(N__42493));
    InMux I__9145 (
            .O(N__42552),
            .I(N__42493));
    InMux I__9144 (
            .O(N__42551),
            .I(N__42493));
    InMux I__9143 (
            .O(N__42550),
            .I(N__42490));
    InMux I__9142 (
            .O(N__42549),
            .I(N__42483));
    InMux I__9141 (
            .O(N__42546),
            .I(N__42483));
    InMux I__9140 (
            .O(N__42545),
            .I(N__42483));
    LocalMux I__9139 (
            .O(N__42538),
            .I(N__42478));
    LocalMux I__9138 (
            .O(N__42533),
            .I(N__42478));
    LocalMux I__9137 (
            .O(N__42530),
            .I(N__42475));
    InMux I__9136 (
            .O(N__42529),
            .I(N__42470));
    InMux I__9135 (
            .O(N__42528),
            .I(N__42470));
    InMux I__9134 (
            .O(N__42527),
            .I(N__42465));
    InMux I__9133 (
            .O(N__42526),
            .I(N__42465));
    InMux I__9132 (
            .O(N__42525),
            .I(N__42462));
    InMux I__9131 (
            .O(N__42524),
            .I(N__42455));
    InMux I__9130 (
            .O(N__42523),
            .I(N__42455));
    InMux I__9129 (
            .O(N__42522),
            .I(N__42455));
    InMux I__9128 (
            .O(N__42521),
            .I(N__42452));
    Span4Mux_v I__9127 (
            .O(N__42516),
            .I(N__42449));
    InMux I__9126 (
            .O(N__42515),
            .I(N__42446));
    InMux I__9125 (
            .O(N__42514),
            .I(N__42441));
    InMux I__9124 (
            .O(N__42513),
            .I(N__42441));
    InMux I__9123 (
            .O(N__42512),
            .I(N__42434));
    InMux I__9122 (
            .O(N__42511),
            .I(N__42434));
    InMux I__9121 (
            .O(N__42510),
            .I(N__42434));
    LocalMux I__9120 (
            .O(N__42507),
            .I(N__42418));
    LocalMux I__9119 (
            .O(N__42500),
            .I(N__42415));
    LocalMux I__9118 (
            .O(N__42493),
            .I(N__42412));
    LocalMux I__9117 (
            .O(N__42490),
            .I(N__42408));
    LocalMux I__9116 (
            .O(N__42483),
            .I(N__42403));
    Span4Mux_v I__9115 (
            .O(N__42478),
            .I(N__42403));
    Span4Mux_v I__9114 (
            .O(N__42475),
            .I(N__42400));
    LocalMux I__9113 (
            .O(N__42470),
            .I(N__42395));
    LocalMux I__9112 (
            .O(N__42465),
            .I(N__42395));
    LocalMux I__9111 (
            .O(N__42462),
            .I(N__42388));
    LocalMux I__9110 (
            .O(N__42455),
            .I(N__42388));
    LocalMux I__9109 (
            .O(N__42452),
            .I(N__42388));
    Span4Mux_h I__9108 (
            .O(N__42449),
            .I(N__42379));
    LocalMux I__9107 (
            .O(N__42446),
            .I(N__42379));
    LocalMux I__9106 (
            .O(N__42441),
            .I(N__42379));
    LocalMux I__9105 (
            .O(N__42434),
            .I(N__42379));
    InMux I__9104 (
            .O(N__42433),
            .I(N__42376));
    InMux I__9103 (
            .O(N__42432),
            .I(N__42373));
    InMux I__9102 (
            .O(N__42431),
            .I(N__42370));
    InMux I__9101 (
            .O(N__42430),
            .I(N__42367));
    InMux I__9100 (
            .O(N__42429),
            .I(N__42360));
    InMux I__9099 (
            .O(N__42428),
            .I(N__42360));
    InMux I__9098 (
            .O(N__42427),
            .I(N__42360));
    InMux I__9097 (
            .O(N__42426),
            .I(N__42357));
    InMux I__9096 (
            .O(N__42425),
            .I(N__42352));
    InMux I__9095 (
            .O(N__42424),
            .I(N__42352));
    InMux I__9094 (
            .O(N__42423),
            .I(N__42347));
    InMux I__9093 (
            .O(N__42422),
            .I(N__42347));
    InMux I__9092 (
            .O(N__42421),
            .I(N__42344));
    Span4Mux_h I__9091 (
            .O(N__42418),
            .I(N__42337));
    Span4Mux_v I__9090 (
            .O(N__42415),
            .I(N__42337));
    Span4Mux_v I__9089 (
            .O(N__42412),
            .I(N__42337));
    InMux I__9088 (
            .O(N__42411),
            .I(N__42334));
    Span4Mux_v I__9087 (
            .O(N__42408),
            .I(N__42325));
    Span4Mux_h I__9086 (
            .O(N__42403),
            .I(N__42325));
    Span4Mux_h I__9085 (
            .O(N__42400),
            .I(N__42325));
    Span4Mux_v I__9084 (
            .O(N__42395),
            .I(N__42325));
    Span4Mux_v I__9083 (
            .O(N__42388),
            .I(N__42320));
    Span4Mux_v I__9082 (
            .O(N__42379),
            .I(N__42320));
    LocalMux I__9081 (
            .O(N__42376),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9080 (
            .O(N__42373),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9079 (
            .O(N__42370),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9078 (
            .O(N__42367),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9077 (
            .O(N__42360),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9076 (
            .O(N__42357),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9075 (
            .O(N__42352),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9074 (
            .O(N__42347),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9073 (
            .O(N__42344),
            .I(sDAC_mem_pointerZ0Z_5));
    Odrv4 I__9072 (
            .O(N__42337),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9071 (
            .O(N__42334),
            .I(sDAC_mem_pointerZ0Z_5));
    Odrv4 I__9070 (
            .O(N__42325),
            .I(sDAC_mem_pointerZ0Z_5));
    Odrv4 I__9069 (
            .O(N__42320),
            .I(sDAC_mem_pointerZ0Z_5));
    InMux I__9068 (
            .O(N__42293),
            .I(N__42290));
    LocalMux I__9067 (
            .O(N__42290),
            .I(N__42287));
    Span4Mux_v I__9066 (
            .O(N__42287),
            .I(N__42284));
    Span4Mux_v I__9065 (
            .O(N__42284),
            .I(N__42281));
    Odrv4 I__9064 (
            .O(N__42281),
            .I(sDAC_mem_36Z0Z_2));
    InMux I__9063 (
            .O(N__42278),
            .I(N__42275));
    LocalMux I__9062 (
            .O(N__42275),
            .I(N__42272));
    Span12Mux_s11_h I__9061 (
            .O(N__42272),
            .I(N__42269));
    Odrv12 I__9060 (
            .O(N__42269),
            .I(sDAC_mem_4Z0Z_2));
    CascadeMux I__9059 (
            .O(N__42266),
            .I(N__42260));
    CascadeMux I__9058 (
            .O(N__42265),
            .I(N__42256));
    CascadeMux I__9057 (
            .O(N__42264),
            .I(N__42253));
    CascadeMux I__9056 (
            .O(N__42263),
            .I(N__42250));
    InMux I__9055 (
            .O(N__42260),
            .I(N__42235));
    InMux I__9054 (
            .O(N__42259),
            .I(N__42222));
    InMux I__9053 (
            .O(N__42256),
            .I(N__42222));
    InMux I__9052 (
            .O(N__42253),
            .I(N__42222));
    InMux I__9051 (
            .O(N__42250),
            .I(N__42219));
    CascadeMux I__9050 (
            .O(N__42249),
            .I(N__42215));
    CascadeMux I__9049 (
            .O(N__42248),
            .I(N__42206));
    CascadeMux I__9048 (
            .O(N__42247),
            .I(N__42199));
    CascadeMux I__9047 (
            .O(N__42246),
            .I(N__42194));
    CascadeMux I__9046 (
            .O(N__42245),
            .I(N__42185));
    CascadeMux I__9045 (
            .O(N__42244),
            .I(N__42182));
    InMux I__9044 (
            .O(N__42243),
            .I(N__42176));
    InMux I__9043 (
            .O(N__42242),
            .I(N__42176));
    CascadeMux I__9042 (
            .O(N__42241),
            .I(N__42162));
    CascadeMux I__9041 (
            .O(N__42240),
            .I(N__42158));
    CascadeMux I__9040 (
            .O(N__42239),
            .I(N__42154));
    CascadeMux I__9039 (
            .O(N__42238),
            .I(N__42150));
    LocalMux I__9038 (
            .O(N__42235),
            .I(N__42139));
    InMux I__9037 (
            .O(N__42234),
            .I(N__42132));
    InMux I__9036 (
            .O(N__42233),
            .I(N__42132));
    InMux I__9035 (
            .O(N__42232),
            .I(N__42132));
    InMux I__9034 (
            .O(N__42231),
            .I(N__42125));
    InMux I__9033 (
            .O(N__42230),
            .I(N__42125));
    InMux I__9032 (
            .O(N__42229),
            .I(N__42125));
    LocalMux I__9031 (
            .O(N__42222),
            .I(N__42120));
    LocalMux I__9030 (
            .O(N__42219),
            .I(N__42120));
    InMux I__9029 (
            .O(N__42218),
            .I(N__42115));
    InMux I__9028 (
            .O(N__42215),
            .I(N__42115));
    CascadeMux I__9027 (
            .O(N__42214),
            .I(N__42106));
    CascadeMux I__9026 (
            .O(N__42213),
            .I(N__42101));
    CascadeMux I__9025 (
            .O(N__42212),
            .I(N__42098));
    InMux I__9024 (
            .O(N__42211),
            .I(N__42090));
    InMux I__9023 (
            .O(N__42210),
            .I(N__42083));
    InMux I__9022 (
            .O(N__42209),
            .I(N__42083));
    InMux I__9021 (
            .O(N__42206),
            .I(N__42083));
    CascadeMux I__9020 (
            .O(N__42205),
            .I(N__42077));
    CascadeMux I__9019 (
            .O(N__42204),
            .I(N__42069));
    CascadeMux I__9018 (
            .O(N__42203),
            .I(N__42064));
    InMux I__9017 (
            .O(N__42202),
            .I(N__42053));
    InMux I__9016 (
            .O(N__42199),
            .I(N__42053));
    InMux I__9015 (
            .O(N__42198),
            .I(N__42053));
    InMux I__9014 (
            .O(N__42197),
            .I(N__42053));
    InMux I__9013 (
            .O(N__42194),
            .I(N__42053));
    CascadeMux I__9012 (
            .O(N__42193),
            .I(N__42049));
    CascadeMux I__9011 (
            .O(N__42192),
            .I(N__42046));
    InMux I__9010 (
            .O(N__42191),
            .I(N__42039));
    InMux I__9009 (
            .O(N__42190),
            .I(N__42039));
    InMux I__9008 (
            .O(N__42189),
            .I(N__42039));
    InMux I__9007 (
            .O(N__42188),
            .I(N__42029));
    InMux I__9006 (
            .O(N__42185),
            .I(N__42022));
    InMux I__9005 (
            .O(N__42182),
            .I(N__42022));
    InMux I__9004 (
            .O(N__42181),
            .I(N__42022));
    LocalMux I__9003 (
            .O(N__42176),
            .I(N__42019));
    CascadeMux I__9002 (
            .O(N__42175),
            .I(N__42007));
    CascadeMux I__9001 (
            .O(N__42174),
            .I(N__42003));
    CascadeMux I__9000 (
            .O(N__42173),
            .I(N__41997));
    CascadeMux I__8999 (
            .O(N__42172),
            .I(N__41994));
    CascadeMux I__8998 (
            .O(N__42171),
            .I(N__41991));
    CascadeMux I__8997 (
            .O(N__42170),
            .I(N__41979));
    CascadeMux I__8996 (
            .O(N__42169),
            .I(N__41976));
    InMux I__8995 (
            .O(N__42168),
            .I(N__41972));
    InMux I__8994 (
            .O(N__42167),
            .I(N__41965));
    InMux I__8993 (
            .O(N__42166),
            .I(N__41965));
    InMux I__8992 (
            .O(N__42165),
            .I(N__41965));
    InMux I__8991 (
            .O(N__42162),
            .I(N__41958));
    InMux I__8990 (
            .O(N__42161),
            .I(N__41958));
    InMux I__8989 (
            .O(N__42158),
            .I(N__41958));
    InMux I__8988 (
            .O(N__42157),
            .I(N__41953));
    InMux I__8987 (
            .O(N__42154),
            .I(N__41953));
    InMux I__8986 (
            .O(N__42153),
            .I(N__41944));
    InMux I__8985 (
            .O(N__42150),
            .I(N__41944));
    InMux I__8984 (
            .O(N__42149),
            .I(N__41944));
    InMux I__8983 (
            .O(N__42148),
            .I(N__41944));
    InMux I__8982 (
            .O(N__42147),
            .I(N__41937));
    InMux I__8981 (
            .O(N__42146),
            .I(N__41937));
    InMux I__8980 (
            .O(N__42145),
            .I(N__41937));
    InMux I__8979 (
            .O(N__42144),
            .I(N__41932));
    InMux I__8978 (
            .O(N__42143),
            .I(N__41932));
    InMux I__8977 (
            .O(N__42142),
            .I(N__41929));
    Span4Mux_v I__8976 (
            .O(N__42139),
            .I(N__41918));
    LocalMux I__8975 (
            .O(N__42132),
            .I(N__41918));
    LocalMux I__8974 (
            .O(N__42125),
            .I(N__41918));
    Span4Mux_h I__8973 (
            .O(N__42120),
            .I(N__41918));
    LocalMux I__8972 (
            .O(N__42115),
            .I(N__41918));
    InMux I__8971 (
            .O(N__42114),
            .I(N__41911));
    InMux I__8970 (
            .O(N__42113),
            .I(N__41911));
    InMux I__8969 (
            .O(N__42112),
            .I(N__41911));
    InMux I__8968 (
            .O(N__42111),
            .I(N__41898));
    InMux I__8967 (
            .O(N__42110),
            .I(N__41898));
    InMux I__8966 (
            .O(N__42109),
            .I(N__41898));
    InMux I__8965 (
            .O(N__42106),
            .I(N__41898));
    InMux I__8964 (
            .O(N__42105),
            .I(N__41898));
    InMux I__8963 (
            .O(N__42104),
            .I(N__41898));
    InMux I__8962 (
            .O(N__42101),
            .I(N__41893));
    InMux I__8961 (
            .O(N__42098),
            .I(N__41893));
    CascadeMux I__8960 (
            .O(N__42097),
            .I(N__41888));
    InMux I__8959 (
            .O(N__42096),
            .I(N__41879));
    InMux I__8958 (
            .O(N__42095),
            .I(N__41879));
    InMux I__8957 (
            .O(N__42094),
            .I(N__41876));
    InMux I__8956 (
            .O(N__42093),
            .I(N__41869));
    LocalMux I__8955 (
            .O(N__42090),
            .I(N__41856));
    LocalMux I__8954 (
            .O(N__42083),
            .I(N__41856));
    InMux I__8953 (
            .O(N__42082),
            .I(N__41851));
    InMux I__8952 (
            .O(N__42081),
            .I(N__41851));
    InMux I__8951 (
            .O(N__42080),
            .I(N__41842));
    InMux I__8950 (
            .O(N__42077),
            .I(N__41842));
    InMux I__8949 (
            .O(N__42076),
            .I(N__41842));
    InMux I__8948 (
            .O(N__42075),
            .I(N__41842));
    CascadeMux I__8947 (
            .O(N__42074),
            .I(N__41838));
    InMux I__8946 (
            .O(N__42073),
            .I(N__41831));
    InMux I__8945 (
            .O(N__42072),
            .I(N__41831));
    InMux I__8944 (
            .O(N__42069),
            .I(N__41831));
    InMux I__8943 (
            .O(N__42068),
            .I(N__41824));
    InMux I__8942 (
            .O(N__42067),
            .I(N__41824));
    InMux I__8941 (
            .O(N__42064),
            .I(N__41824));
    LocalMux I__8940 (
            .O(N__42053),
            .I(N__41821));
    InMux I__8939 (
            .O(N__42052),
            .I(N__41814));
    InMux I__8938 (
            .O(N__42049),
            .I(N__41814));
    InMux I__8937 (
            .O(N__42046),
            .I(N__41814));
    LocalMux I__8936 (
            .O(N__42039),
            .I(N__41801));
    InMux I__8935 (
            .O(N__42038),
            .I(N__41792));
    InMux I__8934 (
            .O(N__42037),
            .I(N__41792));
    InMux I__8933 (
            .O(N__42036),
            .I(N__41792));
    InMux I__8932 (
            .O(N__42035),
            .I(N__41792));
    InMux I__8931 (
            .O(N__42034),
            .I(N__41785));
    InMux I__8930 (
            .O(N__42033),
            .I(N__41785));
    InMux I__8929 (
            .O(N__42032),
            .I(N__41785));
    LocalMux I__8928 (
            .O(N__42029),
            .I(N__41780));
    LocalMux I__8927 (
            .O(N__42022),
            .I(N__41780));
    Span4Mux_v I__8926 (
            .O(N__42019),
            .I(N__41777));
    InMux I__8925 (
            .O(N__42018),
            .I(N__41768));
    InMux I__8924 (
            .O(N__42017),
            .I(N__41768));
    InMux I__8923 (
            .O(N__42016),
            .I(N__41768));
    InMux I__8922 (
            .O(N__42015),
            .I(N__41768));
    InMux I__8921 (
            .O(N__42014),
            .I(N__41763));
    InMux I__8920 (
            .O(N__42013),
            .I(N__41763));
    InMux I__8919 (
            .O(N__42012),
            .I(N__41756));
    InMux I__8918 (
            .O(N__42011),
            .I(N__41756));
    InMux I__8917 (
            .O(N__42010),
            .I(N__41756));
    InMux I__8916 (
            .O(N__42007),
            .I(N__41749));
    InMux I__8915 (
            .O(N__42006),
            .I(N__41749));
    InMux I__8914 (
            .O(N__42003),
            .I(N__41749));
    InMux I__8913 (
            .O(N__42002),
            .I(N__41744));
    InMux I__8912 (
            .O(N__42001),
            .I(N__41744));
    InMux I__8911 (
            .O(N__42000),
            .I(N__41735));
    InMux I__8910 (
            .O(N__41997),
            .I(N__41735));
    InMux I__8909 (
            .O(N__41994),
            .I(N__41735));
    InMux I__8908 (
            .O(N__41991),
            .I(N__41735));
    InMux I__8907 (
            .O(N__41990),
            .I(N__41730));
    InMux I__8906 (
            .O(N__41989),
            .I(N__41730));
    InMux I__8905 (
            .O(N__41988),
            .I(N__41723));
    InMux I__8904 (
            .O(N__41987),
            .I(N__41723));
    InMux I__8903 (
            .O(N__41986),
            .I(N__41723));
    InMux I__8902 (
            .O(N__41985),
            .I(N__41717));
    InMux I__8901 (
            .O(N__41984),
            .I(N__41712));
    InMux I__8900 (
            .O(N__41983),
            .I(N__41712));
    InMux I__8899 (
            .O(N__41982),
            .I(N__41709));
    InMux I__8898 (
            .O(N__41979),
            .I(N__41702));
    InMux I__8897 (
            .O(N__41976),
            .I(N__41702));
    InMux I__8896 (
            .O(N__41975),
            .I(N__41702));
    LocalMux I__8895 (
            .O(N__41972),
            .I(N__41689));
    LocalMux I__8894 (
            .O(N__41965),
            .I(N__41689));
    LocalMux I__8893 (
            .O(N__41958),
            .I(N__41689));
    LocalMux I__8892 (
            .O(N__41953),
            .I(N__41689));
    LocalMux I__8891 (
            .O(N__41944),
            .I(N__41689));
    LocalMux I__8890 (
            .O(N__41937),
            .I(N__41689));
    LocalMux I__8889 (
            .O(N__41932),
            .I(N__41684));
    LocalMux I__8888 (
            .O(N__41929),
            .I(N__41684));
    Span4Mux_h I__8887 (
            .O(N__41918),
            .I(N__41675));
    LocalMux I__8886 (
            .O(N__41911),
            .I(N__41675));
    LocalMux I__8885 (
            .O(N__41898),
            .I(N__41675));
    LocalMux I__8884 (
            .O(N__41893),
            .I(N__41675));
    InMux I__8883 (
            .O(N__41892),
            .I(N__41666));
    InMux I__8882 (
            .O(N__41891),
            .I(N__41666));
    InMux I__8881 (
            .O(N__41888),
            .I(N__41666));
    InMux I__8880 (
            .O(N__41887),
            .I(N__41666));
    InMux I__8879 (
            .O(N__41886),
            .I(N__41659));
    InMux I__8878 (
            .O(N__41885),
            .I(N__41659));
    InMux I__8877 (
            .O(N__41884),
            .I(N__41659));
    LocalMux I__8876 (
            .O(N__41879),
            .I(N__41652));
    LocalMux I__8875 (
            .O(N__41876),
            .I(N__41652));
    InMux I__8874 (
            .O(N__41875),
            .I(N__41643));
    InMux I__8873 (
            .O(N__41874),
            .I(N__41643));
    InMux I__8872 (
            .O(N__41873),
            .I(N__41643));
    InMux I__8871 (
            .O(N__41872),
            .I(N__41643));
    LocalMux I__8870 (
            .O(N__41869),
            .I(N__41640));
    InMux I__8869 (
            .O(N__41868),
            .I(N__41631));
    InMux I__8868 (
            .O(N__41867),
            .I(N__41631));
    InMux I__8867 (
            .O(N__41866),
            .I(N__41631));
    InMux I__8866 (
            .O(N__41865),
            .I(N__41631));
    InMux I__8865 (
            .O(N__41864),
            .I(N__41622));
    InMux I__8864 (
            .O(N__41863),
            .I(N__41622));
    InMux I__8863 (
            .O(N__41862),
            .I(N__41622));
    InMux I__8862 (
            .O(N__41861),
            .I(N__41622));
    Span4Mux_v I__8861 (
            .O(N__41856),
            .I(N__41615));
    LocalMux I__8860 (
            .O(N__41851),
            .I(N__41615));
    LocalMux I__8859 (
            .O(N__41842),
            .I(N__41615));
    InMux I__8858 (
            .O(N__41841),
            .I(N__41610));
    InMux I__8857 (
            .O(N__41838),
            .I(N__41610));
    LocalMux I__8856 (
            .O(N__41831),
            .I(N__41596));
    LocalMux I__8855 (
            .O(N__41824),
            .I(N__41596));
    Span4Mux_v I__8854 (
            .O(N__41821),
            .I(N__41596));
    LocalMux I__8853 (
            .O(N__41814),
            .I(N__41596));
    InMux I__8852 (
            .O(N__41813),
            .I(N__41587));
    InMux I__8851 (
            .O(N__41812),
            .I(N__41587));
    InMux I__8850 (
            .O(N__41811),
            .I(N__41587));
    InMux I__8849 (
            .O(N__41810),
            .I(N__41587));
    InMux I__8848 (
            .O(N__41809),
            .I(N__41582));
    InMux I__8847 (
            .O(N__41808),
            .I(N__41582));
    InMux I__8846 (
            .O(N__41807),
            .I(N__41579));
    InMux I__8845 (
            .O(N__41806),
            .I(N__41572));
    InMux I__8844 (
            .O(N__41805),
            .I(N__41572));
    InMux I__8843 (
            .O(N__41804),
            .I(N__41572));
    Span4Mux_v I__8842 (
            .O(N__41801),
            .I(N__41567));
    LocalMux I__8841 (
            .O(N__41792),
            .I(N__41567));
    LocalMux I__8840 (
            .O(N__41785),
            .I(N__41560));
    Span4Mux_v I__8839 (
            .O(N__41780),
            .I(N__41557));
    Span4Mux_h I__8838 (
            .O(N__41777),
            .I(N__41548));
    LocalMux I__8837 (
            .O(N__41768),
            .I(N__41548));
    LocalMux I__8836 (
            .O(N__41763),
            .I(N__41548));
    LocalMux I__8835 (
            .O(N__41756),
            .I(N__41548));
    LocalMux I__8834 (
            .O(N__41749),
            .I(N__41541));
    LocalMux I__8833 (
            .O(N__41744),
            .I(N__41541));
    LocalMux I__8832 (
            .O(N__41735),
            .I(N__41541));
    LocalMux I__8831 (
            .O(N__41730),
            .I(N__41538));
    LocalMux I__8830 (
            .O(N__41723),
            .I(N__41533));
    InMux I__8829 (
            .O(N__41722),
            .I(N__41526));
    InMux I__8828 (
            .O(N__41721),
            .I(N__41526));
    InMux I__8827 (
            .O(N__41720),
            .I(N__41526));
    LocalMux I__8826 (
            .O(N__41717),
            .I(N__41523));
    LocalMux I__8825 (
            .O(N__41712),
            .I(N__41506));
    LocalMux I__8824 (
            .O(N__41709),
            .I(N__41506));
    LocalMux I__8823 (
            .O(N__41702),
            .I(N__41506));
    Span4Mux_v I__8822 (
            .O(N__41689),
            .I(N__41506));
    Span4Mux_h I__8821 (
            .O(N__41684),
            .I(N__41506));
    Span4Mux_v I__8820 (
            .O(N__41675),
            .I(N__41506));
    LocalMux I__8819 (
            .O(N__41666),
            .I(N__41506));
    LocalMux I__8818 (
            .O(N__41659),
            .I(N__41506));
    InMux I__8817 (
            .O(N__41658),
            .I(N__41501));
    InMux I__8816 (
            .O(N__41657),
            .I(N__41501));
    Span4Mux_h I__8815 (
            .O(N__41652),
            .I(N__41494));
    LocalMux I__8814 (
            .O(N__41643),
            .I(N__41494));
    Span4Mux_v I__8813 (
            .O(N__41640),
            .I(N__41494));
    LocalMux I__8812 (
            .O(N__41631),
            .I(N__41489));
    LocalMux I__8811 (
            .O(N__41622),
            .I(N__41489));
    Span4Mux_h I__8810 (
            .O(N__41615),
            .I(N__41484));
    LocalMux I__8809 (
            .O(N__41610),
            .I(N__41484));
    InMux I__8808 (
            .O(N__41609),
            .I(N__41479));
    InMux I__8807 (
            .O(N__41608),
            .I(N__41479));
    InMux I__8806 (
            .O(N__41607),
            .I(N__41476));
    InMux I__8805 (
            .O(N__41606),
            .I(N__41471));
    InMux I__8804 (
            .O(N__41605),
            .I(N__41471));
    Sp12to4 I__8803 (
            .O(N__41596),
            .I(N__41464));
    LocalMux I__8802 (
            .O(N__41587),
            .I(N__41464));
    LocalMux I__8801 (
            .O(N__41582),
            .I(N__41464));
    LocalMux I__8800 (
            .O(N__41579),
            .I(N__41457));
    LocalMux I__8799 (
            .O(N__41572),
            .I(N__41457));
    Span4Mux_v I__8798 (
            .O(N__41567),
            .I(N__41457));
    InMux I__8797 (
            .O(N__41566),
            .I(N__41448));
    InMux I__8796 (
            .O(N__41565),
            .I(N__41448));
    InMux I__8795 (
            .O(N__41564),
            .I(N__41448));
    InMux I__8794 (
            .O(N__41563),
            .I(N__41448));
    Span4Mux_v I__8793 (
            .O(N__41560),
            .I(N__41441));
    Span4Mux_h I__8792 (
            .O(N__41557),
            .I(N__41441));
    Span4Mux_v I__8791 (
            .O(N__41548),
            .I(N__41441));
    Span12Mux_h I__8790 (
            .O(N__41541),
            .I(N__41436));
    Span12Mux_h I__8789 (
            .O(N__41538),
            .I(N__41436));
    InMux I__8788 (
            .O(N__41537),
            .I(N__41431));
    InMux I__8787 (
            .O(N__41536),
            .I(N__41431));
    Span4Mux_h I__8786 (
            .O(N__41533),
            .I(N__41424));
    LocalMux I__8785 (
            .O(N__41526),
            .I(N__41424));
    Span4Mux_v I__8784 (
            .O(N__41523),
            .I(N__41424));
    Span4Mux_v I__8783 (
            .O(N__41506),
            .I(N__41419));
    LocalMux I__8782 (
            .O(N__41501),
            .I(N__41419));
    Span4Mux_v I__8781 (
            .O(N__41494),
            .I(N__41412));
    Span4Mux_v I__8780 (
            .O(N__41489),
            .I(N__41412));
    Span4Mux_h I__8779 (
            .O(N__41484),
            .I(N__41412));
    LocalMux I__8778 (
            .O(N__41479),
            .I(sDAC_mem_pointerZ0Z_0));
    LocalMux I__8777 (
            .O(N__41476),
            .I(sDAC_mem_pointerZ0Z_0));
    LocalMux I__8776 (
            .O(N__41471),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv12 I__8775 (
            .O(N__41464),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv4 I__8774 (
            .O(N__41457),
            .I(sDAC_mem_pointerZ0Z_0));
    LocalMux I__8773 (
            .O(N__41448),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv4 I__8772 (
            .O(N__41441),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv12 I__8771 (
            .O(N__41436),
            .I(sDAC_mem_pointerZ0Z_0));
    LocalMux I__8770 (
            .O(N__41431),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv4 I__8769 (
            .O(N__41424),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv4 I__8768 (
            .O(N__41419),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv4 I__8767 (
            .O(N__41412),
            .I(sDAC_mem_pointerZ0Z_0));
    InMux I__8766 (
            .O(N__41387),
            .I(N__41384));
    LocalMux I__8765 (
            .O(N__41384),
            .I(N__41381));
    Odrv4 I__8764 (
            .O(N__41381),
            .I(sDAC_mem_37Z0Z_2));
    CascadeMux I__8763 (
            .O(N__41378),
            .I(sDAC_data_2_13_am_1_5_cascade_));
    InMux I__8762 (
            .O(N__41375),
            .I(N__41372));
    LocalMux I__8761 (
            .O(N__41372),
            .I(sDAC_data_RNO_4Z0Z_5));
    InMux I__8760 (
            .O(N__41369),
            .I(N__41366));
    LocalMux I__8759 (
            .O(N__41366),
            .I(N__41363));
    Span4Mux_h I__8758 (
            .O(N__41363),
            .I(N__41360));
    Odrv4 I__8757 (
            .O(N__41360),
            .I(sDAC_mem_25Z0Z_5));
    InMux I__8756 (
            .O(N__41357),
            .I(N__41354));
    LocalMux I__8755 (
            .O(N__41354),
            .I(N__41351));
    Span4Mux_h I__8754 (
            .O(N__41351),
            .I(N__41348));
    Odrv4 I__8753 (
            .O(N__41348),
            .I(sDAC_mem_25Z0Z_2));
    InMux I__8752 (
            .O(N__41345),
            .I(N__41342));
    LocalMux I__8751 (
            .O(N__41342),
            .I(sDAC_mem_25Z0Z_3));
    InMux I__8750 (
            .O(N__41339),
            .I(N__41336));
    LocalMux I__8749 (
            .O(N__41336),
            .I(N__41333));
    Span4Mux_h I__8748 (
            .O(N__41333),
            .I(N__41330));
    Span4Mux_h I__8747 (
            .O(N__41330),
            .I(N__41327));
    Odrv4 I__8746 (
            .O(N__41327),
            .I(sDAC_mem_25Z0Z_4));
    InMux I__8745 (
            .O(N__41324),
            .I(N__41321));
    LocalMux I__8744 (
            .O(N__41321),
            .I(N__41318));
    Span4Mux_h I__8743 (
            .O(N__41318),
            .I(N__41315));
    Odrv4 I__8742 (
            .O(N__41315),
            .I(sDAC_mem_25Z0Z_0));
    InMux I__8741 (
            .O(N__41312),
            .I(N__41309));
    LocalMux I__8740 (
            .O(N__41309),
            .I(N__41306));
    Span4Mux_h I__8739 (
            .O(N__41306),
            .I(N__41303));
    Span4Mux_h I__8738 (
            .O(N__41303),
            .I(N__41300));
    Odrv4 I__8737 (
            .O(N__41300),
            .I(sDAC_mem_25Z0Z_6));
    InMux I__8736 (
            .O(N__41297),
            .I(N__41294));
    LocalMux I__8735 (
            .O(N__41294),
            .I(sDAC_mem_32Z0Z_1));
    CascadeMux I__8734 (
            .O(N__41291),
            .I(sDAC_data_RNO_26Z0Z_5_cascade_));
    InMux I__8733 (
            .O(N__41288),
            .I(N__41285));
    LocalMux I__8732 (
            .O(N__41285),
            .I(sDAC_data_RNO_14Z0Z_5));
    InMux I__8731 (
            .O(N__41282),
            .I(N__41279));
    LocalMux I__8730 (
            .O(N__41279),
            .I(sDAC_mem_32Z0Z_2));
    CEMux I__8729 (
            .O(N__41276),
            .I(N__41272));
    CEMux I__8728 (
            .O(N__41275),
            .I(N__41269));
    LocalMux I__8727 (
            .O(N__41272),
            .I(N__41266));
    LocalMux I__8726 (
            .O(N__41269),
            .I(N__41262));
    Span4Mux_h I__8725 (
            .O(N__41266),
            .I(N__41259));
    CEMux I__8724 (
            .O(N__41265),
            .I(N__41255));
    Span4Mux_h I__8723 (
            .O(N__41262),
            .I(N__41252));
    Span4Mux_v I__8722 (
            .O(N__41259),
            .I(N__41249));
    CEMux I__8721 (
            .O(N__41258),
            .I(N__41246));
    LocalMux I__8720 (
            .O(N__41255),
            .I(N__41243));
    Span4Mux_h I__8719 (
            .O(N__41252),
            .I(N__41240));
    Span4Mux_h I__8718 (
            .O(N__41249),
            .I(N__41237));
    LocalMux I__8717 (
            .O(N__41246),
            .I(N__41234));
    Span4Mux_v I__8716 (
            .O(N__41243),
            .I(N__41231));
    Span4Mux_h I__8715 (
            .O(N__41240),
            .I(N__41226));
    Span4Mux_h I__8714 (
            .O(N__41237),
            .I(N__41226));
    Span12Mux_h I__8713 (
            .O(N__41234),
            .I(N__41223));
    Span4Mux_h I__8712 (
            .O(N__41231),
            .I(N__41220));
    Odrv4 I__8711 (
            .O(N__41226),
            .I(sDAC_mem_32_1_sqmuxa));
    Odrv12 I__8710 (
            .O(N__41223),
            .I(sDAC_mem_32_1_sqmuxa));
    Odrv4 I__8709 (
            .O(N__41220),
            .I(sDAC_mem_32_1_sqmuxa));
    InMux I__8708 (
            .O(N__41213),
            .I(N__41210));
    LocalMux I__8707 (
            .O(N__41210),
            .I(N__41207));
    Span12Mux_h I__8706 (
            .O(N__41207),
            .I(N__41204));
    Odrv12 I__8705 (
            .O(N__41204),
            .I(sDAC_mem_36Z0Z_0));
    InMux I__8704 (
            .O(N__41201),
            .I(N__41198));
    LocalMux I__8703 (
            .O(N__41198),
            .I(N__41195));
    Odrv4 I__8702 (
            .O(N__41195),
            .I(sDAC_mem_37Z0Z_0));
    CascadeMux I__8701 (
            .O(N__41192),
            .I(sDAC_data_2_13_am_1_3_cascade_));
    CascadeMux I__8700 (
            .O(N__41189),
            .I(N__41186));
    InMux I__8699 (
            .O(N__41186),
            .I(N__41183));
    LocalMux I__8698 (
            .O(N__41183),
            .I(N__41180));
    Odrv4 I__8697 (
            .O(N__41180),
            .I(sDAC_data_RNO_4Z0Z_3));
    InMux I__8696 (
            .O(N__41177),
            .I(N__41174));
    LocalMux I__8695 (
            .O(N__41174),
            .I(sDAC_mem_4Z0Z_0));
    InMux I__8694 (
            .O(N__41171),
            .I(N__41168));
    LocalMux I__8693 (
            .O(N__41168),
            .I(N__41165));
    Span4Mux_v I__8692 (
            .O(N__41165),
            .I(N__41162));
    Span4Mux_v I__8691 (
            .O(N__41162),
            .I(N__41159));
    Odrv4 I__8690 (
            .O(N__41159),
            .I(sDAC_mem_36Z0Z_1));
    CascadeMux I__8689 (
            .O(N__41156),
            .I(sDAC_data_2_13_am_1_4_cascade_));
    InMux I__8688 (
            .O(N__41153),
            .I(N__41150));
    LocalMux I__8687 (
            .O(N__41150),
            .I(N__41147));
    Odrv4 I__8686 (
            .O(N__41147),
            .I(sDAC_mem_37Z0Z_1));
    InMux I__8685 (
            .O(N__41144),
            .I(N__41141));
    LocalMux I__8684 (
            .O(N__41141),
            .I(N__41138));
    Span4Mux_v I__8683 (
            .O(N__41138),
            .I(N__41135));
    Odrv4 I__8682 (
            .O(N__41135),
            .I(sDAC_data_RNO_4Z0Z_4));
    InMux I__8681 (
            .O(N__41132),
            .I(N__41129));
    LocalMux I__8680 (
            .O(N__41129),
            .I(N__41126));
    Odrv12 I__8679 (
            .O(N__41126),
            .I(sDAC_mem_37Z0Z_3));
    InMux I__8678 (
            .O(N__41123),
            .I(N__41120));
    LocalMux I__8677 (
            .O(N__41120),
            .I(N__41117));
    Span4Mux_h I__8676 (
            .O(N__41117),
            .I(N__41114));
    Odrv4 I__8675 (
            .O(N__41114),
            .I(sDAC_mem_37Z0Z_4));
    InMux I__8674 (
            .O(N__41111),
            .I(N__41108));
    LocalMux I__8673 (
            .O(N__41108),
            .I(N__41105));
    Span4Mux_h I__8672 (
            .O(N__41105),
            .I(N__41102));
    Odrv4 I__8671 (
            .O(N__41102),
            .I(sDAC_mem_37Z0Z_5));
    InMux I__8670 (
            .O(N__41099),
            .I(N__41096));
    LocalMux I__8669 (
            .O(N__41096),
            .I(N__41093));
    Span4Mux_v I__8668 (
            .O(N__41093),
            .I(N__41090));
    Odrv4 I__8667 (
            .O(N__41090),
            .I(sDAC_mem_37Z0Z_6));
    InMux I__8666 (
            .O(N__41087),
            .I(N__41084));
    LocalMux I__8665 (
            .O(N__41084),
            .I(N__41081));
    Span4Mux_h I__8664 (
            .O(N__41081),
            .I(N__41078));
    Odrv4 I__8663 (
            .O(N__41078),
            .I(sDAC_mem_37Z0Z_7));
    CEMux I__8662 (
            .O(N__41075),
            .I(N__41072));
    LocalMux I__8661 (
            .O(N__41072),
            .I(N__41069));
    Span4Mux_h I__8660 (
            .O(N__41069),
            .I(N__41066));
    Span4Mux_h I__8659 (
            .O(N__41066),
            .I(N__41063));
    Odrv4 I__8658 (
            .O(N__41063),
            .I(sDAC_mem_37_1_sqmuxa));
    InMux I__8657 (
            .O(N__41060),
            .I(N__41057));
    LocalMux I__8656 (
            .O(N__41057),
            .I(sDAC_data_RNO_26Z0Z_3));
    InMux I__8655 (
            .O(N__41054),
            .I(N__41051));
    LocalMux I__8654 (
            .O(N__41051),
            .I(sDAC_data_RNO_14Z0Z_3));
    CascadeMux I__8653 (
            .O(N__41048),
            .I(sDAC_data_RNO_26Z0Z_4_cascade_));
    InMux I__8652 (
            .O(N__41045),
            .I(N__41042));
    LocalMux I__8651 (
            .O(N__41042),
            .I(N__41039));
    Span4Mux_v I__8650 (
            .O(N__41039),
            .I(N__41036));
    Odrv4 I__8649 (
            .O(N__41036),
            .I(sDAC_data_RNO_14Z0Z_4));
    InMux I__8648 (
            .O(N__41033),
            .I(N__41030));
    LocalMux I__8647 (
            .O(N__41030),
            .I(sDAC_mem_32Z0Z_0));
    CascadeMux I__8646 (
            .O(N__41027),
            .I(N__41023));
    InMux I__8645 (
            .O(N__41026),
            .I(N__41018));
    InMux I__8644 (
            .O(N__41023),
            .I(N__41018));
    LocalMux I__8643 (
            .O(N__41018),
            .I(sAddress_RNI6VH7_6Z0Z_1));
    CascadeMux I__8642 (
            .O(N__41015),
            .I(sAddress_RNI6VH7_6Z0Z_1_cascade_));
    CascadeMux I__8641 (
            .O(N__41012),
            .I(N__41007));
    CascadeMux I__8640 (
            .O(N__41011),
            .I(N__41004));
    CascadeMux I__8639 (
            .O(N__41010),
            .I(N__41001));
    InMux I__8638 (
            .O(N__41007),
            .I(N__40991));
    InMux I__8637 (
            .O(N__41004),
            .I(N__40986));
    InMux I__8636 (
            .O(N__41001),
            .I(N__40986));
    CascadeMux I__8635 (
            .O(N__41000),
            .I(N__40982));
    CascadeMux I__8634 (
            .O(N__40999),
            .I(N__40979));
    CascadeMux I__8633 (
            .O(N__40998),
            .I(N__40973));
    CascadeMux I__8632 (
            .O(N__40997),
            .I(N__40970));
    CascadeMux I__8631 (
            .O(N__40996),
            .I(N__40965));
    CascadeMux I__8630 (
            .O(N__40995),
            .I(N__40962));
    CascadeMux I__8629 (
            .O(N__40994),
            .I(N__40957));
    LocalMux I__8628 (
            .O(N__40991),
            .I(N__40951));
    LocalMux I__8627 (
            .O(N__40986),
            .I(N__40951));
    InMux I__8626 (
            .O(N__40985),
            .I(N__40940));
    InMux I__8625 (
            .O(N__40982),
            .I(N__40940));
    InMux I__8624 (
            .O(N__40979),
            .I(N__40940));
    InMux I__8623 (
            .O(N__40978),
            .I(N__40940));
    CascadeMux I__8622 (
            .O(N__40977),
            .I(N__40937));
    CascadeMux I__8621 (
            .O(N__40976),
            .I(N__40934));
    InMux I__8620 (
            .O(N__40973),
            .I(N__40931));
    InMux I__8619 (
            .O(N__40970),
            .I(N__40922));
    InMux I__8618 (
            .O(N__40969),
            .I(N__40922));
    InMux I__8617 (
            .O(N__40968),
            .I(N__40922));
    InMux I__8616 (
            .O(N__40965),
            .I(N__40922));
    InMux I__8615 (
            .O(N__40962),
            .I(N__40915));
    InMux I__8614 (
            .O(N__40961),
            .I(N__40915));
    InMux I__8613 (
            .O(N__40960),
            .I(N__40915));
    InMux I__8612 (
            .O(N__40957),
            .I(N__40910));
    InMux I__8611 (
            .O(N__40956),
            .I(N__40910));
    Span4Mux_v I__8610 (
            .O(N__40951),
            .I(N__40907));
    InMux I__8609 (
            .O(N__40950),
            .I(N__40904));
    InMux I__8608 (
            .O(N__40949),
            .I(N__40901));
    LocalMux I__8607 (
            .O(N__40940),
            .I(N__40897));
    InMux I__8606 (
            .O(N__40937),
            .I(N__40889));
    InMux I__8605 (
            .O(N__40934),
            .I(N__40889));
    LocalMux I__8604 (
            .O(N__40931),
            .I(N__40882));
    LocalMux I__8603 (
            .O(N__40922),
            .I(N__40882));
    LocalMux I__8602 (
            .O(N__40915),
            .I(N__40882));
    LocalMux I__8601 (
            .O(N__40910),
            .I(N__40877));
    Span4Mux_v I__8600 (
            .O(N__40907),
            .I(N__40877));
    LocalMux I__8599 (
            .O(N__40904),
            .I(N__40872));
    LocalMux I__8598 (
            .O(N__40901),
            .I(N__40872));
    CascadeMux I__8597 (
            .O(N__40900),
            .I(N__40868));
    Span4Mux_v I__8596 (
            .O(N__40897),
            .I(N__40865));
    InMux I__8595 (
            .O(N__40896),
            .I(N__40854));
    InMux I__8594 (
            .O(N__40895),
            .I(N__40854));
    InMux I__8593 (
            .O(N__40894),
            .I(N__40854));
    LocalMux I__8592 (
            .O(N__40889),
            .I(N__40851));
    Span4Mux_v I__8591 (
            .O(N__40882),
            .I(N__40844));
    Span4Mux_h I__8590 (
            .O(N__40877),
            .I(N__40844));
    Span4Mux_v I__8589 (
            .O(N__40872),
            .I(N__40844));
    InMux I__8588 (
            .O(N__40871),
            .I(N__40839));
    InMux I__8587 (
            .O(N__40868),
            .I(N__40839));
    Sp12to4 I__8586 (
            .O(N__40865),
            .I(N__40836));
    InMux I__8585 (
            .O(N__40864),
            .I(N__40829));
    InMux I__8584 (
            .O(N__40863),
            .I(N__40829));
    InMux I__8583 (
            .O(N__40862),
            .I(N__40829));
    InMux I__8582 (
            .O(N__40861),
            .I(N__40826));
    LocalMux I__8581 (
            .O(N__40854),
            .I(sAddressZ0Z_5));
    Odrv4 I__8580 (
            .O(N__40851),
            .I(sAddressZ0Z_5));
    Odrv4 I__8579 (
            .O(N__40844),
            .I(sAddressZ0Z_5));
    LocalMux I__8578 (
            .O(N__40839),
            .I(sAddressZ0Z_5));
    Odrv12 I__8577 (
            .O(N__40836),
            .I(sAddressZ0Z_5));
    LocalMux I__8576 (
            .O(N__40829),
            .I(sAddressZ0Z_5));
    LocalMux I__8575 (
            .O(N__40826),
            .I(sAddressZ0Z_5));
    InMux I__8574 (
            .O(N__40811),
            .I(N__40806));
    InMux I__8573 (
            .O(N__40810),
            .I(N__40801));
    InMux I__8572 (
            .O(N__40809),
            .I(N__40801));
    LocalMux I__8571 (
            .O(N__40806),
            .I(N__40790));
    LocalMux I__8570 (
            .O(N__40801),
            .I(N__40787));
    InMux I__8569 (
            .O(N__40800),
            .I(N__40775));
    InMux I__8568 (
            .O(N__40799),
            .I(N__40775));
    InMux I__8567 (
            .O(N__40798),
            .I(N__40775));
    InMux I__8566 (
            .O(N__40797),
            .I(N__40775));
    InMux I__8565 (
            .O(N__40796),
            .I(N__40766));
    InMux I__8564 (
            .O(N__40795),
            .I(N__40766));
    InMux I__8563 (
            .O(N__40794),
            .I(N__40766));
    InMux I__8562 (
            .O(N__40793),
            .I(N__40766));
    Span4Mux_v I__8561 (
            .O(N__40790),
            .I(N__40761));
    Span4Mux_v I__8560 (
            .O(N__40787),
            .I(N__40761));
    InMux I__8559 (
            .O(N__40786),
            .I(N__40754));
    InMux I__8558 (
            .O(N__40785),
            .I(N__40754));
    InMux I__8557 (
            .O(N__40784),
            .I(N__40754));
    LocalMux I__8556 (
            .O(N__40775),
            .I(N__40748));
    LocalMux I__8555 (
            .O(N__40766),
            .I(N__40733));
    Span4Mux_h I__8554 (
            .O(N__40761),
            .I(N__40733));
    LocalMux I__8553 (
            .O(N__40754),
            .I(N__40733));
    InMux I__8552 (
            .O(N__40753),
            .I(N__40726));
    InMux I__8551 (
            .O(N__40752),
            .I(N__40726));
    InMux I__8550 (
            .O(N__40751),
            .I(N__40726));
    Span4Mux_v I__8549 (
            .O(N__40748),
            .I(N__40723));
    InMux I__8548 (
            .O(N__40747),
            .I(N__40720));
    InMux I__8547 (
            .O(N__40746),
            .I(N__40715));
    InMux I__8546 (
            .O(N__40745),
            .I(N__40715));
    InMux I__8545 (
            .O(N__40744),
            .I(N__40708));
    InMux I__8544 (
            .O(N__40743),
            .I(N__40708));
    InMux I__8543 (
            .O(N__40742),
            .I(N__40708));
    InMux I__8542 (
            .O(N__40741),
            .I(N__40705));
    InMux I__8541 (
            .O(N__40740),
            .I(N__40702));
    Span4Mux_v I__8540 (
            .O(N__40733),
            .I(N__40699));
    LocalMux I__8539 (
            .O(N__40726),
            .I(N__40696));
    Sp12to4 I__8538 (
            .O(N__40723),
            .I(N__40693));
    LocalMux I__8537 (
            .O(N__40720),
            .I(sAddress_RNIP2UK1Z0Z_4));
    LocalMux I__8536 (
            .O(N__40715),
            .I(sAddress_RNIP2UK1Z0Z_4));
    LocalMux I__8535 (
            .O(N__40708),
            .I(sAddress_RNIP2UK1Z0Z_4));
    LocalMux I__8534 (
            .O(N__40705),
            .I(sAddress_RNIP2UK1Z0Z_4));
    LocalMux I__8533 (
            .O(N__40702),
            .I(sAddress_RNIP2UK1Z0Z_4));
    Odrv4 I__8532 (
            .O(N__40699),
            .I(sAddress_RNIP2UK1Z0Z_4));
    Odrv4 I__8531 (
            .O(N__40696),
            .I(sAddress_RNIP2UK1Z0Z_4));
    Odrv12 I__8530 (
            .O(N__40693),
            .I(sAddress_RNIP2UK1Z0Z_4));
    CascadeMux I__8529 (
            .O(N__40676),
            .I(N__40670));
    InMux I__8528 (
            .O(N__40675),
            .I(N__40660));
    InMux I__8527 (
            .O(N__40674),
            .I(N__40660));
    InMux I__8526 (
            .O(N__40673),
            .I(N__40660));
    InMux I__8525 (
            .O(N__40670),
            .I(N__40660));
    CascadeMux I__8524 (
            .O(N__40669),
            .I(N__40655));
    LocalMux I__8523 (
            .O(N__40660),
            .I(N__40648));
    InMux I__8522 (
            .O(N__40659),
            .I(N__40642));
    InMux I__8521 (
            .O(N__40658),
            .I(N__40633));
    InMux I__8520 (
            .O(N__40655),
            .I(N__40633));
    InMux I__8519 (
            .O(N__40654),
            .I(N__40633));
    InMux I__8518 (
            .O(N__40653),
            .I(N__40633));
    InMux I__8517 (
            .O(N__40652),
            .I(N__40627));
    InMux I__8516 (
            .O(N__40651),
            .I(N__40627));
    Span4Mux_v I__8515 (
            .O(N__40648),
            .I(N__40624));
    InMux I__8514 (
            .O(N__40647),
            .I(N__40621));
    InMux I__8513 (
            .O(N__40646),
            .I(N__40610));
    InMux I__8512 (
            .O(N__40645),
            .I(N__40610));
    LocalMux I__8511 (
            .O(N__40642),
            .I(N__40605));
    LocalMux I__8510 (
            .O(N__40633),
            .I(N__40605));
    InMux I__8509 (
            .O(N__40632),
            .I(N__40600));
    LocalMux I__8508 (
            .O(N__40627),
            .I(N__40597));
    Span4Mux_h I__8507 (
            .O(N__40624),
            .I(N__40592));
    LocalMux I__8506 (
            .O(N__40621),
            .I(N__40592));
    InMux I__8505 (
            .O(N__40620),
            .I(N__40589));
    InMux I__8504 (
            .O(N__40619),
            .I(N__40580));
    InMux I__8503 (
            .O(N__40618),
            .I(N__40580));
    InMux I__8502 (
            .O(N__40617),
            .I(N__40580));
    InMux I__8501 (
            .O(N__40616),
            .I(N__40580));
    InMux I__8500 (
            .O(N__40615),
            .I(N__40577));
    LocalMux I__8499 (
            .O(N__40610),
            .I(N__40572));
    Span12Mux_h I__8498 (
            .O(N__40605),
            .I(N__40572));
    InMux I__8497 (
            .O(N__40604),
            .I(N__40567));
    InMux I__8496 (
            .O(N__40603),
            .I(N__40567));
    LocalMux I__8495 (
            .O(N__40600),
            .I(N__40562));
    Sp12to4 I__8494 (
            .O(N__40597),
            .I(N__40562));
    Odrv4 I__8493 (
            .O(N__40592),
            .I(sAddressZ0Z_2));
    LocalMux I__8492 (
            .O(N__40589),
            .I(sAddressZ0Z_2));
    LocalMux I__8491 (
            .O(N__40580),
            .I(sAddressZ0Z_2));
    LocalMux I__8490 (
            .O(N__40577),
            .I(sAddressZ0Z_2));
    Odrv12 I__8489 (
            .O(N__40572),
            .I(sAddressZ0Z_2));
    LocalMux I__8488 (
            .O(N__40567),
            .I(sAddressZ0Z_2));
    Odrv12 I__8487 (
            .O(N__40562),
            .I(sAddressZ0Z_2));
    InMux I__8486 (
            .O(N__40547),
            .I(N__40540));
    InMux I__8485 (
            .O(N__40546),
            .I(N__40540));
    InMux I__8484 (
            .O(N__40545),
            .I(N__40537));
    LocalMux I__8483 (
            .O(N__40540),
            .I(N__40534));
    LocalMux I__8482 (
            .O(N__40537),
            .I(N__40528));
    Span4Mux_h I__8481 (
            .O(N__40534),
            .I(N__40525));
    InMux I__8480 (
            .O(N__40533),
            .I(N__40522));
    CascadeMux I__8479 (
            .O(N__40532),
            .I(N__40517));
    CascadeMux I__8478 (
            .O(N__40531),
            .I(N__40513));
    Span4Mux_h I__8477 (
            .O(N__40528),
            .I(N__40510));
    Span4Mux_h I__8476 (
            .O(N__40525),
            .I(N__40504));
    LocalMux I__8475 (
            .O(N__40522),
            .I(N__40501));
    CascadeMux I__8474 (
            .O(N__40521),
            .I(N__40497));
    InMux I__8473 (
            .O(N__40520),
            .I(N__40493));
    InMux I__8472 (
            .O(N__40517),
            .I(N__40488));
    InMux I__8471 (
            .O(N__40516),
            .I(N__40488));
    InMux I__8470 (
            .O(N__40513),
            .I(N__40485));
    Span4Mux_v I__8469 (
            .O(N__40510),
            .I(N__40482));
    InMux I__8468 (
            .O(N__40509),
            .I(N__40479));
    InMux I__8467 (
            .O(N__40508),
            .I(N__40474));
    InMux I__8466 (
            .O(N__40507),
            .I(N__40474));
    Span4Mux_h I__8465 (
            .O(N__40504),
            .I(N__40469));
    Span4Mux_h I__8464 (
            .O(N__40501),
            .I(N__40469));
    InMux I__8463 (
            .O(N__40500),
            .I(N__40466));
    InMux I__8462 (
            .O(N__40497),
            .I(N__40461));
    InMux I__8461 (
            .O(N__40496),
            .I(N__40461));
    LocalMux I__8460 (
            .O(N__40493),
            .I(N__40456));
    LocalMux I__8459 (
            .O(N__40488),
            .I(N__40456));
    LocalMux I__8458 (
            .O(N__40485),
            .I(sAddressZ0Z_1));
    Odrv4 I__8457 (
            .O(N__40482),
            .I(sAddressZ0Z_1));
    LocalMux I__8456 (
            .O(N__40479),
            .I(sAddressZ0Z_1));
    LocalMux I__8455 (
            .O(N__40474),
            .I(sAddressZ0Z_1));
    Odrv4 I__8454 (
            .O(N__40469),
            .I(sAddressZ0Z_1));
    LocalMux I__8453 (
            .O(N__40466),
            .I(sAddressZ0Z_1));
    LocalMux I__8452 (
            .O(N__40461),
            .I(sAddressZ0Z_1));
    Odrv12 I__8451 (
            .O(N__40456),
            .I(sAddressZ0Z_1));
    CascadeMux I__8450 (
            .O(N__40439),
            .I(N__40434));
    CascadeMux I__8449 (
            .O(N__40438),
            .I(N__40430));
    InMux I__8448 (
            .O(N__40437),
            .I(N__40419));
    InMux I__8447 (
            .O(N__40434),
            .I(N__40419));
    InMux I__8446 (
            .O(N__40433),
            .I(N__40419));
    InMux I__8445 (
            .O(N__40430),
            .I(N__40419));
    CascadeMux I__8444 (
            .O(N__40429),
            .I(N__40413));
    InMux I__8443 (
            .O(N__40428),
            .I(N__40399));
    LocalMux I__8442 (
            .O(N__40419),
            .I(N__40396));
    InMux I__8441 (
            .O(N__40418),
            .I(N__40391));
    InMux I__8440 (
            .O(N__40417),
            .I(N__40391));
    InMux I__8439 (
            .O(N__40416),
            .I(N__40386));
    InMux I__8438 (
            .O(N__40413),
            .I(N__40386));
    CascadeMux I__8437 (
            .O(N__40412),
            .I(N__40381));
    CascadeMux I__8436 (
            .O(N__40411),
            .I(N__40378));
    InMux I__8435 (
            .O(N__40410),
            .I(N__40374));
    InMux I__8434 (
            .O(N__40409),
            .I(N__40367));
    InMux I__8433 (
            .O(N__40408),
            .I(N__40367));
    InMux I__8432 (
            .O(N__40407),
            .I(N__40367));
    InMux I__8431 (
            .O(N__40406),
            .I(N__40364));
    InMux I__8430 (
            .O(N__40405),
            .I(N__40357));
    InMux I__8429 (
            .O(N__40404),
            .I(N__40357));
    InMux I__8428 (
            .O(N__40403),
            .I(N__40357));
    InMux I__8427 (
            .O(N__40402),
            .I(N__40354));
    LocalMux I__8426 (
            .O(N__40399),
            .I(N__40351));
    Span4Mux_v I__8425 (
            .O(N__40396),
            .I(N__40348));
    LocalMux I__8424 (
            .O(N__40391),
            .I(N__40343));
    LocalMux I__8423 (
            .O(N__40386),
            .I(N__40343));
    InMux I__8422 (
            .O(N__40385),
            .I(N__40340));
    InMux I__8421 (
            .O(N__40384),
            .I(N__40337));
    InMux I__8420 (
            .O(N__40381),
            .I(N__40329));
    InMux I__8419 (
            .O(N__40378),
            .I(N__40329));
    CascadeMux I__8418 (
            .O(N__40377),
            .I(N__40326));
    LocalMux I__8417 (
            .O(N__40374),
            .I(N__40315));
    LocalMux I__8416 (
            .O(N__40367),
            .I(N__40315));
    LocalMux I__8415 (
            .O(N__40364),
            .I(N__40315));
    LocalMux I__8414 (
            .O(N__40357),
            .I(N__40315));
    LocalMux I__8413 (
            .O(N__40354),
            .I(N__40315));
    Span4Mux_v I__8412 (
            .O(N__40351),
            .I(N__40308));
    Span4Mux_v I__8411 (
            .O(N__40348),
            .I(N__40308));
    Span4Mux_h I__8410 (
            .O(N__40343),
            .I(N__40308));
    LocalMux I__8409 (
            .O(N__40340),
            .I(N__40289));
    LocalMux I__8408 (
            .O(N__40337),
            .I(N__40289));
    InMux I__8407 (
            .O(N__40336),
            .I(N__40286));
    InMux I__8406 (
            .O(N__40335),
            .I(N__40281));
    InMux I__8405 (
            .O(N__40334),
            .I(N__40281));
    LocalMux I__8404 (
            .O(N__40329),
            .I(N__40278));
    InMux I__8403 (
            .O(N__40326),
            .I(N__40275));
    Span4Mux_v I__8402 (
            .O(N__40315),
            .I(N__40270));
    Span4Mux_h I__8401 (
            .O(N__40308),
            .I(N__40270));
    InMux I__8400 (
            .O(N__40307),
            .I(N__40264));
    InMux I__8399 (
            .O(N__40306),
            .I(N__40264));
    InMux I__8398 (
            .O(N__40305),
            .I(N__40255));
    InMux I__8397 (
            .O(N__40304),
            .I(N__40255));
    InMux I__8396 (
            .O(N__40303),
            .I(N__40255));
    InMux I__8395 (
            .O(N__40302),
            .I(N__40255));
    InMux I__8394 (
            .O(N__40301),
            .I(N__40252));
    InMux I__8393 (
            .O(N__40300),
            .I(N__40241));
    InMux I__8392 (
            .O(N__40299),
            .I(N__40241));
    InMux I__8391 (
            .O(N__40298),
            .I(N__40241));
    InMux I__8390 (
            .O(N__40297),
            .I(N__40241));
    InMux I__8389 (
            .O(N__40296),
            .I(N__40241));
    InMux I__8388 (
            .O(N__40295),
            .I(N__40236));
    InMux I__8387 (
            .O(N__40294),
            .I(N__40236));
    Span4Mux_v I__8386 (
            .O(N__40289),
            .I(N__40233));
    LocalMux I__8385 (
            .O(N__40286),
            .I(N__40224));
    LocalMux I__8384 (
            .O(N__40281),
            .I(N__40224));
    Span4Mux_v I__8383 (
            .O(N__40278),
            .I(N__40224));
    LocalMux I__8382 (
            .O(N__40275),
            .I(N__40224));
    Span4Mux_h I__8381 (
            .O(N__40270),
            .I(N__40221));
    InMux I__8380 (
            .O(N__40269),
            .I(N__40218));
    LocalMux I__8379 (
            .O(N__40264),
            .I(sAddressZ0Z_3));
    LocalMux I__8378 (
            .O(N__40255),
            .I(sAddressZ0Z_3));
    LocalMux I__8377 (
            .O(N__40252),
            .I(sAddressZ0Z_3));
    LocalMux I__8376 (
            .O(N__40241),
            .I(sAddressZ0Z_3));
    LocalMux I__8375 (
            .O(N__40236),
            .I(sAddressZ0Z_3));
    Odrv4 I__8374 (
            .O(N__40233),
            .I(sAddressZ0Z_3));
    Odrv4 I__8373 (
            .O(N__40224),
            .I(sAddressZ0Z_3));
    Odrv4 I__8372 (
            .O(N__40221),
            .I(sAddressZ0Z_3));
    LocalMux I__8371 (
            .O(N__40218),
            .I(sAddressZ0Z_3));
    CascadeMux I__8370 (
            .O(N__40199),
            .I(N__40192));
    CascadeMux I__8369 (
            .O(N__40198),
            .I(N__40186));
    InMux I__8368 (
            .O(N__40197),
            .I(N__40181));
    InMux I__8367 (
            .O(N__40196),
            .I(N__40181));
    CascadeMux I__8366 (
            .O(N__40195),
            .I(N__40177));
    InMux I__8365 (
            .O(N__40192),
            .I(N__40164));
    InMux I__8364 (
            .O(N__40191),
            .I(N__40164));
    InMux I__8363 (
            .O(N__40190),
            .I(N__40164));
    InMux I__8362 (
            .O(N__40189),
            .I(N__40164));
    InMux I__8361 (
            .O(N__40186),
            .I(N__40164));
    LocalMux I__8360 (
            .O(N__40181),
            .I(N__40154));
    InMux I__8359 (
            .O(N__40180),
            .I(N__40151));
    InMux I__8358 (
            .O(N__40177),
            .I(N__40148));
    InMux I__8357 (
            .O(N__40176),
            .I(N__40143));
    InMux I__8356 (
            .O(N__40175),
            .I(N__40143));
    LocalMux I__8355 (
            .O(N__40164),
            .I(N__40140));
    InMux I__8354 (
            .O(N__40163),
            .I(N__40134));
    InMux I__8353 (
            .O(N__40162),
            .I(N__40134));
    InMux I__8352 (
            .O(N__40161),
            .I(N__40129));
    InMux I__8351 (
            .O(N__40160),
            .I(N__40129));
    InMux I__8350 (
            .O(N__40159),
            .I(N__40124));
    InMux I__8349 (
            .O(N__40158),
            .I(N__40124));
    CascadeMux I__8348 (
            .O(N__40157),
            .I(N__40121));
    Span4Mux_v I__8347 (
            .O(N__40154),
            .I(N__40117));
    LocalMux I__8346 (
            .O(N__40151),
            .I(N__40110));
    LocalMux I__8345 (
            .O(N__40148),
            .I(N__40110));
    LocalMux I__8344 (
            .O(N__40143),
            .I(N__40110));
    Span4Mux_v I__8343 (
            .O(N__40140),
            .I(N__40107));
    InMux I__8342 (
            .O(N__40139),
            .I(N__40104));
    LocalMux I__8341 (
            .O(N__40134),
            .I(N__40097));
    LocalMux I__8340 (
            .O(N__40129),
            .I(N__40097));
    LocalMux I__8339 (
            .O(N__40124),
            .I(N__40097));
    InMux I__8338 (
            .O(N__40121),
            .I(N__40092));
    InMux I__8337 (
            .O(N__40120),
            .I(N__40092));
    Sp12to4 I__8336 (
            .O(N__40117),
            .I(N__40089));
    Span4Mux_v I__8335 (
            .O(N__40110),
            .I(N__40084));
    Span4Mux_v I__8334 (
            .O(N__40107),
            .I(N__40084));
    LocalMux I__8333 (
            .O(N__40104),
            .I(sAddressZ0Z_0));
    Odrv12 I__8332 (
            .O(N__40097),
            .I(sAddressZ0Z_0));
    LocalMux I__8331 (
            .O(N__40092),
            .I(sAddressZ0Z_0));
    Odrv12 I__8330 (
            .O(N__40089),
            .I(sAddressZ0Z_0));
    Odrv4 I__8329 (
            .O(N__40084),
            .I(sAddressZ0Z_0));
    InMux I__8328 (
            .O(N__40073),
            .I(N__40069));
    InMux I__8327 (
            .O(N__40072),
            .I(N__40066));
    LocalMux I__8326 (
            .O(N__40069),
            .I(N__40063));
    LocalMux I__8325 (
            .O(N__40066),
            .I(N__40060));
    Span4Mux_v I__8324 (
            .O(N__40063),
            .I(N__40057));
    Span4Mux_h I__8323 (
            .O(N__40060),
            .I(N__40054));
    Span4Mux_h I__8322 (
            .O(N__40057),
            .I(N__40049));
    Span4Mux_v I__8321 (
            .O(N__40054),
            .I(N__40046));
    InMux I__8320 (
            .O(N__40053),
            .I(N__40041));
    InMux I__8319 (
            .O(N__40052),
            .I(N__40041));
    Span4Mux_h I__8318 (
            .O(N__40049),
            .I(N__40034));
    Span4Mux_v I__8317 (
            .O(N__40046),
            .I(N__40034));
    LocalMux I__8316 (
            .O(N__40041),
            .I(N__40034));
    Odrv4 I__8315 (
            .O(N__40034),
            .I(sAddress_RNIAM2A_1Z0Z_1));
    CascadeMux I__8314 (
            .O(N__40031),
            .I(sAddress_RNIAM2A_1Z0Z_1_cascade_));
    InMux I__8313 (
            .O(N__40028),
            .I(N__40021));
    InMux I__8312 (
            .O(N__40027),
            .I(N__40016));
    InMux I__8311 (
            .O(N__40026),
            .I(N__40016));
    InMux I__8310 (
            .O(N__40025),
            .I(N__40011));
    InMux I__8309 (
            .O(N__40024),
            .I(N__40011));
    LocalMux I__8308 (
            .O(N__40021),
            .I(N__40006));
    LocalMux I__8307 (
            .O(N__40016),
            .I(N__40003));
    LocalMux I__8306 (
            .O(N__40011),
            .I(N__39999));
    InMux I__8305 (
            .O(N__40010),
            .I(N__39992));
    InMux I__8304 (
            .O(N__40009),
            .I(N__39992));
    Span4Mux_v I__8303 (
            .O(N__40006),
            .I(N__39988));
    Span4Mux_v I__8302 (
            .O(N__40003),
            .I(N__39985));
    InMux I__8301 (
            .O(N__40002),
            .I(N__39982));
    Span4Mux_v I__8300 (
            .O(N__39999),
            .I(N__39979));
    InMux I__8299 (
            .O(N__39998),
            .I(N__39974));
    InMux I__8298 (
            .O(N__39997),
            .I(N__39974));
    LocalMux I__8297 (
            .O(N__39992),
            .I(N__39966));
    InMux I__8296 (
            .O(N__39991),
            .I(N__39963));
    Sp12to4 I__8295 (
            .O(N__39988),
            .I(N__39958));
    Sp12to4 I__8294 (
            .O(N__39985),
            .I(N__39958));
    LocalMux I__8293 (
            .O(N__39982),
            .I(N__39951));
    Span4Mux_h I__8292 (
            .O(N__39979),
            .I(N__39951));
    LocalMux I__8291 (
            .O(N__39974),
            .I(N__39951));
    InMux I__8290 (
            .O(N__39973),
            .I(N__39948));
    InMux I__8289 (
            .O(N__39972),
            .I(N__39945));
    InMux I__8288 (
            .O(N__39971),
            .I(N__39940));
    InMux I__8287 (
            .O(N__39970),
            .I(N__39940));
    InMux I__8286 (
            .O(N__39969),
            .I(N__39937));
    Odrv4 I__8285 (
            .O(N__39966),
            .I(sAddress_RNIVREN1Z0Z_4));
    LocalMux I__8284 (
            .O(N__39963),
            .I(sAddress_RNIVREN1Z0Z_4));
    Odrv12 I__8283 (
            .O(N__39958),
            .I(sAddress_RNIVREN1Z0Z_4));
    Odrv4 I__8282 (
            .O(N__39951),
            .I(sAddress_RNIVREN1Z0Z_4));
    LocalMux I__8281 (
            .O(N__39948),
            .I(sAddress_RNIVREN1Z0Z_4));
    LocalMux I__8280 (
            .O(N__39945),
            .I(sAddress_RNIVREN1Z0Z_4));
    LocalMux I__8279 (
            .O(N__39940),
            .I(sAddress_RNIVREN1Z0Z_4));
    LocalMux I__8278 (
            .O(N__39937),
            .I(sAddress_RNIVREN1Z0Z_4));
    CEMux I__8277 (
            .O(N__39920),
            .I(N__39917));
    LocalMux I__8276 (
            .O(N__39917),
            .I(N__39914));
    Sp12to4 I__8275 (
            .O(N__39914),
            .I(N__39911));
    Odrv12 I__8274 (
            .O(N__39911),
            .I(sDAC_mem_17_1_sqmuxa));
    InMux I__8273 (
            .O(N__39908),
            .I(N__39905));
    LocalMux I__8272 (
            .O(N__39905),
            .I(N__39902));
    Span4Mux_v I__8271 (
            .O(N__39902),
            .I(N__39899));
    Odrv4 I__8270 (
            .O(N__39899),
            .I(sDAC_mem_41Z0Z_0));
    InMux I__8269 (
            .O(N__39896),
            .I(N__39893));
    LocalMux I__8268 (
            .O(N__39893),
            .I(N__39890));
    Span12Mux_v I__8267 (
            .O(N__39890),
            .I(N__39887));
    Odrv12 I__8266 (
            .O(N__39887),
            .I(sDAC_mem_41Z0Z_1));
    InMux I__8265 (
            .O(N__39884),
            .I(N__39881));
    LocalMux I__8264 (
            .O(N__39881),
            .I(N__39878));
    Span4Mux_v I__8263 (
            .O(N__39878),
            .I(N__39875));
    Odrv4 I__8262 (
            .O(N__39875),
            .I(sDAC_mem_41Z0Z_2));
    InMux I__8261 (
            .O(N__39872),
            .I(N__39869));
    LocalMux I__8260 (
            .O(N__39869),
            .I(N__39866));
    Span4Mux_v I__8259 (
            .O(N__39866),
            .I(N__39863));
    Span4Mux_h I__8258 (
            .O(N__39863),
            .I(N__39860));
    Odrv4 I__8257 (
            .O(N__39860),
            .I(sDAC_mem_41Z0Z_3));
    InMux I__8256 (
            .O(N__39857),
            .I(N__39854));
    LocalMux I__8255 (
            .O(N__39854),
            .I(N__39851));
    Span4Mux_h I__8254 (
            .O(N__39851),
            .I(N__39848));
    Span4Mux_h I__8253 (
            .O(N__39848),
            .I(N__39845));
    Odrv4 I__8252 (
            .O(N__39845),
            .I(sDAC_mem_41Z0Z_5));
    InMux I__8251 (
            .O(N__39842),
            .I(N__39839));
    LocalMux I__8250 (
            .O(N__39839),
            .I(N__39836));
    Span4Mux_h I__8249 (
            .O(N__39836),
            .I(N__39833));
    Odrv4 I__8248 (
            .O(N__39833),
            .I(sDAC_mem_41Z0Z_6));
    InMux I__8247 (
            .O(N__39830),
            .I(N__39827));
    LocalMux I__8246 (
            .O(N__39827),
            .I(N__39824));
    Span4Mux_v I__8245 (
            .O(N__39824),
            .I(N__39821));
    Odrv4 I__8244 (
            .O(N__39821),
            .I(sDAC_mem_41Z0Z_7));
    CEMux I__8243 (
            .O(N__39818),
            .I(N__39815));
    LocalMux I__8242 (
            .O(N__39815),
            .I(N__39812));
    Span4Mux_v I__8241 (
            .O(N__39812),
            .I(N__39809));
    Odrv4 I__8240 (
            .O(N__39809),
            .I(sDAC_mem_9_1_sqmuxa));
    CEMux I__8239 (
            .O(N__39806),
            .I(N__39803));
    LocalMux I__8238 (
            .O(N__39803),
            .I(N__39799));
    CEMux I__8237 (
            .O(N__39802),
            .I(N__39796));
    Span4Mux_v I__8236 (
            .O(N__39799),
            .I(N__39791));
    LocalMux I__8235 (
            .O(N__39796),
            .I(N__39791));
    Span4Mux_v I__8234 (
            .O(N__39791),
            .I(N__39788));
    Odrv4 I__8233 (
            .O(N__39788),
            .I(sDAC_mem_41_1_sqmuxa));
    IoInMux I__8232 (
            .O(N__39785),
            .I(N__39782));
    LocalMux I__8231 (
            .O(N__39782),
            .I(N__39779));
    IoSpan4Mux I__8230 (
            .O(N__39779),
            .I(N__39776));
    Span4Mux_s3_v I__8229 (
            .O(N__39776),
            .I(N__39773));
    Span4Mux_h I__8228 (
            .O(N__39773),
            .I(N__39769));
    CascadeMux I__8227 (
            .O(N__39772),
            .I(N__39766));
    Span4Mux_v I__8226 (
            .O(N__39769),
            .I(N__39763));
    InMux I__8225 (
            .O(N__39766),
            .I(N__39760));
    Odrv4 I__8224 (
            .O(N__39763),
            .I(RAM_DATA_cl_8Z0Z_15));
    LocalMux I__8223 (
            .O(N__39760),
            .I(RAM_DATA_cl_8Z0Z_15));
    IoInMux I__8222 (
            .O(N__39755),
            .I(N__39752));
    LocalMux I__8221 (
            .O(N__39752),
            .I(N__39749));
    Span4Mux_s3_v I__8220 (
            .O(N__39749),
            .I(N__39746));
    Span4Mux_h I__8219 (
            .O(N__39746),
            .I(N__39743));
    Span4Mux_h I__8218 (
            .O(N__39743),
            .I(N__39739));
    CascadeMux I__8217 (
            .O(N__39742),
            .I(N__39736));
    Span4Mux_v I__8216 (
            .O(N__39739),
            .I(N__39733));
    InMux I__8215 (
            .O(N__39736),
            .I(N__39730));
    Odrv4 I__8214 (
            .O(N__39733),
            .I(RAM_DATA_cl_9Z0Z_15));
    LocalMux I__8213 (
            .O(N__39730),
            .I(RAM_DATA_cl_9Z0Z_15));
    IoInMux I__8212 (
            .O(N__39725),
            .I(N__39722));
    LocalMux I__8211 (
            .O(N__39722),
            .I(N__39719));
    Span4Mux_s3_v I__8210 (
            .O(N__39719),
            .I(N__39716));
    Span4Mux_h I__8209 (
            .O(N__39716),
            .I(N__39713));
    Span4Mux_v I__8208 (
            .O(N__39713),
            .I(N__39709));
    InMux I__8207 (
            .O(N__39712),
            .I(N__39706));
    Odrv4 I__8206 (
            .O(N__39709),
            .I(RAM_DATA_clZ0Z_15));
    LocalMux I__8205 (
            .O(N__39706),
            .I(RAM_DATA_clZ0Z_15));
    IoInMux I__8204 (
            .O(N__39701),
            .I(N__39698));
    LocalMux I__8203 (
            .O(N__39698),
            .I(N__39695));
    IoSpan4Mux I__8202 (
            .O(N__39695),
            .I(N__39692));
    IoSpan4Mux I__8201 (
            .O(N__39692),
            .I(N__39689));
    IoSpan4Mux I__8200 (
            .O(N__39689),
            .I(N__39686));
    Span4Mux_s3_v I__8199 (
            .O(N__39686),
            .I(N__39683));
    Odrv4 I__8198 (
            .O(N__39683),
            .I(RAM_DATA_1Z0Z_7));
    InMux I__8197 (
            .O(N__39680),
            .I(N__39677));
    LocalMux I__8196 (
            .O(N__39677),
            .I(N__39674));
    Span4Mux_h I__8195 (
            .O(N__39674),
            .I(N__39671));
    Odrv4 I__8194 (
            .O(N__39671),
            .I(sDAC_mem_41Z0Z_4));
    InMux I__8193 (
            .O(N__39668),
            .I(N__39665));
    LocalMux I__8192 (
            .O(N__39665),
            .I(N__39662));
    Span4Mux_v I__8191 (
            .O(N__39662),
            .I(N__39659));
    Odrv4 I__8190 (
            .O(N__39659),
            .I(sDAC_mem_36Z0Z_3));
    InMux I__8189 (
            .O(N__39656),
            .I(N__39653));
    LocalMux I__8188 (
            .O(N__39653),
            .I(N__39650));
    Span4Mux_h I__8187 (
            .O(N__39650),
            .I(N__39647));
    Odrv4 I__8186 (
            .O(N__39647),
            .I(sDAC_mem_4Z0Z_3));
    CascadeMux I__8185 (
            .O(N__39644),
            .I(sDAC_data_2_13_am_1_6_cascade_));
    InMux I__8184 (
            .O(N__39641),
            .I(N__39638));
    LocalMux I__8183 (
            .O(N__39638),
            .I(N__39635));
    Odrv12 I__8182 (
            .O(N__39635),
            .I(sDAC_data_RNO_4Z0Z_6));
    InMux I__8181 (
            .O(N__39632),
            .I(N__39629));
    LocalMux I__8180 (
            .O(N__39629),
            .I(N__39626));
    Odrv4 I__8179 (
            .O(N__39626),
            .I(sDAC_mem_32Z0Z_5));
    InMux I__8178 (
            .O(N__39623),
            .I(N__39620));
    LocalMux I__8177 (
            .O(N__39620),
            .I(N__39617));
    Span4Mux_h I__8176 (
            .O(N__39617),
            .I(N__39614));
    Span4Mux_v I__8175 (
            .O(N__39614),
            .I(N__39611));
    Odrv4 I__8174 (
            .O(N__39611),
            .I(sDAC_mem_32Z0Z_7));
    CascadeMux I__8173 (
            .O(N__39608),
            .I(N__39605));
    InMux I__8172 (
            .O(N__39605),
            .I(N__39602));
    LocalMux I__8171 (
            .O(N__39602),
            .I(N__39598));
    InMux I__8170 (
            .O(N__39601),
            .I(N__39595));
    Span4Mux_h I__8169 (
            .O(N__39598),
            .I(N__39592));
    LocalMux I__8168 (
            .O(N__39595),
            .I(sCounterRAMZ0Z_2));
    Odrv4 I__8167 (
            .O(N__39592),
            .I(sCounterRAMZ0Z_2));
    InMux I__8166 (
            .O(N__39587),
            .I(sCounterRAM_cry_1));
    InMux I__8165 (
            .O(N__39584),
            .I(N__39580));
    InMux I__8164 (
            .O(N__39583),
            .I(N__39577));
    LocalMux I__8163 (
            .O(N__39580),
            .I(N__39574));
    LocalMux I__8162 (
            .O(N__39577),
            .I(sCounterRAMZ0Z_3));
    Odrv4 I__8161 (
            .O(N__39574),
            .I(sCounterRAMZ0Z_3));
    InMux I__8160 (
            .O(N__39569),
            .I(sCounterRAM_cry_2));
    InMux I__8159 (
            .O(N__39566),
            .I(N__39562));
    InMux I__8158 (
            .O(N__39565),
            .I(N__39559));
    LocalMux I__8157 (
            .O(N__39562),
            .I(N__39556));
    LocalMux I__8156 (
            .O(N__39559),
            .I(sCounterRAMZ0Z_4));
    Odrv4 I__8155 (
            .O(N__39556),
            .I(sCounterRAMZ0Z_4));
    InMux I__8154 (
            .O(N__39551),
            .I(sCounterRAM_cry_3));
    InMux I__8153 (
            .O(N__39548),
            .I(N__39544));
    InMux I__8152 (
            .O(N__39547),
            .I(N__39541));
    LocalMux I__8151 (
            .O(N__39544),
            .I(N__39538));
    LocalMux I__8150 (
            .O(N__39541),
            .I(sCounterRAMZ0Z_5));
    Odrv4 I__8149 (
            .O(N__39538),
            .I(sCounterRAMZ0Z_5));
    InMux I__8148 (
            .O(N__39533),
            .I(sCounterRAM_cry_4));
    InMux I__8147 (
            .O(N__39530),
            .I(N__39526));
    InMux I__8146 (
            .O(N__39529),
            .I(N__39523));
    LocalMux I__8145 (
            .O(N__39526),
            .I(N__39520));
    LocalMux I__8144 (
            .O(N__39523),
            .I(sCounterRAMZ0Z_6));
    Odrv4 I__8143 (
            .O(N__39520),
            .I(sCounterRAMZ0Z_6));
    InMux I__8142 (
            .O(N__39515),
            .I(sCounterRAM_cry_5));
    InMux I__8141 (
            .O(N__39512),
            .I(N__39496));
    InMux I__8140 (
            .O(N__39511),
            .I(N__39496));
    InMux I__8139 (
            .O(N__39510),
            .I(N__39496));
    InMux I__8138 (
            .O(N__39509),
            .I(N__39496));
    InMux I__8137 (
            .O(N__39508),
            .I(N__39487));
    InMux I__8136 (
            .O(N__39507),
            .I(N__39487));
    InMux I__8135 (
            .O(N__39506),
            .I(N__39487));
    InMux I__8134 (
            .O(N__39505),
            .I(N__39487));
    LocalMux I__8133 (
            .O(N__39496),
            .I(N_70_i));
    LocalMux I__8132 (
            .O(N__39487),
            .I(N_70_i));
    InMux I__8131 (
            .O(N__39482),
            .I(sCounterRAM_cry_6));
    CascadeMux I__8130 (
            .O(N__39479),
            .I(N__39476));
    InMux I__8129 (
            .O(N__39476),
            .I(N__39472));
    InMux I__8128 (
            .O(N__39475),
            .I(N__39469));
    LocalMux I__8127 (
            .O(N__39472),
            .I(N__39466));
    LocalMux I__8126 (
            .O(N__39469),
            .I(sCounterRAMZ0Z_7));
    Odrv4 I__8125 (
            .O(N__39466),
            .I(sCounterRAMZ0Z_7));
    IoInMux I__8124 (
            .O(N__39461),
            .I(N__39458));
    LocalMux I__8123 (
            .O(N__39458),
            .I(N__39455));
    IoSpan4Mux I__8122 (
            .O(N__39455),
            .I(N__39452));
    Span4Mux_s3_h I__8121 (
            .O(N__39452),
            .I(N__39449));
    Sp12to4 I__8120 (
            .O(N__39449),
            .I(N__39446));
    Span12Mux_v I__8119 (
            .O(N__39446),
            .I(N__39442));
    CascadeMux I__8118 (
            .O(N__39445),
            .I(N__39439));
    Span12Mux_v I__8117 (
            .O(N__39442),
            .I(N__39436));
    InMux I__8116 (
            .O(N__39439),
            .I(N__39433));
    Odrv12 I__8115 (
            .O(N__39436),
            .I(RAM_DATA_cl_6Z0Z_15));
    LocalMux I__8114 (
            .O(N__39433),
            .I(RAM_DATA_cl_6Z0Z_15));
    IoInMux I__8113 (
            .O(N__39428),
            .I(N__39425));
    LocalMux I__8112 (
            .O(N__39425),
            .I(N__39422));
    Span12Mux_s11_h I__8111 (
            .O(N__39422),
            .I(N__39418));
    InMux I__8110 (
            .O(N__39421),
            .I(N__39415));
    Odrv12 I__8109 (
            .O(N__39418),
            .I(RAM_DATA_cl_7Z0Z_15));
    LocalMux I__8108 (
            .O(N__39415),
            .I(RAM_DATA_cl_7Z0Z_15));
    InMux I__8107 (
            .O(N__39410),
            .I(N__39378));
    InMux I__8106 (
            .O(N__39409),
            .I(N__39378));
    InMux I__8105 (
            .O(N__39408),
            .I(N__39378));
    InMux I__8104 (
            .O(N__39407),
            .I(N__39378));
    InMux I__8103 (
            .O(N__39406),
            .I(N__39369));
    InMux I__8102 (
            .O(N__39405),
            .I(N__39369));
    InMux I__8101 (
            .O(N__39404),
            .I(N__39369));
    InMux I__8100 (
            .O(N__39403),
            .I(N__39369));
    InMux I__8099 (
            .O(N__39402),
            .I(N__39360));
    InMux I__8098 (
            .O(N__39401),
            .I(N__39360));
    InMux I__8097 (
            .O(N__39400),
            .I(N__39360));
    InMux I__8096 (
            .O(N__39399),
            .I(N__39360));
    InMux I__8095 (
            .O(N__39398),
            .I(N__39351));
    InMux I__8094 (
            .O(N__39397),
            .I(N__39351));
    InMux I__8093 (
            .O(N__39396),
            .I(N__39348));
    InMux I__8092 (
            .O(N__39395),
            .I(N__39331));
    InMux I__8091 (
            .O(N__39394),
            .I(N__39331));
    InMux I__8090 (
            .O(N__39393),
            .I(N__39331));
    InMux I__8089 (
            .O(N__39392),
            .I(N__39331));
    InMux I__8088 (
            .O(N__39391),
            .I(N__39322));
    InMux I__8087 (
            .O(N__39390),
            .I(N__39322));
    InMux I__8086 (
            .O(N__39389),
            .I(N__39322));
    InMux I__8085 (
            .O(N__39388),
            .I(N__39322));
    CascadeMux I__8084 (
            .O(N__39387),
            .I(N__39319));
    LocalMux I__8083 (
            .O(N__39378),
            .I(N__39312));
    LocalMux I__8082 (
            .O(N__39369),
            .I(N__39312));
    LocalMux I__8081 (
            .O(N__39360),
            .I(N__39312));
    InMux I__8080 (
            .O(N__39359),
            .I(N__39303));
    InMux I__8079 (
            .O(N__39358),
            .I(N__39303));
    InMux I__8078 (
            .O(N__39357),
            .I(N__39303));
    InMux I__8077 (
            .O(N__39356),
            .I(N__39303));
    LocalMux I__8076 (
            .O(N__39351),
            .I(N__39298));
    LocalMux I__8075 (
            .O(N__39348),
            .I(N__39298));
    InMux I__8074 (
            .O(N__39347),
            .I(N__39286));
    InMux I__8073 (
            .O(N__39346),
            .I(N__39286));
    InMux I__8072 (
            .O(N__39345),
            .I(N__39286));
    InMux I__8071 (
            .O(N__39344),
            .I(N__39286));
    InMux I__8070 (
            .O(N__39343),
            .I(N__39277));
    InMux I__8069 (
            .O(N__39342),
            .I(N__39277));
    InMux I__8068 (
            .O(N__39341),
            .I(N__39277));
    InMux I__8067 (
            .O(N__39340),
            .I(N__39277));
    LocalMux I__8066 (
            .O(N__39331),
            .I(N__39272));
    LocalMux I__8065 (
            .O(N__39322),
            .I(N__39272));
    InMux I__8064 (
            .O(N__39319),
            .I(N__39269));
    Span4Mux_v I__8063 (
            .O(N__39312),
            .I(N__39262));
    LocalMux I__8062 (
            .O(N__39303),
            .I(N__39262));
    Span4Mux_v I__8061 (
            .O(N__39298),
            .I(N__39262));
    InMux I__8060 (
            .O(N__39297),
            .I(N__39257));
    InMux I__8059 (
            .O(N__39296),
            .I(N__39257));
    InMux I__8058 (
            .O(N__39295),
            .I(N__39254));
    LocalMux I__8057 (
            .O(N__39286),
            .I(N__39249));
    LocalMux I__8056 (
            .O(N__39277),
            .I(N__39249));
    Span4Mux_h I__8055 (
            .O(N__39272),
            .I(N__39243));
    LocalMux I__8054 (
            .O(N__39269),
            .I(N__39243));
    Span4Mux_h I__8053 (
            .O(N__39262),
            .I(N__39240));
    LocalMux I__8052 (
            .O(N__39257),
            .I(N__39235));
    LocalMux I__8051 (
            .O(N__39254),
            .I(N__39235));
    Span4Mux_h I__8050 (
            .O(N__39249),
            .I(N__39232));
    InMux I__8049 (
            .O(N__39248),
            .I(N__39229));
    Span4Mux_v I__8048 (
            .O(N__39243),
            .I(N__39226));
    Sp12to4 I__8047 (
            .O(N__39240),
            .I(N__39220));
    Span12Mux_h I__8046 (
            .O(N__39235),
            .I(N__39220));
    Sp12to4 I__8045 (
            .O(N__39232),
            .I(N__39215));
    LocalMux I__8044 (
            .O(N__39229),
            .I(N__39215));
    Span4Mux_h I__8043 (
            .O(N__39226),
            .I(N__39212));
    InMux I__8042 (
            .O(N__39225),
            .I(N__39209));
    Span12Mux_v I__8041 (
            .O(N__39220),
            .I(N__39204));
    Span12Mux_v I__8040 (
            .O(N__39215),
            .I(N__39204));
    Span4Mux_v I__8039 (
            .O(N__39212),
            .I(N__39201));
    LocalMux I__8038 (
            .O(N__39209),
            .I(sEEPointerResetZ0));
    Odrv12 I__8037 (
            .O(N__39204),
            .I(sEEPointerResetZ0));
    Odrv4 I__8036 (
            .O(N__39201),
            .I(sEEPointerResetZ0));
    CascadeMux I__8035 (
            .O(N__39194),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3_cascade_));
    IoInMux I__8034 (
            .O(N__39191),
            .I(N__39188));
    LocalMux I__8033 (
            .O(N__39188),
            .I(N__39185));
    IoSpan4Mux I__8032 (
            .O(N__39185),
            .I(N__39182));
    Span4Mux_s2_v I__8031 (
            .O(N__39182),
            .I(N__39179));
    Span4Mux_v I__8030 (
            .O(N__39179),
            .I(N__39176));
    Odrv4 I__8029 (
            .O(N__39176),
            .I(N_28));
    CascadeMux I__8028 (
            .O(N__39173),
            .I(N__39169));
    CascadeMux I__8027 (
            .O(N__39172),
            .I(N__39166));
    InMux I__8026 (
            .O(N__39169),
            .I(N__39160));
    InMux I__8025 (
            .O(N__39166),
            .I(N__39155));
    InMux I__8024 (
            .O(N__39165),
            .I(N__39155));
    InMux I__8023 (
            .O(N__39164),
            .I(N__39150));
    InMux I__8022 (
            .O(N__39163),
            .I(N__39150));
    LocalMux I__8021 (
            .O(N__39160),
            .I(N__39145));
    LocalMux I__8020 (
            .O(N__39155),
            .I(N__39145));
    LocalMux I__8019 (
            .O(N__39150),
            .I(sSPI_MSB0LSBZ0Z1));
    Odrv12 I__8018 (
            .O(N__39145),
            .I(sSPI_MSB0LSBZ0Z1));
    InMux I__8017 (
            .O(N__39140),
            .I(N__39134));
    InMux I__8016 (
            .O(N__39139),
            .I(N__39134));
    LocalMux I__8015 (
            .O(N__39134),
            .I(N__39131));
    Span4Mux_v I__8014 (
            .O(N__39131),
            .I(N__39124));
    InMux I__8013 (
            .O(N__39130),
            .I(N__39115));
    InMux I__8012 (
            .O(N__39129),
            .I(N__39115));
    InMux I__8011 (
            .O(N__39128),
            .I(N__39115));
    InMux I__8010 (
            .O(N__39127),
            .I(N__39115));
    Span4Mux_v I__8009 (
            .O(N__39124),
            .I(N__39112));
    LocalMux I__8008 (
            .O(N__39115),
            .I(N__39109));
    Sp12to4 I__8007 (
            .O(N__39112),
            .I(N__39104));
    Span12Mux_v I__8006 (
            .O(N__39109),
            .I(N__39104));
    Odrv12 I__8005 (
            .O(N__39104),
            .I(spi_mosi_ready_prev3_RNILKERZ0));
    IoInMux I__8004 (
            .O(N__39101),
            .I(N__39098));
    LocalMux I__8003 (
            .O(N__39098),
            .I(N__39095));
    IoSpan4Mux I__8002 (
            .O(N__39095),
            .I(N__39092));
    IoSpan4Mux I__8001 (
            .O(N__39092),
            .I(N__39089));
    Span4Mux_s1_h I__8000 (
            .O(N__39089),
            .I(N__39086));
    Sp12to4 I__7999 (
            .O(N__39086),
            .I(N__39083));
    Span12Mux_v I__7998 (
            .O(N__39083),
            .I(N__39079));
    InMux I__7997 (
            .O(N__39082),
            .I(N__39076));
    Odrv12 I__7996 (
            .O(N__39079),
            .I(RAM_DATA_cl_11Z0Z_15));
    LocalMux I__7995 (
            .O(N__39076),
            .I(RAM_DATA_cl_11Z0Z_15));
    IoInMux I__7994 (
            .O(N__39071),
            .I(N__39068));
    LocalMux I__7993 (
            .O(N__39068),
            .I(N__39065));
    Span4Mux_s2_v I__7992 (
            .O(N__39065),
            .I(N__39062));
    Sp12to4 I__7991 (
            .O(N__39062),
            .I(N__39059));
    Span12Mux_s11_h I__7990 (
            .O(N__39059),
            .I(N__39055));
    InMux I__7989 (
            .O(N__39058),
            .I(N__39052));
    Odrv12 I__7988 (
            .O(N__39055),
            .I(RAM_DATA_cl_12Z0Z_15));
    LocalMux I__7987 (
            .O(N__39052),
            .I(RAM_DATA_cl_12Z0Z_15));
    InMux I__7986 (
            .O(N__39047),
            .I(N__39043));
    InMux I__7985 (
            .O(N__39046),
            .I(N__39040));
    LocalMux I__7984 (
            .O(N__39043),
            .I(N__39037));
    LocalMux I__7983 (
            .O(N__39040),
            .I(sCounterRAMZ0Z_0));
    Odrv4 I__7982 (
            .O(N__39037),
            .I(sCounterRAMZ0Z_0));
    InMux I__7981 (
            .O(N__39032),
            .I(bfn_17_18_0_));
    InMux I__7980 (
            .O(N__39029),
            .I(N__39026));
    LocalMux I__7979 (
            .O(N__39026),
            .I(N__39022));
    InMux I__7978 (
            .O(N__39025),
            .I(N__39019));
    Span4Mux_v I__7977 (
            .O(N__39022),
            .I(N__39016));
    LocalMux I__7976 (
            .O(N__39019),
            .I(sCounterRAMZ0Z_1));
    Odrv4 I__7975 (
            .O(N__39016),
            .I(sCounterRAMZ0Z_1));
    InMux I__7974 (
            .O(N__39011),
            .I(sCounterRAM_cry_0));
    InMux I__7973 (
            .O(N__39008),
            .I(N__39005));
    LocalMux I__7972 (
            .O(N__39005),
            .I(N__39002));
    Span4Mux_v I__7971 (
            .O(N__39002),
            .I(N__38999));
    Span4Mux_v I__7970 (
            .O(N__38999),
            .I(N__38996));
    Odrv4 I__7969 (
            .O(N__38996),
            .I(sDAC_mem_17Z0Z_4));
    InMux I__7968 (
            .O(N__38993),
            .I(N__38990));
    LocalMux I__7967 (
            .O(N__38990),
            .I(N__38987));
    Span4Mux_v I__7966 (
            .O(N__38987),
            .I(N__38984));
    Span4Mux_h I__7965 (
            .O(N__38984),
            .I(N__38981));
    Odrv4 I__7964 (
            .O(N__38981),
            .I(sDAC_mem_17Z0Z_5));
    InMux I__7963 (
            .O(N__38978),
            .I(N__38975));
    LocalMux I__7962 (
            .O(N__38975),
            .I(N__38972));
    Span4Mux_h I__7961 (
            .O(N__38972),
            .I(N__38969));
    Span4Mux_v I__7960 (
            .O(N__38969),
            .I(N__38966));
    Odrv4 I__7959 (
            .O(N__38966),
            .I(sDAC_mem_17Z0Z_6));
    InMux I__7958 (
            .O(N__38963),
            .I(N__38960));
    LocalMux I__7957 (
            .O(N__38960),
            .I(N__38957));
    Span4Mux_h I__7956 (
            .O(N__38957),
            .I(N__38954));
    Odrv4 I__7955 (
            .O(N__38954),
            .I(sDAC_mem_17Z0Z_7));
    InMux I__7954 (
            .O(N__38951),
            .I(N__38948));
    LocalMux I__7953 (
            .O(N__38948),
            .I(N__38945));
    Span4Mux_v I__7952 (
            .O(N__38945),
            .I(N__38942));
    Span4Mux_h I__7951 (
            .O(N__38942),
            .I(N__38939));
    Span4Mux_h I__7950 (
            .O(N__38939),
            .I(N__38936));
    Span4Mux_v I__7949 (
            .O(N__38936),
            .I(N__38933));
    Odrv4 I__7948 (
            .O(N__38933),
            .I(RAM_DATA_in_14));
    CascadeMux I__7947 (
            .O(N__38930),
            .I(N__38927));
    InMux I__7946 (
            .O(N__38927),
            .I(N__38924));
    LocalMux I__7945 (
            .O(N__38924),
            .I(N__38921));
    Span4Mux_v I__7944 (
            .O(N__38921),
            .I(N__38918));
    Sp12to4 I__7943 (
            .O(N__38918),
            .I(N__38915));
    Span12Mux_h I__7942 (
            .O(N__38915),
            .I(N__38912));
    Span12Mux_v I__7941 (
            .O(N__38912),
            .I(N__38909));
    Odrv12 I__7940 (
            .O(N__38909),
            .I(RAM_DATA_in_6));
    InMux I__7939 (
            .O(N__38906),
            .I(N__38902));
    InMux I__7938 (
            .O(N__38905),
            .I(N__38899));
    LocalMux I__7937 (
            .O(N__38902),
            .I(N__38896));
    LocalMux I__7936 (
            .O(N__38899),
            .I(button_debounce_counterZ0Z_13));
    Odrv4 I__7935 (
            .O(N__38896),
            .I(button_debounce_counterZ0Z_13));
    InMux I__7934 (
            .O(N__38891),
            .I(N__38887));
    InMux I__7933 (
            .O(N__38890),
            .I(N__38884));
    LocalMux I__7932 (
            .O(N__38887),
            .I(N__38881));
    LocalMux I__7931 (
            .O(N__38884),
            .I(button_debounce_counterZ0Z_12));
    Odrv4 I__7930 (
            .O(N__38881),
            .I(button_debounce_counterZ0Z_12));
    CascadeMux I__7929 (
            .O(N__38876),
            .I(N__38873));
    InMux I__7928 (
            .O(N__38873),
            .I(N__38869));
    InMux I__7927 (
            .O(N__38872),
            .I(N__38866));
    LocalMux I__7926 (
            .O(N__38869),
            .I(N__38863));
    LocalMux I__7925 (
            .O(N__38866),
            .I(button_debounce_counterZ0Z_14));
    Odrv4 I__7924 (
            .O(N__38863),
            .I(button_debounce_counterZ0Z_14));
    InMux I__7923 (
            .O(N__38858),
            .I(N__38854));
    InMux I__7922 (
            .O(N__38857),
            .I(N__38851));
    LocalMux I__7921 (
            .O(N__38854),
            .I(N__38848));
    LocalMux I__7920 (
            .O(N__38851),
            .I(button_debounce_counterZ0Z_11));
    Odrv4 I__7919 (
            .O(N__38848),
            .I(button_debounce_counterZ0Z_11));
    InMux I__7918 (
            .O(N__38843),
            .I(N__38840));
    LocalMux I__7917 (
            .O(N__38840),
            .I(N__38837));
    Odrv4 I__7916 (
            .O(N__38837),
            .I(sbuttonModeStatus_0_sqmuxa_15));
    InMux I__7915 (
            .O(N__38834),
            .I(N__38831));
    LocalMux I__7914 (
            .O(N__38831),
            .I(N__38827));
    InMux I__7913 (
            .O(N__38830),
            .I(N__38824));
    Span4Mux_h I__7912 (
            .O(N__38827),
            .I(N__38821));
    LocalMux I__7911 (
            .O(N__38824),
            .I(button_debounce_counterZ0Z_9));
    Odrv4 I__7910 (
            .O(N__38821),
            .I(button_debounce_counterZ0Z_9));
    InMux I__7909 (
            .O(N__38816),
            .I(N__38812));
    InMux I__7908 (
            .O(N__38815),
            .I(N__38809));
    LocalMux I__7907 (
            .O(N__38812),
            .I(N__38806));
    LocalMux I__7906 (
            .O(N__38809),
            .I(button_debounce_counterZ0Z_7));
    Odrv4 I__7905 (
            .O(N__38806),
            .I(button_debounce_counterZ0Z_7));
    CascadeMux I__7904 (
            .O(N__38801),
            .I(N__38798));
    InMux I__7903 (
            .O(N__38798),
            .I(N__38795));
    LocalMux I__7902 (
            .O(N__38795),
            .I(N__38791));
    InMux I__7901 (
            .O(N__38794),
            .I(N__38788));
    Span4Mux_v I__7900 (
            .O(N__38791),
            .I(N__38785));
    LocalMux I__7899 (
            .O(N__38788),
            .I(button_debounce_counterZ0Z_10));
    Odrv4 I__7898 (
            .O(N__38785),
            .I(button_debounce_counterZ0Z_10));
    InMux I__7897 (
            .O(N__38780),
            .I(N__38776));
    InMux I__7896 (
            .O(N__38779),
            .I(N__38773));
    LocalMux I__7895 (
            .O(N__38776),
            .I(N__38770));
    LocalMux I__7894 (
            .O(N__38773),
            .I(button_debounce_counterZ0Z_8));
    Odrv4 I__7893 (
            .O(N__38770),
            .I(button_debounce_counterZ0Z_8));
    InMux I__7892 (
            .O(N__38765),
            .I(N__38762));
    LocalMux I__7891 (
            .O(N__38762),
            .I(N__38759));
    Odrv12 I__7890 (
            .O(N__38759),
            .I(sbuttonModeStatus_0_sqmuxa_16));
    InMux I__7889 (
            .O(N__38756),
            .I(N__38753));
    LocalMux I__7888 (
            .O(N__38753),
            .I(N__38750));
    Span4Mux_v I__7887 (
            .O(N__38750),
            .I(N__38747));
    Sp12to4 I__7886 (
            .O(N__38747),
            .I(N__38744));
    Span12Mux_h I__7885 (
            .O(N__38744),
            .I(N__38741));
    Odrv12 I__7884 (
            .O(N__38741),
            .I(RAM_DATA_in_0));
    CascadeMux I__7883 (
            .O(N__38738),
            .I(N__38735));
    InMux I__7882 (
            .O(N__38735),
            .I(N__38732));
    LocalMux I__7881 (
            .O(N__38732),
            .I(N__38729));
    Span4Mux_v I__7880 (
            .O(N__38729),
            .I(N__38726));
    Span4Mux_h I__7879 (
            .O(N__38726),
            .I(N__38723));
    Sp12to4 I__7878 (
            .O(N__38723),
            .I(N__38720));
    Span12Mux_v I__7877 (
            .O(N__38720),
            .I(N__38717));
    Odrv12 I__7876 (
            .O(N__38717),
            .I(RAM_DATA_in_8));
    InMux I__7875 (
            .O(N__38714),
            .I(N__38711));
    LocalMux I__7874 (
            .O(N__38711),
            .I(N__38708));
    Span4Mux_v I__7873 (
            .O(N__38708),
            .I(N__38705));
    Span4Mux_h I__7872 (
            .O(N__38705),
            .I(N__38702));
    Span4Mux_h I__7871 (
            .O(N__38702),
            .I(N__38699));
    IoSpan4Mux I__7870 (
            .O(N__38699),
            .I(N__38696));
    Odrv4 I__7869 (
            .O(N__38696),
            .I(RAM_DATA_in_12));
    CascadeMux I__7868 (
            .O(N__38693),
            .I(N__38690));
    InMux I__7867 (
            .O(N__38690),
            .I(N__38687));
    LocalMux I__7866 (
            .O(N__38687),
            .I(N__38684));
    Span4Mux_v I__7865 (
            .O(N__38684),
            .I(N__38681));
    Sp12to4 I__7864 (
            .O(N__38681),
            .I(N__38678));
    Span12Mux_h I__7863 (
            .O(N__38678),
            .I(N__38675));
    Odrv12 I__7862 (
            .O(N__38675),
            .I(RAM_DATA_in_4));
    InMux I__7861 (
            .O(N__38672),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0 ));
    InMux I__7860 (
            .O(N__38669),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1 ));
    InMux I__7859 (
            .O(N__38666),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2 ));
    InMux I__7858 (
            .O(N__38663),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3 ));
    InMux I__7857 (
            .O(N__38660),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4 ));
    InMux I__7856 (
            .O(N__38657),
            .I(N__38654));
    LocalMux I__7855 (
            .O(N__38654),
            .I(N__38650));
    InMux I__7854 (
            .O(N__38653),
            .I(N__38647));
    Span4Mux_h I__7853 (
            .O(N__38650),
            .I(N__38644));
    LocalMux I__7852 (
            .O(N__38647),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5 ));
    Odrv4 I__7851 (
            .O(N__38644),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5 ));
    InMux I__7850 (
            .O(N__38639),
            .I(N__38636));
    LocalMux I__7849 (
            .O(N__38636),
            .I(N__38633));
    Odrv12 I__7848 (
            .O(N__38633),
            .I(sDAC_mem_17Z0Z_0));
    InMux I__7847 (
            .O(N__38630),
            .I(N__38627));
    LocalMux I__7846 (
            .O(N__38627),
            .I(N__38624));
    Odrv12 I__7845 (
            .O(N__38624),
            .I(sDAC_mem_17Z0Z_1));
    InMux I__7844 (
            .O(N__38621),
            .I(N__38618));
    LocalMux I__7843 (
            .O(N__38618),
            .I(N__38615));
    Odrv4 I__7842 (
            .O(N__38615),
            .I(sDAC_mem_17Z0Z_2));
    InMux I__7841 (
            .O(N__38612),
            .I(N__38609));
    LocalMux I__7840 (
            .O(N__38609),
            .I(N__38606));
    Span4Mux_h I__7839 (
            .O(N__38606),
            .I(N__38603));
    Span4Mux_v I__7838 (
            .O(N__38603),
            .I(N__38600));
    Odrv4 I__7837 (
            .O(N__38600),
            .I(sDAC_mem_17Z0Z_3));
    InMux I__7836 (
            .O(N__38597),
            .I(N__38594));
    LocalMux I__7835 (
            .O(N__38594),
            .I(N__38591));
    Span4Mux_h I__7834 (
            .O(N__38591),
            .I(N__38588));
    Span4Mux_h I__7833 (
            .O(N__38588),
            .I(N__38585));
    Span4Mux_h I__7832 (
            .O(N__38585),
            .I(N__38582));
    Odrv4 I__7831 (
            .O(N__38582),
            .I(sDAC_mem_29Z0Z_2));
    InMux I__7830 (
            .O(N__38579),
            .I(N__38576));
    LocalMux I__7829 (
            .O(N__38576),
            .I(sDAC_data_RNO_23Z0Z_5));
    InMux I__7828 (
            .O(N__38573),
            .I(N__38570));
    LocalMux I__7827 (
            .O(N__38570),
            .I(N__38567));
    Span4Mux_v I__7826 (
            .O(N__38567),
            .I(N__38564));
    Span4Mux_h I__7825 (
            .O(N__38564),
            .I(N__38561));
    Odrv4 I__7824 (
            .O(N__38561),
            .I(sDAC_mem_24Z0Z_3));
    InMux I__7823 (
            .O(N__38558),
            .I(N__38547));
    InMux I__7822 (
            .O(N__38557),
            .I(N__38542));
    InMux I__7821 (
            .O(N__38556),
            .I(N__38542));
    InMux I__7820 (
            .O(N__38555),
            .I(N__38539));
    InMux I__7819 (
            .O(N__38554),
            .I(N__38534));
    InMux I__7818 (
            .O(N__38553),
            .I(N__38534));
    CascadeMux I__7817 (
            .O(N__38552),
            .I(N__38527));
    InMux I__7816 (
            .O(N__38551),
            .I(N__38521));
    InMux I__7815 (
            .O(N__38550),
            .I(N__38521));
    LocalMux I__7814 (
            .O(N__38547),
            .I(N__38512));
    LocalMux I__7813 (
            .O(N__38542),
            .I(N__38512));
    LocalMux I__7812 (
            .O(N__38539),
            .I(N__38512));
    LocalMux I__7811 (
            .O(N__38534),
            .I(N__38512));
    InMux I__7810 (
            .O(N__38533),
            .I(N__38501));
    InMux I__7809 (
            .O(N__38532),
            .I(N__38501));
    CascadeMux I__7808 (
            .O(N__38531),
            .I(N__38497));
    InMux I__7807 (
            .O(N__38530),
            .I(N__38494));
    InMux I__7806 (
            .O(N__38527),
            .I(N__38491));
    InMux I__7805 (
            .O(N__38526),
            .I(N__38486));
    LocalMux I__7804 (
            .O(N__38521),
            .I(N__38481));
    Span4Mux_v I__7803 (
            .O(N__38512),
            .I(N__38481));
    InMux I__7802 (
            .O(N__38511),
            .I(N__38478));
    CascadeMux I__7801 (
            .O(N__38510),
            .I(N__38473));
    InMux I__7800 (
            .O(N__38509),
            .I(N__38470));
    InMux I__7799 (
            .O(N__38508),
            .I(N__38467));
    InMux I__7798 (
            .O(N__38507),
            .I(N__38464));
    InMux I__7797 (
            .O(N__38506),
            .I(N__38461));
    LocalMux I__7796 (
            .O(N__38501),
            .I(N__38456));
    InMux I__7795 (
            .O(N__38500),
            .I(N__38453));
    InMux I__7794 (
            .O(N__38497),
            .I(N__38449));
    LocalMux I__7793 (
            .O(N__38494),
            .I(N__38445));
    LocalMux I__7792 (
            .O(N__38491),
            .I(N__38442));
    InMux I__7791 (
            .O(N__38490),
            .I(N__38437));
    InMux I__7790 (
            .O(N__38489),
            .I(N__38437));
    LocalMux I__7789 (
            .O(N__38486),
            .I(N__38430));
    Span4Mux_v I__7788 (
            .O(N__38481),
            .I(N__38430));
    LocalMux I__7787 (
            .O(N__38478),
            .I(N__38430));
    InMux I__7786 (
            .O(N__38477),
            .I(N__38427));
    InMux I__7785 (
            .O(N__38476),
            .I(N__38420));
    InMux I__7784 (
            .O(N__38473),
            .I(N__38420));
    LocalMux I__7783 (
            .O(N__38470),
            .I(N__38415));
    LocalMux I__7782 (
            .O(N__38467),
            .I(N__38415));
    LocalMux I__7781 (
            .O(N__38464),
            .I(N__38409));
    LocalMux I__7780 (
            .O(N__38461),
            .I(N__38409));
    InMux I__7779 (
            .O(N__38460),
            .I(N__38404));
    InMux I__7778 (
            .O(N__38459),
            .I(N__38404));
    Span4Mux_v I__7777 (
            .O(N__38456),
            .I(N__38397));
    LocalMux I__7776 (
            .O(N__38453),
            .I(N__38397));
    InMux I__7775 (
            .O(N__38452),
            .I(N__38394));
    LocalMux I__7774 (
            .O(N__38449),
            .I(N__38391));
    InMux I__7773 (
            .O(N__38448),
            .I(N__38388));
    Span4Mux_v I__7772 (
            .O(N__38445),
            .I(N__38384));
    Span4Mux_h I__7771 (
            .O(N__38442),
            .I(N__38375));
    LocalMux I__7770 (
            .O(N__38437),
            .I(N__38375));
    Span4Mux_h I__7769 (
            .O(N__38430),
            .I(N__38375));
    LocalMux I__7768 (
            .O(N__38427),
            .I(N__38375));
    InMux I__7767 (
            .O(N__38426),
            .I(N__38372));
    InMux I__7766 (
            .O(N__38425),
            .I(N__38369));
    LocalMux I__7765 (
            .O(N__38420),
            .I(N__38364));
    Span4Mux_h I__7764 (
            .O(N__38415),
            .I(N__38364));
    InMux I__7763 (
            .O(N__38414),
            .I(N__38361));
    Span4Mux_v I__7762 (
            .O(N__38409),
            .I(N__38356));
    LocalMux I__7761 (
            .O(N__38404),
            .I(N__38356));
    InMux I__7760 (
            .O(N__38403),
            .I(N__38353));
    InMux I__7759 (
            .O(N__38402),
            .I(N__38350));
    Span4Mux_v I__7758 (
            .O(N__38397),
            .I(N__38347));
    LocalMux I__7757 (
            .O(N__38394),
            .I(N__38340));
    Span4Mux_v I__7756 (
            .O(N__38391),
            .I(N__38340));
    LocalMux I__7755 (
            .O(N__38388),
            .I(N__38340));
    InMux I__7754 (
            .O(N__38387),
            .I(N__38337));
    Span4Mux_h I__7753 (
            .O(N__38384),
            .I(N__38332));
    Span4Mux_v I__7752 (
            .O(N__38375),
            .I(N__38332));
    LocalMux I__7751 (
            .O(N__38372),
            .I(N__38321));
    LocalMux I__7750 (
            .O(N__38369),
            .I(N__38321));
    Span4Mux_v I__7749 (
            .O(N__38364),
            .I(N__38321));
    LocalMux I__7748 (
            .O(N__38361),
            .I(N__38321));
    Span4Mux_h I__7747 (
            .O(N__38356),
            .I(N__38321));
    LocalMux I__7746 (
            .O(N__38353),
            .I(sDAC_mem_pointerZ0Z_1));
    LocalMux I__7745 (
            .O(N__38350),
            .I(sDAC_mem_pointerZ0Z_1));
    Odrv4 I__7744 (
            .O(N__38347),
            .I(sDAC_mem_pointerZ0Z_1));
    Odrv4 I__7743 (
            .O(N__38340),
            .I(sDAC_mem_pointerZ0Z_1));
    LocalMux I__7742 (
            .O(N__38337),
            .I(sDAC_mem_pointerZ0Z_1));
    Odrv4 I__7741 (
            .O(N__38332),
            .I(sDAC_mem_pointerZ0Z_1));
    Odrv4 I__7740 (
            .O(N__38321),
            .I(sDAC_mem_pointerZ0Z_1));
    CascadeMux I__7739 (
            .O(N__38306),
            .I(sDAC_data_RNO_30Z0Z_6_cascade_));
    InMux I__7738 (
            .O(N__38303),
            .I(N__38297));
    InMux I__7737 (
            .O(N__38302),
            .I(N__38292));
    InMux I__7736 (
            .O(N__38301),
            .I(N__38292));
    InMux I__7735 (
            .O(N__38300),
            .I(N__38282));
    LocalMux I__7734 (
            .O(N__38297),
            .I(N__38277));
    LocalMux I__7733 (
            .O(N__38292),
            .I(N__38277));
    InMux I__7732 (
            .O(N__38291),
            .I(N__38272));
    InMux I__7731 (
            .O(N__38290),
            .I(N__38272));
    InMux I__7730 (
            .O(N__38289),
            .I(N__38263));
    InMux I__7729 (
            .O(N__38288),
            .I(N__38263));
    InMux I__7728 (
            .O(N__38287),
            .I(N__38263));
    InMux I__7727 (
            .O(N__38286),
            .I(N__38263));
    CascadeMux I__7726 (
            .O(N__38285),
            .I(N__38259));
    LocalMux I__7725 (
            .O(N__38282),
            .I(N__38246));
    Span4Mux_v I__7724 (
            .O(N__38277),
            .I(N__38239));
    LocalMux I__7723 (
            .O(N__38272),
            .I(N__38239));
    LocalMux I__7722 (
            .O(N__38263),
            .I(N__38239));
    InMux I__7721 (
            .O(N__38262),
            .I(N__38234));
    InMux I__7720 (
            .O(N__38259),
            .I(N__38234));
    CascadeMux I__7719 (
            .O(N__38258),
            .I(N__38227));
    CascadeMux I__7718 (
            .O(N__38257),
            .I(N__38224));
    CascadeMux I__7717 (
            .O(N__38256),
            .I(N__38221));
    CascadeMux I__7716 (
            .O(N__38255),
            .I(N__38218));
    CascadeMux I__7715 (
            .O(N__38254),
            .I(N__38213));
    CascadeMux I__7714 (
            .O(N__38253),
            .I(N__38204));
    InMux I__7713 (
            .O(N__38252),
            .I(N__38197));
    CascadeMux I__7712 (
            .O(N__38251),
            .I(N__38191));
    InMux I__7711 (
            .O(N__38250),
            .I(N__38185));
    InMux I__7710 (
            .O(N__38249),
            .I(N__38185));
    Span4Mux_h I__7709 (
            .O(N__38246),
            .I(N__38178));
    Span4Mux_v I__7708 (
            .O(N__38239),
            .I(N__38178));
    LocalMux I__7707 (
            .O(N__38234),
            .I(N__38178));
    CascadeMux I__7706 (
            .O(N__38233),
            .I(N__38174));
    CascadeMux I__7705 (
            .O(N__38232),
            .I(N__38171));
    InMux I__7704 (
            .O(N__38231),
            .I(N__38163));
    InMux I__7703 (
            .O(N__38230),
            .I(N__38156));
    InMux I__7702 (
            .O(N__38227),
            .I(N__38156));
    InMux I__7701 (
            .O(N__38224),
            .I(N__38156));
    InMux I__7700 (
            .O(N__38221),
            .I(N__38151));
    InMux I__7699 (
            .O(N__38218),
            .I(N__38151));
    InMux I__7698 (
            .O(N__38217),
            .I(N__38144));
    InMux I__7697 (
            .O(N__38216),
            .I(N__38144));
    InMux I__7696 (
            .O(N__38213),
            .I(N__38144));
    CascadeMux I__7695 (
            .O(N__38212),
            .I(N__38141));
    CascadeMux I__7694 (
            .O(N__38211),
            .I(N__38138));
    CascadeMux I__7693 (
            .O(N__38210),
            .I(N__38135));
    CascadeMux I__7692 (
            .O(N__38209),
            .I(N__38132));
    CascadeMux I__7691 (
            .O(N__38208),
            .I(N__38126));
    CascadeMux I__7690 (
            .O(N__38207),
            .I(N__38123));
    InMux I__7689 (
            .O(N__38204),
            .I(N__38118));
    CascadeMux I__7688 (
            .O(N__38203),
            .I(N__38112));
    InMux I__7687 (
            .O(N__38202),
            .I(N__38108));
    CascadeMux I__7686 (
            .O(N__38201),
            .I(N__38105));
    CascadeMux I__7685 (
            .O(N__38200),
            .I(N__38101));
    LocalMux I__7684 (
            .O(N__38197),
            .I(N__38098));
    CascadeMux I__7683 (
            .O(N__38196),
            .I(N__38092));
    CascadeMux I__7682 (
            .O(N__38195),
            .I(N__38088));
    InMux I__7681 (
            .O(N__38194),
            .I(N__38083));
    InMux I__7680 (
            .O(N__38191),
            .I(N__38083));
    InMux I__7679 (
            .O(N__38190),
            .I(N__38080));
    LocalMux I__7678 (
            .O(N__38185),
            .I(N__38075));
    Span4Mux_v I__7677 (
            .O(N__38178),
            .I(N__38075));
    InMux I__7676 (
            .O(N__38177),
            .I(N__38066));
    InMux I__7675 (
            .O(N__38174),
            .I(N__38066));
    InMux I__7674 (
            .O(N__38171),
            .I(N__38066));
    InMux I__7673 (
            .O(N__38170),
            .I(N__38066));
    InMux I__7672 (
            .O(N__38169),
            .I(N__38061));
    InMux I__7671 (
            .O(N__38168),
            .I(N__38061));
    InMux I__7670 (
            .O(N__38167),
            .I(N__38056));
    InMux I__7669 (
            .O(N__38166),
            .I(N__38056));
    LocalMux I__7668 (
            .O(N__38163),
            .I(N__38053));
    LocalMux I__7667 (
            .O(N__38156),
            .I(N__38048));
    LocalMux I__7666 (
            .O(N__38151),
            .I(N__38048));
    LocalMux I__7665 (
            .O(N__38144),
            .I(N__38045));
    InMux I__7664 (
            .O(N__38141),
            .I(N__38042));
    InMux I__7663 (
            .O(N__38138),
            .I(N__38035));
    InMux I__7662 (
            .O(N__38135),
            .I(N__38035));
    InMux I__7661 (
            .O(N__38132),
            .I(N__38035));
    InMux I__7660 (
            .O(N__38131),
            .I(N__38032));
    InMux I__7659 (
            .O(N__38130),
            .I(N__38025));
    InMux I__7658 (
            .O(N__38129),
            .I(N__38025));
    InMux I__7657 (
            .O(N__38126),
            .I(N__38020));
    InMux I__7656 (
            .O(N__38123),
            .I(N__38020));
    InMux I__7655 (
            .O(N__38122),
            .I(N__38015));
    InMux I__7654 (
            .O(N__38121),
            .I(N__38015));
    LocalMux I__7653 (
            .O(N__38118),
            .I(N__38012));
    InMux I__7652 (
            .O(N__38117),
            .I(N__38009));
    InMux I__7651 (
            .O(N__38116),
            .I(N__38002));
    InMux I__7650 (
            .O(N__38115),
            .I(N__38002));
    InMux I__7649 (
            .O(N__38112),
            .I(N__38002));
    InMux I__7648 (
            .O(N__38111),
            .I(N__37998));
    LocalMux I__7647 (
            .O(N__38108),
            .I(N__37994));
    InMux I__7646 (
            .O(N__38105),
            .I(N__37989));
    InMux I__7645 (
            .O(N__38104),
            .I(N__37989));
    InMux I__7644 (
            .O(N__38101),
            .I(N__37986));
    Span4Mux_v I__7643 (
            .O(N__38098),
            .I(N__37983));
    InMux I__7642 (
            .O(N__38097),
            .I(N__37980));
    InMux I__7641 (
            .O(N__38096),
            .I(N__37975));
    InMux I__7640 (
            .O(N__38095),
            .I(N__37975));
    InMux I__7639 (
            .O(N__38092),
            .I(N__37968));
    InMux I__7638 (
            .O(N__38091),
            .I(N__37968));
    InMux I__7637 (
            .O(N__38088),
            .I(N__37968));
    LocalMux I__7636 (
            .O(N__38083),
            .I(N__37959));
    LocalMux I__7635 (
            .O(N__38080),
            .I(N__37959));
    Span4Mux_h I__7634 (
            .O(N__38075),
            .I(N__37959));
    LocalMux I__7633 (
            .O(N__38066),
            .I(N__37959));
    LocalMux I__7632 (
            .O(N__38061),
            .I(N__37948));
    LocalMux I__7631 (
            .O(N__38056),
            .I(N__37948));
    Span4Mux_h I__7630 (
            .O(N__38053),
            .I(N__37948));
    Span4Mux_v I__7629 (
            .O(N__38048),
            .I(N__37948));
    Span4Mux_h I__7628 (
            .O(N__38045),
            .I(N__37948));
    LocalMux I__7627 (
            .O(N__38042),
            .I(N__37943));
    LocalMux I__7626 (
            .O(N__38035),
            .I(N__37943));
    LocalMux I__7625 (
            .O(N__38032),
            .I(N__37940));
    InMux I__7624 (
            .O(N__38031),
            .I(N__37937));
    InMux I__7623 (
            .O(N__38030),
            .I(N__37934));
    LocalMux I__7622 (
            .O(N__38025),
            .I(N__37929));
    LocalMux I__7621 (
            .O(N__38020),
            .I(N__37929));
    LocalMux I__7620 (
            .O(N__38015),
            .I(N__37926));
    Span4Mux_h I__7619 (
            .O(N__38012),
            .I(N__37919));
    LocalMux I__7618 (
            .O(N__38009),
            .I(N__37919));
    LocalMux I__7617 (
            .O(N__38002),
            .I(N__37919));
    InMux I__7616 (
            .O(N__38001),
            .I(N__37916));
    LocalMux I__7615 (
            .O(N__37998),
            .I(N__37913));
    InMux I__7614 (
            .O(N__37997),
            .I(N__37910));
    Span4Mux_v I__7613 (
            .O(N__37994),
            .I(N__37907));
    LocalMux I__7612 (
            .O(N__37989),
            .I(N__37902));
    LocalMux I__7611 (
            .O(N__37986),
            .I(N__37902));
    Span4Mux_h I__7610 (
            .O(N__37983),
            .I(N__37891));
    LocalMux I__7609 (
            .O(N__37980),
            .I(N__37891));
    LocalMux I__7608 (
            .O(N__37975),
            .I(N__37891));
    LocalMux I__7607 (
            .O(N__37968),
            .I(N__37891));
    Span4Mux_v I__7606 (
            .O(N__37959),
            .I(N__37891));
    Span4Mux_v I__7605 (
            .O(N__37948),
            .I(N__37886));
    Span4Mux_h I__7604 (
            .O(N__37943),
            .I(N__37886));
    Span12Mux_h I__7603 (
            .O(N__37940),
            .I(N__37873));
    LocalMux I__7602 (
            .O(N__37937),
            .I(N__37873));
    LocalMux I__7601 (
            .O(N__37934),
            .I(N__37873));
    Span12Mux_h I__7600 (
            .O(N__37929),
            .I(N__37873));
    Sp12to4 I__7599 (
            .O(N__37926),
            .I(N__37873));
    Sp12to4 I__7598 (
            .O(N__37919),
            .I(N__37873));
    LocalMux I__7597 (
            .O(N__37916),
            .I(sDAC_mem_pointerZ0Z_2));
    Odrv12 I__7596 (
            .O(N__37913),
            .I(sDAC_mem_pointerZ0Z_2));
    LocalMux I__7595 (
            .O(N__37910),
            .I(sDAC_mem_pointerZ0Z_2));
    Odrv4 I__7594 (
            .O(N__37907),
            .I(sDAC_mem_pointerZ0Z_2));
    Odrv4 I__7593 (
            .O(N__37902),
            .I(sDAC_mem_pointerZ0Z_2));
    Odrv4 I__7592 (
            .O(N__37891),
            .I(sDAC_mem_pointerZ0Z_2));
    Odrv4 I__7591 (
            .O(N__37886),
            .I(sDAC_mem_pointerZ0Z_2));
    Odrv12 I__7590 (
            .O(N__37873),
            .I(sDAC_mem_pointerZ0Z_2));
    InMux I__7589 (
            .O(N__37856),
            .I(N__37853));
    LocalMux I__7588 (
            .O(N__37853),
            .I(N__37850));
    Span4Mux_v I__7587 (
            .O(N__37850),
            .I(N__37847));
    Odrv4 I__7586 (
            .O(N__37847),
            .I(sDAC_data_RNO_24Z0Z_6));
    CascadeMux I__7585 (
            .O(N__37844),
            .I(sDAC_data_2_39_ns_1_6_cascade_));
    InMux I__7584 (
            .O(N__37841),
            .I(N__37838));
    LocalMux I__7583 (
            .O(N__37838),
            .I(N__37835));
    Span4Mux_h I__7582 (
            .O(N__37835),
            .I(N__37832));
    Odrv4 I__7581 (
            .O(N__37832),
            .I(sDAC_data_RNO_23Z0Z_6));
    InMux I__7580 (
            .O(N__37829),
            .I(N__37826));
    LocalMux I__7579 (
            .O(N__37826),
            .I(N__37823));
    Span4Mux_v I__7578 (
            .O(N__37823),
            .I(N__37820));
    Span4Mux_h I__7577 (
            .O(N__37820),
            .I(N__37817));
    Odrv4 I__7576 (
            .O(N__37817),
            .I(sDAC_data_RNO_11Z0Z_6));
    InMux I__7575 (
            .O(N__37814),
            .I(N__37811));
    LocalMux I__7574 (
            .O(N__37811),
            .I(sDAC_mem_28Z0Z_2));
    CEMux I__7573 (
            .O(N__37808),
            .I(N__37803));
    CEMux I__7572 (
            .O(N__37807),
            .I(N__37800));
    CEMux I__7571 (
            .O(N__37806),
            .I(N__37797));
    LocalMux I__7570 (
            .O(N__37803),
            .I(N__37793));
    LocalMux I__7569 (
            .O(N__37800),
            .I(N__37790));
    LocalMux I__7568 (
            .O(N__37797),
            .I(N__37786));
    CEMux I__7567 (
            .O(N__37796),
            .I(N__37783));
    Span4Mux_h I__7566 (
            .O(N__37793),
            .I(N__37780));
    Span4Mux_v I__7565 (
            .O(N__37790),
            .I(N__37777));
    CEMux I__7564 (
            .O(N__37789),
            .I(N__37774));
    Span4Mux_v I__7563 (
            .O(N__37786),
            .I(N__37771));
    LocalMux I__7562 (
            .O(N__37783),
            .I(N__37768));
    Span4Mux_h I__7561 (
            .O(N__37780),
            .I(N__37765));
    Span4Mux_h I__7560 (
            .O(N__37777),
            .I(N__37760));
    LocalMux I__7559 (
            .O(N__37774),
            .I(N__37760));
    Span4Mux_h I__7558 (
            .O(N__37771),
            .I(N__37755));
    Span4Mux_v I__7557 (
            .O(N__37768),
            .I(N__37755));
    Span4Mux_v I__7556 (
            .O(N__37765),
            .I(N__37752));
    Span4Mux_v I__7555 (
            .O(N__37760),
            .I(N__37749));
    Span4Mux_h I__7554 (
            .O(N__37755),
            .I(N__37746));
    Odrv4 I__7553 (
            .O(N__37752),
            .I(sDAC_mem_28_1_sqmuxa));
    Odrv4 I__7552 (
            .O(N__37749),
            .I(sDAC_mem_28_1_sqmuxa));
    Odrv4 I__7551 (
            .O(N__37746),
            .I(sDAC_mem_28_1_sqmuxa));
    InMux I__7550 (
            .O(N__37739),
            .I(N__37736));
    LocalMux I__7549 (
            .O(N__37736),
            .I(N__37733));
    Span4Mux_h I__7548 (
            .O(N__37733),
            .I(N__37730));
    Span4Mux_h I__7547 (
            .O(N__37730),
            .I(N__37727));
    Odrv4 I__7546 (
            .O(N__37727),
            .I(sDAC_mem_30Z0Z_2));
    InMux I__7545 (
            .O(N__37724),
            .I(N__37721));
    LocalMux I__7544 (
            .O(N__37721),
            .I(N__37718));
    Span12Mux_h I__7543 (
            .O(N__37718),
            .I(N__37715));
    Odrv12 I__7542 (
            .O(N__37715),
            .I(sDAC_mem_31Z0Z_2));
    InMux I__7541 (
            .O(N__37712),
            .I(N__37709));
    LocalMux I__7540 (
            .O(N__37709),
            .I(sDAC_data_RNO_24Z0Z_5));
    InMux I__7539 (
            .O(N__37706),
            .I(N__37703));
    LocalMux I__7538 (
            .O(N__37703),
            .I(N__37700));
    Span12Mux_h I__7537 (
            .O(N__37700),
            .I(N__37697));
    Odrv12 I__7536 (
            .O(N__37697),
            .I(sDAC_mem_26Z0Z_3));
    InMux I__7535 (
            .O(N__37694),
            .I(N__37691));
    LocalMux I__7534 (
            .O(N__37691),
            .I(N__37688));
    Span4Mux_h I__7533 (
            .O(N__37688),
            .I(N__37685));
    Odrv4 I__7532 (
            .O(N__37685),
            .I(sDAC_mem_27Z0Z_3));
    InMux I__7531 (
            .O(N__37682),
            .I(N__37679));
    LocalMux I__7530 (
            .O(N__37679),
            .I(sDAC_data_RNO_31Z0Z_6));
    InMux I__7529 (
            .O(N__37676),
            .I(N__37673));
    LocalMux I__7528 (
            .O(N__37673),
            .I(N__37670));
    Span4Mux_h I__7527 (
            .O(N__37670),
            .I(N__37667));
    Odrv4 I__7526 (
            .O(N__37667),
            .I(sDAC_data_RNO_5Z0Z_3));
    InMux I__7525 (
            .O(N__37664),
            .I(N__37661));
    LocalMux I__7524 (
            .O(N__37661),
            .I(sDAC_data_RNO_2Z0Z_3));
    CascadeMux I__7523 (
            .O(N__37658),
            .I(sDAC_data_RNO_1Z0Z_3_cascade_));
    InMux I__7522 (
            .O(N__37655),
            .I(N__37652));
    LocalMux I__7521 (
            .O(N__37652),
            .I(N__37649));
    Span4Mux_v I__7520 (
            .O(N__37649),
            .I(N__37646));
    Span4Mux_v I__7519 (
            .O(N__37646),
            .I(N__37643));
    Odrv4 I__7518 (
            .O(N__37643),
            .I(sEEDACZ0Z_0));
    CascadeMux I__7517 (
            .O(N__37640),
            .I(sDAC_data_2_3_cascade_));
    InMux I__7516 (
            .O(N__37637),
            .I(N__37624));
    InMux I__7515 (
            .O(N__37636),
            .I(N__37621));
    InMux I__7514 (
            .O(N__37635),
            .I(N__37618));
    InMux I__7513 (
            .O(N__37634),
            .I(N__37611));
    InMux I__7512 (
            .O(N__37633),
            .I(N__37611));
    InMux I__7511 (
            .O(N__37632),
            .I(N__37611));
    InMux I__7510 (
            .O(N__37631),
            .I(N__37608));
    InMux I__7509 (
            .O(N__37630),
            .I(N__37605));
    InMux I__7508 (
            .O(N__37629),
            .I(N__37602));
    InMux I__7507 (
            .O(N__37628),
            .I(N__37599));
    InMux I__7506 (
            .O(N__37627),
            .I(N__37596));
    LocalMux I__7505 (
            .O(N__37624),
            .I(N__37593));
    LocalMux I__7504 (
            .O(N__37621),
            .I(N__37590));
    LocalMux I__7503 (
            .O(N__37618),
            .I(N__37585));
    LocalMux I__7502 (
            .O(N__37611),
            .I(N__37585));
    LocalMux I__7501 (
            .O(N__37608),
            .I(N__37579));
    LocalMux I__7500 (
            .O(N__37605),
            .I(N__37576));
    LocalMux I__7499 (
            .O(N__37602),
            .I(N__37573));
    LocalMux I__7498 (
            .O(N__37599),
            .I(N__37564));
    LocalMux I__7497 (
            .O(N__37596),
            .I(N__37564));
    Span4Mux_h I__7496 (
            .O(N__37593),
            .I(N__37564));
    Span4Mux_h I__7495 (
            .O(N__37590),
            .I(N__37564));
    Span4Mux_v I__7494 (
            .O(N__37585),
            .I(N__37561));
    InMux I__7493 (
            .O(N__37584),
            .I(N__37554));
    InMux I__7492 (
            .O(N__37583),
            .I(N__37554));
    InMux I__7491 (
            .O(N__37582),
            .I(N__37554));
    Span4Mux_h I__7490 (
            .O(N__37579),
            .I(N__37551));
    Span4Mux_v I__7489 (
            .O(N__37576),
            .I(N__37548));
    Span4Mux_v I__7488 (
            .O(N__37573),
            .I(N__37545));
    Span4Mux_v I__7487 (
            .O(N__37564),
            .I(N__37542));
    Span4Mux_v I__7486 (
            .O(N__37561),
            .I(N__37539));
    LocalMux I__7485 (
            .O(N__37554),
            .I(un5_sdacdyn_cry_23_c_RNIELGZ0Z28));
    Odrv4 I__7484 (
            .O(N__37551),
            .I(un5_sdacdyn_cry_23_c_RNIELGZ0Z28));
    Odrv4 I__7483 (
            .O(N__37548),
            .I(un5_sdacdyn_cry_23_c_RNIELGZ0Z28));
    Odrv4 I__7482 (
            .O(N__37545),
            .I(un5_sdacdyn_cry_23_c_RNIELGZ0Z28));
    Odrv4 I__7481 (
            .O(N__37542),
            .I(un5_sdacdyn_cry_23_c_RNIELGZ0Z28));
    Odrv4 I__7480 (
            .O(N__37539),
            .I(un5_sdacdyn_cry_23_c_RNIELGZ0Z28));
    InMux I__7479 (
            .O(N__37526),
            .I(N__37523));
    LocalMux I__7478 (
            .O(N__37523),
            .I(N__37520));
    Span4Mux_h I__7477 (
            .O(N__37520),
            .I(N__37517));
    Span4Mux_v I__7476 (
            .O(N__37517),
            .I(N__37514));
    Odrv4 I__7475 (
            .O(N__37514),
            .I(sDAC_dataZ0Z_3));
    InMux I__7474 (
            .O(N__37511),
            .I(N__37508));
    LocalMux I__7473 (
            .O(N__37508),
            .I(N__37505));
    Span4Mux_v I__7472 (
            .O(N__37505),
            .I(N__37502));
    Odrv4 I__7471 (
            .O(N__37502),
            .I(sDAC_data_RNO_21Z0Z_3));
    InMux I__7470 (
            .O(N__37499),
            .I(N__37496));
    LocalMux I__7469 (
            .O(N__37496),
            .I(N__37493));
    Span4Mux_v I__7468 (
            .O(N__37493),
            .I(N__37490));
    Odrv4 I__7467 (
            .O(N__37490),
            .I(sDAC_data_RNO_20Z0Z_3));
    CascadeMux I__7466 (
            .O(N__37487),
            .I(N__37482));
    InMux I__7465 (
            .O(N__37486),
            .I(N__37478));
    InMux I__7464 (
            .O(N__37485),
            .I(N__37473));
    InMux I__7463 (
            .O(N__37482),
            .I(N__37473));
    CascadeMux I__7462 (
            .O(N__37481),
            .I(N__37468));
    LocalMux I__7461 (
            .O(N__37478),
            .I(N__37463));
    LocalMux I__7460 (
            .O(N__37473),
            .I(N__37463));
    CascadeMux I__7459 (
            .O(N__37472),
            .I(N__37458));
    InMux I__7458 (
            .O(N__37471),
            .I(N__37449));
    InMux I__7457 (
            .O(N__37468),
            .I(N__37449));
    Span4Mux_v I__7456 (
            .O(N__37463),
            .I(N__37446));
    InMux I__7455 (
            .O(N__37462),
            .I(N__37443));
    InMux I__7454 (
            .O(N__37461),
            .I(N__37436));
    InMux I__7453 (
            .O(N__37458),
            .I(N__37433));
    InMux I__7452 (
            .O(N__37457),
            .I(N__37428));
    InMux I__7451 (
            .O(N__37456),
            .I(N__37428));
    InMux I__7450 (
            .O(N__37455),
            .I(N__37423));
    InMux I__7449 (
            .O(N__37454),
            .I(N__37423));
    LocalMux I__7448 (
            .O(N__37449),
            .I(N__37420));
    Span4Mux_h I__7447 (
            .O(N__37446),
            .I(N__37416));
    LocalMux I__7446 (
            .O(N__37443),
            .I(N__37413));
    InMux I__7445 (
            .O(N__37442),
            .I(N__37408));
    InMux I__7444 (
            .O(N__37441),
            .I(N__37408));
    InMux I__7443 (
            .O(N__37440),
            .I(N__37403));
    InMux I__7442 (
            .O(N__37439),
            .I(N__37403));
    LocalMux I__7441 (
            .O(N__37436),
            .I(N__37396));
    LocalMux I__7440 (
            .O(N__37433),
            .I(N__37396));
    LocalMux I__7439 (
            .O(N__37428),
            .I(N__37396));
    LocalMux I__7438 (
            .O(N__37423),
            .I(N__37391));
    Span4Mux_h I__7437 (
            .O(N__37420),
            .I(N__37391));
    InMux I__7436 (
            .O(N__37419),
            .I(N__37387));
    Sp12to4 I__7435 (
            .O(N__37416),
            .I(N__37382));
    Sp12to4 I__7434 (
            .O(N__37413),
            .I(N__37382));
    LocalMux I__7433 (
            .O(N__37408),
            .I(N__37379));
    LocalMux I__7432 (
            .O(N__37403),
            .I(N__37376));
    Span4Mux_v I__7431 (
            .O(N__37396),
            .I(N__37371));
    Span4Mux_v I__7430 (
            .O(N__37391),
            .I(N__37371));
    InMux I__7429 (
            .O(N__37390),
            .I(N__37368));
    LocalMux I__7428 (
            .O(N__37387),
            .I(sDAC_mem_pointerZ0Z_4));
    Odrv12 I__7427 (
            .O(N__37382),
            .I(sDAC_mem_pointerZ0Z_4));
    Odrv4 I__7426 (
            .O(N__37379),
            .I(sDAC_mem_pointerZ0Z_4));
    Odrv12 I__7425 (
            .O(N__37376),
            .I(sDAC_mem_pointerZ0Z_4));
    Odrv4 I__7424 (
            .O(N__37371),
            .I(sDAC_mem_pointerZ0Z_4));
    LocalMux I__7423 (
            .O(N__37368),
            .I(sDAC_mem_pointerZ0Z_4));
    InMux I__7422 (
            .O(N__37355),
            .I(N__37352));
    LocalMux I__7421 (
            .O(N__37352),
            .I(N__37348));
    InMux I__7420 (
            .O(N__37351),
            .I(N__37345));
    Span4Mux_v I__7419 (
            .O(N__37348),
            .I(N__37336));
    LocalMux I__7418 (
            .O(N__37345),
            .I(N__37336));
    InMux I__7417 (
            .O(N__37344),
            .I(N__37331));
    InMux I__7416 (
            .O(N__37343),
            .I(N__37328));
    InMux I__7415 (
            .O(N__37342),
            .I(N__37324));
    InMux I__7414 (
            .O(N__37341),
            .I(N__37321));
    Span4Mux_h I__7413 (
            .O(N__37336),
            .I(N__37318));
    InMux I__7412 (
            .O(N__37335),
            .I(N__37315));
    InMux I__7411 (
            .O(N__37334),
            .I(N__37312));
    LocalMux I__7410 (
            .O(N__37331),
            .I(N__37309));
    LocalMux I__7409 (
            .O(N__37328),
            .I(N__37306));
    InMux I__7408 (
            .O(N__37327),
            .I(N__37302));
    LocalMux I__7407 (
            .O(N__37324),
            .I(N__37297));
    LocalMux I__7406 (
            .O(N__37321),
            .I(N__37297));
    Span4Mux_h I__7405 (
            .O(N__37318),
            .I(N__37290));
    LocalMux I__7404 (
            .O(N__37315),
            .I(N__37290));
    LocalMux I__7403 (
            .O(N__37312),
            .I(N__37290));
    Span4Mux_h I__7402 (
            .O(N__37309),
            .I(N__37285));
    Span4Mux_v I__7401 (
            .O(N__37306),
            .I(N__37285));
    InMux I__7400 (
            .O(N__37305),
            .I(N__37282));
    LocalMux I__7399 (
            .O(N__37302),
            .I(sDAC_mem_pointerZ0Z_3));
    Odrv4 I__7398 (
            .O(N__37297),
            .I(sDAC_mem_pointerZ0Z_3));
    Odrv4 I__7397 (
            .O(N__37290),
            .I(sDAC_mem_pointerZ0Z_3));
    Odrv4 I__7396 (
            .O(N__37285),
            .I(sDAC_mem_pointerZ0Z_3));
    LocalMux I__7395 (
            .O(N__37282),
            .I(sDAC_mem_pointerZ0Z_3));
    CascadeMux I__7394 (
            .O(N__37271),
            .I(sDAC_data_RNO_10Z0Z_3_cascade_));
    InMux I__7393 (
            .O(N__37268),
            .I(N__37265));
    LocalMux I__7392 (
            .O(N__37265),
            .I(N__37262));
    Span4Mux_h I__7391 (
            .O(N__37262),
            .I(N__37259));
    Odrv4 I__7390 (
            .O(N__37259),
            .I(sDAC_data_RNO_11Z0Z_3));
    InMux I__7389 (
            .O(N__37256),
            .I(N__37253));
    LocalMux I__7388 (
            .O(N__37253),
            .I(sDAC_data_2_41_ns_1_3));
    InMux I__7387 (
            .O(N__37250),
            .I(N__37247));
    LocalMux I__7386 (
            .O(N__37247),
            .I(sDAC_data_RNO_15Z0Z_3));
    InMux I__7385 (
            .O(N__37244),
            .I(N__37241));
    LocalMux I__7384 (
            .O(N__37241),
            .I(sDAC_data_2_14_ns_1_3));
    InMux I__7383 (
            .O(N__37238),
            .I(N__37235));
    LocalMux I__7382 (
            .O(N__37235),
            .I(N__37232));
    Span4Mux_v I__7381 (
            .O(N__37232),
            .I(N__37229));
    Odrv4 I__7380 (
            .O(N__37229),
            .I(sDAC_data_RNO_28Z0Z_3));
    InMux I__7379 (
            .O(N__37226),
            .I(N__37223));
    LocalMux I__7378 (
            .O(N__37223),
            .I(sDAC_data_RNO_29Z0Z_3));
    InMux I__7377 (
            .O(N__37220),
            .I(N__37217));
    LocalMux I__7376 (
            .O(N__37217),
            .I(sDAC_data_2_32_ns_1_3));
    InMux I__7375 (
            .O(N__37214),
            .I(N__37211));
    LocalMux I__7374 (
            .O(N__37211),
            .I(N__37208));
    Odrv12 I__7373 (
            .O(N__37208),
            .I(sDAC_data_2_39_ns_1_5));
    InMux I__7372 (
            .O(N__37205),
            .I(N__37202));
    LocalMux I__7371 (
            .O(N__37202),
            .I(N__37199));
    Odrv4 I__7370 (
            .O(N__37199),
            .I(sDAC_data_RNO_11Z0Z_5));
    InMux I__7369 (
            .O(N__37196),
            .I(N__37193));
    LocalMux I__7368 (
            .O(N__37193),
            .I(N__37190));
    Span4Mux_v I__7367 (
            .O(N__37190),
            .I(N__37187));
    Span4Mux_v I__7366 (
            .O(N__37187),
            .I(N__37184));
    Odrv4 I__7365 (
            .O(N__37184),
            .I(sDAC_mem_pointerZ0Z_7));
    InMux I__7364 (
            .O(N__37181),
            .I(N__37178));
    LocalMux I__7363 (
            .O(N__37178),
            .I(N__37175));
    Odrv12 I__7362 (
            .O(N__37175),
            .I(sDAC_mem_pointerZ0Z_6));
    InMux I__7361 (
            .O(N__37172),
            .I(N__37169));
    LocalMux I__7360 (
            .O(N__37169),
            .I(un17_sdacdyn_0));
    InMux I__7359 (
            .O(N__37166),
            .I(N__37163));
    LocalMux I__7358 (
            .O(N__37163),
            .I(N__37160));
    Span4Mux_v I__7357 (
            .O(N__37160),
            .I(N__37157));
    Odrv4 I__7356 (
            .O(N__37157),
            .I(sDAC_data_RNO_5Z0Z_5));
    InMux I__7355 (
            .O(N__37154),
            .I(N__37151));
    LocalMux I__7354 (
            .O(N__37151),
            .I(sDAC_data_RNO_2Z0Z_5));
    CascadeMux I__7353 (
            .O(N__37148),
            .I(sDAC_data_RNO_1Z0Z_5_cascade_));
    InMux I__7352 (
            .O(N__37145),
            .I(N__37142));
    LocalMux I__7351 (
            .O(N__37142),
            .I(N__37139));
    Span4Mux_v I__7350 (
            .O(N__37139),
            .I(N__37136));
    Span4Mux_v I__7349 (
            .O(N__37136),
            .I(N__37133));
    Odrv4 I__7348 (
            .O(N__37133),
            .I(sEEDACZ0Z_2));
    CascadeMux I__7347 (
            .O(N__37130),
            .I(sDAC_data_2_5_cascade_));
    InMux I__7346 (
            .O(N__37127),
            .I(N__37124));
    LocalMux I__7345 (
            .O(N__37124),
            .I(N__37121));
    Span4Mux_h I__7344 (
            .O(N__37121),
            .I(N__37118));
    Span4Mux_v I__7343 (
            .O(N__37118),
            .I(N__37115));
    Span4Mux_h I__7342 (
            .O(N__37115),
            .I(N__37112));
    Span4Mux_h I__7341 (
            .O(N__37112),
            .I(N__37109));
    Odrv4 I__7340 (
            .O(N__37109),
            .I(sDAC_dataZ0Z_5));
    InMux I__7339 (
            .O(N__37106),
            .I(N__37103));
    LocalMux I__7338 (
            .O(N__37103),
            .I(sDAC_data_RNO_15Z0Z_5));
    InMux I__7337 (
            .O(N__37100),
            .I(N__37097));
    LocalMux I__7336 (
            .O(N__37097),
            .I(sDAC_data_2_14_ns_1_5));
    InMux I__7335 (
            .O(N__37094),
            .I(N__37091));
    LocalMux I__7334 (
            .O(N__37091),
            .I(sDAC_data_RNO_29Z0Z_5));
    InMux I__7333 (
            .O(N__37088),
            .I(N__37085));
    LocalMux I__7332 (
            .O(N__37085),
            .I(N__37082));
    Span4Mux_h I__7331 (
            .O(N__37082),
            .I(N__37079));
    Span4Mux_v I__7330 (
            .O(N__37079),
            .I(N__37076));
    Odrv4 I__7329 (
            .O(N__37076),
            .I(sDAC_data_RNO_28Z0Z_5));
    InMux I__7328 (
            .O(N__37073),
            .I(N__37070));
    LocalMux I__7327 (
            .O(N__37070),
            .I(N__37067));
    Odrv4 I__7326 (
            .O(N__37067),
            .I(sDAC_data_RNO_20Z0Z_5));
    CascadeMux I__7325 (
            .O(N__37064),
            .I(sDAC_data_2_32_ns_1_5_cascade_));
    InMux I__7324 (
            .O(N__37061),
            .I(N__37058));
    LocalMux I__7323 (
            .O(N__37058),
            .I(N__37055));
    Span4Mux_h I__7322 (
            .O(N__37055),
            .I(N__37052));
    Odrv4 I__7321 (
            .O(N__37052),
            .I(sDAC_data_RNO_21Z0Z_5));
    CascadeMux I__7320 (
            .O(N__37049),
            .I(sDAC_data_RNO_10Z0Z_5_cascade_));
    InMux I__7319 (
            .O(N__37046),
            .I(N__37043));
    LocalMux I__7318 (
            .O(N__37043),
            .I(sDAC_data_2_41_ns_1_5));
    InMux I__7317 (
            .O(N__37040),
            .I(N__37037));
    LocalMux I__7316 (
            .O(N__37037),
            .I(N__37034));
    Span4Mux_h I__7315 (
            .O(N__37034),
            .I(N__37031));
    Odrv4 I__7314 (
            .O(N__37031),
            .I(sDAC_mem_9Z0Z_6));
    InMux I__7313 (
            .O(N__37028),
            .I(N__37025));
    LocalMux I__7312 (
            .O(N__37025),
            .I(N__37022));
    Span4Mux_h I__7311 (
            .O(N__37022),
            .I(N__37019));
    Odrv4 I__7310 (
            .O(N__37019),
            .I(sDAC_mem_9Z0Z_7));
    InMux I__7309 (
            .O(N__37016),
            .I(N__37013));
    LocalMux I__7308 (
            .O(N__37013),
            .I(N__37010));
    Odrv12 I__7307 (
            .O(N__37010),
            .I(sDAC_mem_15Z0Z_6));
    InMux I__7306 (
            .O(N__37007),
            .I(N__37004));
    LocalMux I__7305 (
            .O(N__37004),
            .I(N__37001));
    Span4Mux_h I__7304 (
            .O(N__37001),
            .I(N__36998));
    Span4Mux_h I__7303 (
            .O(N__36998),
            .I(N__36995));
    Odrv4 I__7302 (
            .O(N__36995),
            .I(sDAC_mem_14Z0Z_6));
    CascadeMux I__7301 (
            .O(N__36992),
            .I(sDAC_data_RNO_18Z0Z_9_cascade_));
    InMux I__7300 (
            .O(N__36989),
            .I(N__36986));
    LocalMux I__7299 (
            .O(N__36986),
            .I(sDAC_data_RNO_19Z0Z_9));
    InMux I__7298 (
            .O(N__36983),
            .I(N__36980));
    LocalMux I__7297 (
            .O(N__36980),
            .I(N__36977));
    Span4Mux_h I__7296 (
            .O(N__36977),
            .I(N__36974));
    Odrv4 I__7295 (
            .O(N__36974),
            .I(sDAC_data_2_24_ns_1_9));
    InMux I__7294 (
            .O(N__36971),
            .I(N__36968));
    LocalMux I__7293 (
            .O(N__36968),
            .I(sDAC_mem_12Z0Z_6));
    CEMux I__7292 (
            .O(N__36965),
            .I(N__36961));
    CEMux I__7291 (
            .O(N__36964),
            .I(N__36956));
    LocalMux I__7290 (
            .O(N__36961),
            .I(N__36953));
    CEMux I__7289 (
            .O(N__36960),
            .I(N__36949));
    CEMux I__7288 (
            .O(N__36959),
            .I(N__36946));
    LocalMux I__7287 (
            .O(N__36956),
            .I(N__36943));
    Span4Mux_h I__7286 (
            .O(N__36953),
            .I(N__36940));
    CEMux I__7285 (
            .O(N__36952),
            .I(N__36937));
    LocalMux I__7284 (
            .O(N__36949),
            .I(N__36934));
    LocalMux I__7283 (
            .O(N__36946),
            .I(N__36931));
    Span4Mux_h I__7282 (
            .O(N__36943),
            .I(N__36924));
    Span4Mux_v I__7281 (
            .O(N__36940),
            .I(N__36924));
    LocalMux I__7280 (
            .O(N__36937),
            .I(N__36924));
    Span4Mux_v I__7279 (
            .O(N__36934),
            .I(N__36921));
    Span4Mux_h I__7278 (
            .O(N__36931),
            .I(N__36918));
    Span4Mux_h I__7277 (
            .O(N__36924),
            .I(N__36915));
    Span4Mux_h I__7276 (
            .O(N__36921),
            .I(N__36910));
    Span4Mux_h I__7275 (
            .O(N__36918),
            .I(N__36910));
    Span4Mux_h I__7274 (
            .O(N__36915),
            .I(N__36907));
    Odrv4 I__7273 (
            .O(N__36910),
            .I(sDAC_mem_12_1_sqmuxa));
    Odrv4 I__7272 (
            .O(N__36907),
            .I(sDAC_mem_12_1_sqmuxa));
    CascadeMux I__7271 (
            .O(N__36902),
            .I(op_le_op_le_un15_sdacdynlt4_cascade_));
    InMux I__7270 (
            .O(N__36899),
            .I(N__36896));
    LocalMux I__7269 (
            .O(N__36896),
            .I(N__36893));
    Span4Mux_h I__7268 (
            .O(N__36893),
            .I(N__36890));
    Sp12to4 I__7267 (
            .O(N__36890),
            .I(N__36887));
    Odrv12 I__7266 (
            .O(N__36887),
            .I(un17_sdacdyn_1));
    CascadeMux I__7265 (
            .O(N__36884),
            .I(sDAC_data_RNO_26Z0Z_7_cascade_));
    InMux I__7264 (
            .O(N__36881),
            .I(N__36878));
    LocalMux I__7263 (
            .O(N__36878),
            .I(N__36875));
    Span4Mux_h I__7262 (
            .O(N__36875),
            .I(N__36872));
    Odrv4 I__7261 (
            .O(N__36872),
            .I(sDAC_data_RNO_14Z0Z_7));
    InMux I__7260 (
            .O(N__36869),
            .I(N__36866));
    LocalMux I__7259 (
            .O(N__36866),
            .I(sDAC_mem_32Z0Z_4));
    CascadeMux I__7258 (
            .O(N__36863),
            .I(sDAC_data_RNO_26Z0Z_8_cascade_));
    CascadeMux I__7257 (
            .O(N__36860),
            .I(N__36857));
    InMux I__7256 (
            .O(N__36857),
            .I(N__36854));
    LocalMux I__7255 (
            .O(N__36854),
            .I(N__36851));
    Span4Mux_h I__7254 (
            .O(N__36851),
            .I(N__36848));
    Odrv4 I__7253 (
            .O(N__36848),
            .I(sDAC_data_RNO_14Z0Z_8));
    InMux I__7252 (
            .O(N__36845),
            .I(N__36842));
    LocalMux I__7251 (
            .O(N__36842),
            .I(N__36839));
    Span4Mux_v I__7250 (
            .O(N__36839),
            .I(N__36836));
    Odrv4 I__7249 (
            .O(N__36836),
            .I(sDAC_mem_9Z0Z_0));
    InMux I__7248 (
            .O(N__36833),
            .I(N__36830));
    LocalMux I__7247 (
            .O(N__36830),
            .I(N__36827));
    Span4Mux_h I__7246 (
            .O(N__36827),
            .I(N__36824));
    Odrv4 I__7245 (
            .O(N__36824),
            .I(sDAC_mem_9Z0Z_1));
    InMux I__7244 (
            .O(N__36821),
            .I(N__36818));
    LocalMux I__7243 (
            .O(N__36818),
            .I(sDAC_mem_9Z0Z_2));
    InMux I__7242 (
            .O(N__36815),
            .I(N__36812));
    LocalMux I__7241 (
            .O(N__36812),
            .I(N__36809));
    Span4Mux_h I__7240 (
            .O(N__36809),
            .I(N__36806));
    Span4Mux_h I__7239 (
            .O(N__36806),
            .I(N__36803));
    Odrv4 I__7238 (
            .O(N__36803),
            .I(sDAC_mem_9Z0Z_3));
    InMux I__7237 (
            .O(N__36800),
            .I(N__36797));
    LocalMux I__7236 (
            .O(N__36797),
            .I(N__36794));
    Sp12to4 I__7235 (
            .O(N__36794),
            .I(N__36791));
    Odrv12 I__7234 (
            .O(N__36791),
            .I(sDAC_mem_9Z0Z_4));
    InMux I__7233 (
            .O(N__36788),
            .I(N__36785));
    LocalMux I__7232 (
            .O(N__36785),
            .I(N__36782));
    Span4Mux_v I__7231 (
            .O(N__36782),
            .I(N__36779));
    Odrv4 I__7230 (
            .O(N__36779),
            .I(sDAC_mem_9Z0Z_5));
    InMux I__7229 (
            .O(N__36776),
            .I(N__36773));
    LocalMux I__7228 (
            .O(N__36773),
            .I(N__36770));
    Span4Mux_h I__7227 (
            .O(N__36770),
            .I(N__36767));
    Odrv4 I__7226 (
            .O(N__36767),
            .I(sDAC_mem_23Z0Z_3));
    InMux I__7225 (
            .O(N__36764),
            .I(N__36761));
    LocalMux I__7224 (
            .O(N__36761),
            .I(N__36758));
    Span4Mux_v I__7223 (
            .O(N__36758),
            .I(N__36755));
    Span4Mux_v I__7222 (
            .O(N__36755),
            .I(N__36752));
    Span4Mux_v I__7221 (
            .O(N__36752),
            .I(N__36749));
    Odrv4 I__7220 (
            .O(N__36749),
            .I(sDAC_mem_23Z0Z_4));
    InMux I__7219 (
            .O(N__36746),
            .I(N__36743));
    LocalMux I__7218 (
            .O(N__36743),
            .I(N__36740));
    Span4Mux_v I__7217 (
            .O(N__36740),
            .I(N__36737));
    Sp12to4 I__7216 (
            .O(N__36737),
            .I(N__36734));
    Span12Mux_h I__7215 (
            .O(N__36734),
            .I(N__36731));
    Odrv12 I__7214 (
            .O(N__36731),
            .I(sDAC_mem_23Z0Z_5));
    InMux I__7213 (
            .O(N__36728),
            .I(N__36725));
    LocalMux I__7212 (
            .O(N__36725),
            .I(N__36722));
    Span12Mux_v I__7211 (
            .O(N__36722),
            .I(N__36719));
    Odrv12 I__7210 (
            .O(N__36719),
            .I(sDAC_mem_23Z0Z_6));
    InMux I__7209 (
            .O(N__36716),
            .I(N__36713));
    LocalMux I__7208 (
            .O(N__36713),
            .I(N__36710));
    Span4Mux_h I__7207 (
            .O(N__36710),
            .I(N__36707));
    Span4Mux_v I__7206 (
            .O(N__36707),
            .I(N__36704));
    Odrv4 I__7205 (
            .O(N__36704),
            .I(sDAC_mem_23Z0Z_7));
    CEMux I__7204 (
            .O(N__36701),
            .I(N__36698));
    LocalMux I__7203 (
            .O(N__36698),
            .I(N__36695));
    Span4Mux_v I__7202 (
            .O(N__36695),
            .I(N__36692));
    Span4Mux_h I__7201 (
            .O(N__36692),
            .I(N__36689));
    Span4Mux_h I__7200 (
            .O(N__36689),
            .I(N__36686));
    Odrv4 I__7199 (
            .O(N__36686),
            .I(sDAC_mem_23_1_sqmuxa));
    CascadeMux I__7198 (
            .O(N__36683),
            .I(sDAC_data_RNO_26Z0Z_6_cascade_));
    InMux I__7197 (
            .O(N__36680),
            .I(N__36677));
    LocalMux I__7196 (
            .O(N__36677),
            .I(sDAC_mem_32Z0Z_3));
    InMux I__7195 (
            .O(N__36674),
            .I(N__36671));
    LocalMux I__7194 (
            .O(N__36671),
            .I(N__36668));
    Span4Mux_v I__7193 (
            .O(N__36668),
            .I(N__36665));
    Odrv4 I__7192 (
            .O(N__36665),
            .I(sDAC_data_RNO_14Z0Z_6));
    InMux I__7191 (
            .O(N__36662),
            .I(N__36659));
    LocalMux I__7190 (
            .O(N__36659),
            .I(N__36656));
    Odrv4 I__7189 (
            .O(N__36656),
            .I(sDAC_mem_20Z0Z_4));
    InMux I__7188 (
            .O(N__36653),
            .I(N__36650));
    LocalMux I__7187 (
            .O(N__36650),
            .I(N__36647));
    Sp12to4 I__7186 (
            .O(N__36647),
            .I(N__36644));
    Span12Mux_v I__7185 (
            .O(N__36644),
            .I(N__36641));
    Odrv12 I__7184 (
            .O(N__36641),
            .I(sDAC_mem_20Z0Z_7));
    CEMux I__7183 (
            .O(N__36638),
            .I(N__36634));
    CEMux I__7182 (
            .O(N__36637),
            .I(N__36631));
    LocalMux I__7181 (
            .O(N__36634),
            .I(N__36628));
    LocalMux I__7180 (
            .O(N__36631),
            .I(N__36625));
    Span4Mux_h I__7179 (
            .O(N__36628),
            .I(N__36622));
    Span12Mux_v I__7178 (
            .O(N__36625),
            .I(N__36619));
    Span4Mux_v I__7177 (
            .O(N__36622),
            .I(N__36616));
    Odrv12 I__7176 (
            .O(N__36619),
            .I(sDAC_mem_20_1_sqmuxa));
    Odrv4 I__7175 (
            .O(N__36616),
            .I(sDAC_mem_20_1_sqmuxa));
    InMux I__7174 (
            .O(N__36611),
            .I(N__36608));
    LocalMux I__7173 (
            .O(N__36608),
            .I(N__36605));
    Span4Mux_h I__7172 (
            .O(N__36605),
            .I(N__36602));
    Span4Mux_v I__7171 (
            .O(N__36602),
            .I(N__36599));
    Odrv4 I__7170 (
            .O(N__36599),
            .I(sDAC_mem_6Z0Z_0));
    InMux I__7169 (
            .O(N__36596),
            .I(N__36593));
    LocalMux I__7168 (
            .O(N__36593),
            .I(N__36590));
    Span4Mux_h I__7167 (
            .O(N__36590),
            .I(N__36587));
    Span4Mux_v I__7166 (
            .O(N__36587),
            .I(N__36584));
    Odrv4 I__7165 (
            .O(N__36584),
            .I(sDAC_mem_6Z0Z_1));
    InMux I__7164 (
            .O(N__36581),
            .I(N__36578));
    LocalMux I__7163 (
            .O(N__36578),
            .I(N__36575));
    Span4Mux_h I__7162 (
            .O(N__36575),
            .I(N__36572));
    Odrv4 I__7161 (
            .O(N__36572),
            .I(sDAC_mem_6Z0Z_4));
    InMux I__7160 (
            .O(N__36569),
            .I(N__36566));
    LocalMux I__7159 (
            .O(N__36566),
            .I(N__36563));
    Span4Mux_h I__7158 (
            .O(N__36563),
            .I(N__36560));
    Span4Mux_v I__7157 (
            .O(N__36560),
            .I(N__36557));
    Odrv4 I__7156 (
            .O(N__36557),
            .I(sDAC_mem_6Z0Z_7));
    CEMux I__7155 (
            .O(N__36554),
            .I(N__36550));
    CEMux I__7154 (
            .O(N__36553),
            .I(N__36546));
    LocalMux I__7153 (
            .O(N__36550),
            .I(N__36543));
    CEMux I__7152 (
            .O(N__36549),
            .I(N__36540));
    LocalMux I__7151 (
            .O(N__36546),
            .I(N__36537));
    Span4Mux_v I__7150 (
            .O(N__36543),
            .I(N__36532));
    LocalMux I__7149 (
            .O(N__36540),
            .I(N__36532));
    Span4Mux_v I__7148 (
            .O(N__36537),
            .I(N__36529));
    Span4Mux_h I__7147 (
            .O(N__36532),
            .I(N__36526));
    Span4Mux_h I__7146 (
            .O(N__36529),
            .I(N__36523));
    Span4Mux_h I__7145 (
            .O(N__36526),
            .I(N__36520));
    Odrv4 I__7144 (
            .O(N__36523),
            .I(sDAC_mem_6_1_sqmuxa));
    Odrv4 I__7143 (
            .O(N__36520),
            .I(sDAC_mem_6_1_sqmuxa));
    InMux I__7142 (
            .O(N__36515),
            .I(N__36512));
    LocalMux I__7141 (
            .O(N__36512),
            .I(N__36509));
    Span4Mux_h I__7140 (
            .O(N__36509),
            .I(N__36506));
    Odrv4 I__7139 (
            .O(N__36506),
            .I(sDAC_mem_23Z0Z_0));
    InMux I__7138 (
            .O(N__36503),
            .I(N__36500));
    LocalMux I__7137 (
            .O(N__36500),
            .I(N__36497));
    Span4Mux_v I__7136 (
            .O(N__36497),
            .I(N__36494));
    Odrv4 I__7135 (
            .O(N__36494),
            .I(sDAC_mem_23Z0Z_1));
    InMux I__7134 (
            .O(N__36491),
            .I(N__36488));
    LocalMux I__7133 (
            .O(N__36488),
            .I(N__36485));
    Span4Mux_h I__7132 (
            .O(N__36485),
            .I(N__36482));
    Odrv4 I__7131 (
            .O(N__36482),
            .I(sDAC_mem_23Z0Z_2));
    CascadeMux I__7130 (
            .O(N__36479),
            .I(N__36476));
    InMux I__7129 (
            .O(N__36476),
            .I(N__36473));
    LocalMux I__7128 (
            .O(N__36473),
            .I(N__36470));
    Span4Mux_h I__7127 (
            .O(N__36470),
            .I(N__36467));
    Span4Mux_v I__7126 (
            .O(N__36467),
            .I(N__36464));
    Odrv4 I__7125 (
            .O(N__36464),
            .I(sDAC_mem_4Z0Z_5));
    InMux I__7124 (
            .O(N__36461),
            .I(N__36458));
    LocalMux I__7123 (
            .O(N__36458),
            .I(N__36455));
    Sp12to4 I__7122 (
            .O(N__36455),
            .I(N__36452));
    Odrv12 I__7121 (
            .O(N__36452),
            .I(sDAC_mem_4Z0Z_7));
    InMux I__7120 (
            .O(N__36449),
            .I(N__36446));
    LocalMux I__7119 (
            .O(N__36446),
            .I(N__36443));
    Span4Mux_v I__7118 (
            .O(N__36443),
            .I(N__36440));
    Odrv4 I__7117 (
            .O(N__36440),
            .I(sDAC_mem_20Z0Z_0));
    InMux I__7116 (
            .O(N__36437),
            .I(N__36434));
    LocalMux I__7115 (
            .O(N__36434),
            .I(N__36431));
    Span4Mux_v I__7114 (
            .O(N__36431),
            .I(N__36428));
    Odrv4 I__7113 (
            .O(N__36428),
            .I(sDAC_mem_20Z0Z_1));
    InMux I__7112 (
            .O(N__36425),
            .I(N__36422));
    LocalMux I__7111 (
            .O(N__36422),
            .I(N__36419));
    Span4Mux_h I__7110 (
            .O(N__36419),
            .I(N__36416));
    Odrv4 I__7109 (
            .O(N__36416),
            .I(sDAC_mem_20Z0Z_2));
    InMux I__7108 (
            .O(N__36413),
            .I(N__36410));
    LocalMux I__7107 (
            .O(N__36410),
            .I(N__36407));
    Odrv4 I__7106 (
            .O(N__36407),
            .I(sDAC_mem_20Z0Z_3));
    InMux I__7105 (
            .O(N__36404),
            .I(N__36401));
    LocalMux I__7104 (
            .O(N__36401),
            .I(N__36398));
    Span4Mux_h I__7103 (
            .O(N__36398),
            .I(N__36395));
    Sp12to4 I__7102 (
            .O(N__36395),
            .I(N__36392));
    Span12Mux_v I__7101 (
            .O(N__36392),
            .I(N__36389));
    Span12Mux_h I__7100 (
            .O(N__36389),
            .I(N__36385));
    InMux I__7099 (
            .O(N__36388),
            .I(N__36382));
    Odrv12 I__7098 (
            .O(N__36385),
            .I(sRAM_pointer_writeZ0Z_17));
    LocalMux I__7097 (
            .O(N__36382),
            .I(sRAM_pointer_writeZ0Z_17));
    CascadeMux I__7096 (
            .O(N__36377),
            .I(N__36374));
    InMux I__7095 (
            .O(N__36374),
            .I(N__36371));
    LocalMux I__7094 (
            .O(N__36371),
            .I(N__36368));
    Span4Mux_h I__7093 (
            .O(N__36368),
            .I(N__36364));
    InMux I__7092 (
            .O(N__36367),
            .I(N__36361));
    Odrv4 I__7091 (
            .O(N__36364),
            .I(sRAM_pointer_readZ0Z_17));
    LocalMux I__7090 (
            .O(N__36361),
            .I(sRAM_pointer_readZ0Z_17));
    IoInMux I__7089 (
            .O(N__36356),
            .I(N__36353));
    LocalMux I__7088 (
            .O(N__36353),
            .I(N__36350));
    IoSpan4Mux I__7087 (
            .O(N__36350),
            .I(N__36347));
    Span4Mux_s3_h I__7086 (
            .O(N__36347),
            .I(N__36344));
    Sp12to4 I__7085 (
            .O(N__36344),
            .I(N__36341));
    Odrv12 I__7084 (
            .O(N__36341),
            .I(RAM_ADD_c_17));
    InMux I__7083 (
            .O(N__36338),
            .I(N__36335));
    LocalMux I__7082 (
            .O(N__36335),
            .I(N__36332));
    Span4Mux_v I__7081 (
            .O(N__36332),
            .I(N__36329));
    Span4Mux_v I__7080 (
            .O(N__36329),
            .I(N__36326));
    Sp12to4 I__7079 (
            .O(N__36326),
            .I(N__36323));
    Span12Mux_h I__7078 (
            .O(N__36323),
            .I(N__36319));
    InMux I__7077 (
            .O(N__36322),
            .I(N__36316));
    Odrv12 I__7076 (
            .O(N__36319),
            .I(sRAM_pointer_writeZ0Z_18));
    LocalMux I__7075 (
            .O(N__36316),
            .I(sRAM_pointer_writeZ0Z_18));
    CascadeMux I__7074 (
            .O(N__36311),
            .I(N__36308));
    InMux I__7073 (
            .O(N__36308),
            .I(N__36305));
    LocalMux I__7072 (
            .O(N__36305),
            .I(N__36302));
    Span12Mux_h I__7071 (
            .O(N__36302),
            .I(N__36298));
    InMux I__7070 (
            .O(N__36301),
            .I(N__36295));
    Odrv12 I__7069 (
            .O(N__36298),
            .I(sRAM_pointer_readZ0Z_18));
    LocalMux I__7068 (
            .O(N__36295),
            .I(sRAM_pointer_readZ0Z_18));
    IoInMux I__7067 (
            .O(N__36290),
            .I(N__36287));
    LocalMux I__7066 (
            .O(N__36287),
            .I(N__36284));
    IoSpan4Mux I__7065 (
            .O(N__36284),
            .I(N__36281));
    Span4Mux_s1_h I__7064 (
            .O(N__36281),
            .I(N__36278));
    Sp12to4 I__7063 (
            .O(N__36278),
            .I(N__36275));
    Span12Mux_h I__7062 (
            .O(N__36275),
            .I(N__36272));
    Span12Mux_v I__7061 (
            .O(N__36272),
            .I(N__36269));
    Odrv12 I__7060 (
            .O(N__36269),
            .I(RAM_ADD_c_18));
    InMux I__7059 (
            .O(N__36266),
            .I(N__36263));
    LocalMux I__7058 (
            .O(N__36263),
            .I(N__36260));
    Span4Mux_v I__7057 (
            .O(N__36260),
            .I(N__36257));
    Span4Mux_h I__7056 (
            .O(N__36257),
            .I(N__36254));
    Sp12to4 I__7055 (
            .O(N__36254),
            .I(N__36251));
    Span12Mux_h I__7054 (
            .O(N__36251),
            .I(N__36247));
    InMux I__7053 (
            .O(N__36250),
            .I(N__36244));
    Odrv12 I__7052 (
            .O(N__36247),
            .I(sRAM_pointer_writeZ0Z_9));
    LocalMux I__7051 (
            .O(N__36244),
            .I(sRAM_pointer_writeZ0Z_9));
    CascadeMux I__7050 (
            .O(N__36239),
            .I(N__36236));
    InMux I__7049 (
            .O(N__36236),
            .I(N__36233));
    LocalMux I__7048 (
            .O(N__36233),
            .I(N__36230));
    Span4Mux_v I__7047 (
            .O(N__36230),
            .I(N__36226));
    InMux I__7046 (
            .O(N__36229),
            .I(N__36223));
    Odrv4 I__7045 (
            .O(N__36226),
            .I(sRAM_pointer_readZ0Z_9));
    LocalMux I__7044 (
            .O(N__36223),
            .I(sRAM_pointer_readZ0Z_9));
    IoInMux I__7043 (
            .O(N__36218),
            .I(N__36215));
    LocalMux I__7042 (
            .O(N__36215),
            .I(N__36212));
    Span4Mux_s3_h I__7041 (
            .O(N__36212),
            .I(N__36209));
    Span4Mux_h I__7040 (
            .O(N__36209),
            .I(N__36206));
    Span4Mux_h I__7039 (
            .O(N__36206),
            .I(N__36203));
    Span4Mux_v I__7038 (
            .O(N__36203),
            .I(N__36200));
    Odrv4 I__7037 (
            .O(N__36200),
            .I(RAM_ADD_c_9));
    InMux I__7036 (
            .O(N__36197),
            .I(N__36194));
    LocalMux I__7035 (
            .O(N__36194),
            .I(N__36191));
    Span4Mux_h I__7034 (
            .O(N__36191),
            .I(N__36188));
    Span4Mux_h I__7033 (
            .O(N__36188),
            .I(N__36185));
    Sp12to4 I__7032 (
            .O(N__36185),
            .I(N__36182));
    Span12Mux_v I__7031 (
            .O(N__36182),
            .I(N__36178));
    InMux I__7030 (
            .O(N__36181),
            .I(N__36175));
    Odrv12 I__7029 (
            .O(N__36178),
            .I(sRAM_pointer_writeZ0Z_7));
    LocalMux I__7028 (
            .O(N__36175),
            .I(sRAM_pointer_writeZ0Z_7));
    CascadeMux I__7027 (
            .O(N__36170),
            .I(N__36167));
    InMux I__7026 (
            .O(N__36167),
            .I(N__36164));
    LocalMux I__7025 (
            .O(N__36164),
            .I(N__36160));
    InMux I__7024 (
            .O(N__36163),
            .I(N__36157));
    Odrv12 I__7023 (
            .O(N__36160),
            .I(sRAM_pointer_readZ0Z_7));
    LocalMux I__7022 (
            .O(N__36157),
            .I(sRAM_pointer_readZ0Z_7));
    IoInMux I__7021 (
            .O(N__36152),
            .I(N__36149));
    LocalMux I__7020 (
            .O(N__36149),
            .I(N__36146));
    Span4Mux_s0_h I__7019 (
            .O(N__36146),
            .I(N__36143));
    Sp12to4 I__7018 (
            .O(N__36143),
            .I(N__36140));
    Span12Mux_s8_v I__7017 (
            .O(N__36140),
            .I(N__36137));
    Odrv12 I__7016 (
            .O(N__36137),
            .I(RAM_ADD_c_7));
    InMux I__7015 (
            .O(N__36134),
            .I(N__36131));
    LocalMux I__7014 (
            .O(N__36131),
            .I(N__36127));
    InMux I__7013 (
            .O(N__36130),
            .I(N__36124));
    Odrv4 I__7012 (
            .O(N__36127),
            .I(sRAM_pointer_readZ0Z_2));
    LocalMux I__7011 (
            .O(N__36124),
            .I(sRAM_pointer_readZ0Z_2));
    CascadeMux I__7010 (
            .O(N__36119),
            .I(N__36116));
    InMux I__7009 (
            .O(N__36116),
            .I(N__36113));
    LocalMux I__7008 (
            .O(N__36113),
            .I(N__36110));
    Span4Mux_v I__7007 (
            .O(N__36110),
            .I(N__36107));
    Span4Mux_h I__7006 (
            .O(N__36107),
            .I(N__36104));
    Sp12to4 I__7005 (
            .O(N__36104),
            .I(N__36101));
    Span12Mux_h I__7004 (
            .O(N__36101),
            .I(N__36097));
    InMux I__7003 (
            .O(N__36100),
            .I(N__36094));
    Odrv12 I__7002 (
            .O(N__36097),
            .I(sRAM_pointer_writeZ0Z_2));
    LocalMux I__7001 (
            .O(N__36094),
            .I(sRAM_pointer_writeZ0Z_2));
    IoInMux I__7000 (
            .O(N__36089),
            .I(N__36086));
    LocalMux I__6999 (
            .O(N__36086),
            .I(N__36083));
    Span4Mux_s2_v I__6998 (
            .O(N__36083),
            .I(N__36080));
    Span4Mux_v I__6997 (
            .O(N__36080),
            .I(N__36077));
    Odrv4 I__6996 (
            .O(N__36077),
            .I(RAM_ADD_c_2));
    InMux I__6995 (
            .O(N__36074),
            .I(N__36071));
    LocalMux I__6994 (
            .O(N__36071),
            .I(N__36068));
    Span4Mux_v I__6993 (
            .O(N__36068),
            .I(N__36065));
    Span4Mux_h I__6992 (
            .O(N__36065),
            .I(N__36062));
    Sp12to4 I__6991 (
            .O(N__36062),
            .I(N__36059));
    Span12Mux_h I__6990 (
            .O(N__36059),
            .I(N__36055));
    InMux I__6989 (
            .O(N__36058),
            .I(N__36052));
    Odrv12 I__6988 (
            .O(N__36055),
            .I(sRAM_pointer_writeZ0Z_1));
    LocalMux I__6987 (
            .O(N__36052),
            .I(sRAM_pointer_writeZ0Z_1));
    CascadeMux I__6986 (
            .O(N__36047),
            .I(N__36044));
    InMux I__6985 (
            .O(N__36044),
            .I(N__36041));
    LocalMux I__6984 (
            .O(N__36041),
            .I(N__36037));
    InMux I__6983 (
            .O(N__36040),
            .I(N__36034));
    Odrv4 I__6982 (
            .O(N__36037),
            .I(sRAM_pointer_readZ0Z_1));
    LocalMux I__6981 (
            .O(N__36034),
            .I(sRAM_pointer_readZ0Z_1));
    IoInMux I__6980 (
            .O(N__36029),
            .I(N__36026));
    LocalMux I__6979 (
            .O(N__36026),
            .I(N__36023));
    Span12Mux_s2_v I__6978 (
            .O(N__36023),
            .I(N__36020));
    Odrv12 I__6977 (
            .O(N__36020),
            .I(RAM_ADD_c_1));
    InMux I__6976 (
            .O(N__36017),
            .I(N__36014));
    LocalMux I__6975 (
            .O(N__36014),
            .I(N__36011));
    Span4Mux_v I__6974 (
            .O(N__36011),
            .I(N__36008));
    Span4Mux_h I__6973 (
            .O(N__36008),
            .I(N__36005));
    Span4Mux_v I__6972 (
            .O(N__36005),
            .I(N__36002));
    Sp12to4 I__6971 (
            .O(N__36002),
            .I(N__35998));
    InMux I__6970 (
            .O(N__36001),
            .I(N__35995));
    Odrv12 I__6969 (
            .O(N__35998),
            .I(sRAM_pointer_writeZ0Z_6));
    LocalMux I__6968 (
            .O(N__35995),
            .I(sRAM_pointer_writeZ0Z_6));
    CascadeMux I__6967 (
            .O(N__35990),
            .I(N__35987));
    InMux I__6966 (
            .O(N__35987),
            .I(N__35984));
    LocalMux I__6965 (
            .O(N__35984),
            .I(N__35980));
    InMux I__6964 (
            .O(N__35983),
            .I(N__35977));
    Odrv12 I__6963 (
            .O(N__35980),
            .I(sRAM_pointer_readZ0Z_6));
    LocalMux I__6962 (
            .O(N__35977),
            .I(sRAM_pointer_readZ0Z_6));
    IoInMux I__6961 (
            .O(N__35972),
            .I(N__35969));
    LocalMux I__6960 (
            .O(N__35969),
            .I(N__35966));
    IoSpan4Mux I__6959 (
            .O(N__35966),
            .I(N__35963));
    Span4Mux_s3_h I__6958 (
            .O(N__35963),
            .I(N__35960));
    Span4Mux_h I__6957 (
            .O(N__35960),
            .I(N__35957));
    Span4Mux_h I__6956 (
            .O(N__35957),
            .I(N__35954));
    Odrv4 I__6955 (
            .O(N__35954),
            .I(RAM_ADD_c_6));
    InMux I__6954 (
            .O(N__35951),
            .I(N__35948));
    LocalMux I__6953 (
            .O(N__35948),
            .I(N__35945));
    Span4Mux_v I__6952 (
            .O(N__35945),
            .I(N__35942));
    Span4Mux_h I__6951 (
            .O(N__35942),
            .I(N__35939));
    Sp12to4 I__6950 (
            .O(N__35939),
            .I(N__35936));
    Span12Mux_h I__6949 (
            .O(N__35936),
            .I(N__35933));
    Odrv12 I__6948 (
            .O(N__35933),
            .I(ADC4_c));
    IoInMux I__6947 (
            .O(N__35930),
            .I(N__35927));
    LocalMux I__6946 (
            .O(N__35927),
            .I(N__35924));
    Span4Mux_s2_v I__6945 (
            .O(N__35924),
            .I(N__35921));
    Span4Mux_h I__6944 (
            .O(N__35921),
            .I(N__35918));
    Span4Mux_h I__6943 (
            .O(N__35918),
            .I(N__35915));
    Span4Mux_v I__6942 (
            .O(N__35915),
            .I(N__35912));
    Odrv4 I__6941 (
            .O(N__35912),
            .I(RAM_DATA_1Z0Z_4));
    InMux I__6940 (
            .O(N__35909),
            .I(N__35906));
    LocalMux I__6939 (
            .O(N__35906),
            .I(N__35903));
    Span4Mux_v I__6938 (
            .O(N__35903),
            .I(N__35899));
    InMux I__6937 (
            .O(N__35902),
            .I(N__35896));
    Odrv4 I__6936 (
            .O(N__35899),
            .I(sRAM_pointer_readZ0Z_0));
    LocalMux I__6935 (
            .O(N__35896),
            .I(sRAM_pointer_readZ0Z_0));
    CascadeMux I__6934 (
            .O(N__35891),
            .I(N__35888));
    InMux I__6933 (
            .O(N__35888),
            .I(N__35885));
    LocalMux I__6932 (
            .O(N__35885),
            .I(N__35882));
    Span4Mux_h I__6931 (
            .O(N__35882),
            .I(N__35879));
    Sp12to4 I__6930 (
            .O(N__35879),
            .I(N__35876));
    Span12Mux_s7_v I__6929 (
            .O(N__35876),
            .I(N__35873));
    Span12Mux_h I__6928 (
            .O(N__35873),
            .I(N__35869));
    InMux I__6927 (
            .O(N__35872),
            .I(N__35866));
    Odrv12 I__6926 (
            .O(N__35869),
            .I(sRAM_pointer_writeZ0Z_0));
    LocalMux I__6925 (
            .O(N__35866),
            .I(sRAM_pointer_writeZ0Z_0));
    IoInMux I__6924 (
            .O(N__35861),
            .I(N__35858));
    LocalMux I__6923 (
            .O(N__35858),
            .I(N__35855));
    IoSpan4Mux I__6922 (
            .O(N__35855),
            .I(N__35852));
    Sp12to4 I__6921 (
            .O(N__35852),
            .I(N__35849));
    Odrv12 I__6920 (
            .O(N__35849),
            .I(RAM_ADD_c_0));
    InMux I__6919 (
            .O(N__35846),
            .I(N__35843));
    LocalMux I__6918 (
            .O(N__35843),
            .I(N__35840));
    Span4Mux_v I__6917 (
            .O(N__35840),
            .I(N__35836));
    InMux I__6916 (
            .O(N__35839),
            .I(N__35833));
    Odrv4 I__6915 (
            .O(N__35836),
            .I(sRAM_pointer_readZ0Z_10));
    LocalMux I__6914 (
            .O(N__35833),
            .I(sRAM_pointer_readZ0Z_10));
    InMux I__6913 (
            .O(N__35828),
            .I(N__35825));
    LocalMux I__6912 (
            .O(N__35825),
            .I(N__35822));
    Span4Mux_v I__6911 (
            .O(N__35822),
            .I(N__35819));
    Span4Mux_h I__6910 (
            .O(N__35819),
            .I(N__35816));
    Span4Mux_h I__6909 (
            .O(N__35816),
            .I(N__35813));
    Span4Mux_h I__6908 (
            .O(N__35813),
            .I(N__35810));
    Span4Mux_h I__6907 (
            .O(N__35810),
            .I(N__35806));
    InMux I__6906 (
            .O(N__35809),
            .I(N__35803));
    Odrv4 I__6905 (
            .O(N__35806),
            .I(sRAM_pointer_writeZ0Z_10));
    LocalMux I__6904 (
            .O(N__35803),
            .I(sRAM_pointer_writeZ0Z_10));
    IoInMux I__6903 (
            .O(N__35798),
            .I(N__35795));
    LocalMux I__6902 (
            .O(N__35795),
            .I(N__35792));
    IoSpan4Mux I__6901 (
            .O(N__35792),
            .I(N__35789));
    Span4Mux_s1_h I__6900 (
            .O(N__35789),
            .I(N__35786));
    Sp12to4 I__6899 (
            .O(N__35786),
            .I(N__35783));
    Span12Mux_h I__6898 (
            .O(N__35783),
            .I(N__35780));
    Span12Mux_v I__6897 (
            .O(N__35780),
            .I(N__35777));
    Odrv12 I__6896 (
            .O(N__35777),
            .I(RAM_ADD_c_10));
    InMux I__6895 (
            .O(N__35774),
            .I(N__35771));
    LocalMux I__6894 (
            .O(N__35771),
            .I(N__35768));
    Span4Mux_v I__6893 (
            .O(N__35768),
            .I(N__35764));
    InMux I__6892 (
            .O(N__35767),
            .I(N__35761));
    Odrv4 I__6891 (
            .O(N__35764),
            .I(sRAM_pointer_readZ0Z_11));
    LocalMux I__6890 (
            .O(N__35761),
            .I(sRAM_pointer_readZ0Z_11));
    CascadeMux I__6889 (
            .O(N__35756),
            .I(N__35753));
    InMux I__6888 (
            .O(N__35753),
            .I(N__35750));
    LocalMux I__6887 (
            .O(N__35750),
            .I(N__35747));
    Span4Mux_v I__6886 (
            .O(N__35747),
            .I(N__35744));
    Span4Mux_h I__6885 (
            .O(N__35744),
            .I(N__35741));
    Sp12to4 I__6884 (
            .O(N__35741),
            .I(N__35738));
    Span12Mux_h I__6883 (
            .O(N__35738),
            .I(N__35734));
    InMux I__6882 (
            .O(N__35737),
            .I(N__35731));
    Odrv12 I__6881 (
            .O(N__35734),
            .I(sRAM_pointer_writeZ0Z_11));
    LocalMux I__6880 (
            .O(N__35731),
            .I(sRAM_pointer_writeZ0Z_11));
    IoInMux I__6879 (
            .O(N__35726),
            .I(N__35723));
    LocalMux I__6878 (
            .O(N__35723),
            .I(N__35720));
    Span4Mux_s0_h I__6877 (
            .O(N__35720),
            .I(N__35717));
    Sp12to4 I__6876 (
            .O(N__35717),
            .I(N__35714));
    Span12Mux_v I__6875 (
            .O(N__35714),
            .I(N__35711));
    Span12Mux_h I__6874 (
            .O(N__35711),
            .I(N__35708));
    Odrv12 I__6873 (
            .O(N__35708),
            .I(RAM_ADD_c_11));
    InMux I__6872 (
            .O(N__35705),
            .I(N__35702));
    LocalMux I__6871 (
            .O(N__35702),
            .I(N__35699));
    Span4Mux_v I__6870 (
            .O(N__35699),
            .I(N__35696));
    Span4Mux_h I__6869 (
            .O(N__35696),
            .I(N__35693));
    Sp12to4 I__6868 (
            .O(N__35693),
            .I(N__35690));
    Span12Mux_v I__6867 (
            .O(N__35690),
            .I(N__35686));
    InMux I__6866 (
            .O(N__35689),
            .I(N__35683));
    Odrv12 I__6865 (
            .O(N__35686),
            .I(sRAM_pointer_writeZ0Z_12));
    LocalMux I__6864 (
            .O(N__35683),
            .I(sRAM_pointer_writeZ0Z_12));
    InMux I__6863 (
            .O(N__35678),
            .I(N__35675));
    LocalMux I__6862 (
            .O(N__35675),
            .I(N__35672));
    Span4Mux_v I__6861 (
            .O(N__35672),
            .I(N__35668));
    InMux I__6860 (
            .O(N__35671),
            .I(N__35665));
    Odrv4 I__6859 (
            .O(N__35668),
            .I(sRAM_pointer_readZ0Z_12));
    LocalMux I__6858 (
            .O(N__35665),
            .I(sRAM_pointer_readZ0Z_12));
    IoInMux I__6857 (
            .O(N__35660),
            .I(N__35657));
    LocalMux I__6856 (
            .O(N__35657),
            .I(N__35654));
    Span4Mux_s0_h I__6855 (
            .O(N__35654),
            .I(N__35651));
    Sp12to4 I__6854 (
            .O(N__35651),
            .I(N__35648));
    Span12Mux_v I__6853 (
            .O(N__35648),
            .I(N__35645));
    Span12Mux_h I__6852 (
            .O(N__35645),
            .I(N__35642));
    Odrv12 I__6851 (
            .O(N__35642),
            .I(RAM_ADD_c_12));
    InMux I__6850 (
            .O(N__35639),
            .I(N__35636));
    LocalMux I__6849 (
            .O(N__35636),
            .I(N__35633));
    Span4Mux_h I__6848 (
            .O(N__35633),
            .I(N__35629));
    InMux I__6847 (
            .O(N__35632),
            .I(N__35626));
    Odrv4 I__6846 (
            .O(N__35629),
            .I(sRAM_pointer_readZ0Z_13));
    LocalMux I__6845 (
            .O(N__35626),
            .I(sRAM_pointer_readZ0Z_13));
    CascadeMux I__6844 (
            .O(N__35621),
            .I(N__35618));
    InMux I__6843 (
            .O(N__35618),
            .I(N__35615));
    LocalMux I__6842 (
            .O(N__35615),
            .I(N__35612));
    Span4Mux_h I__6841 (
            .O(N__35612),
            .I(N__35609));
    Sp12to4 I__6840 (
            .O(N__35609),
            .I(N__35606));
    Span12Mux_h I__6839 (
            .O(N__35606),
            .I(N__35602));
    InMux I__6838 (
            .O(N__35605),
            .I(N__35599));
    Odrv12 I__6837 (
            .O(N__35602),
            .I(sRAM_pointer_writeZ0Z_13));
    LocalMux I__6836 (
            .O(N__35599),
            .I(sRAM_pointer_writeZ0Z_13));
    IoInMux I__6835 (
            .O(N__35594),
            .I(N__35591));
    LocalMux I__6834 (
            .O(N__35591),
            .I(N__35588));
    Sp12to4 I__6833 (
            .O(N__35588),
            .I(N__35585));
    Span12Mux_h I__6832 (
            .O(N__35585),
            .I(N__35582));
    Span12Mux_v I__6831 (
            .O(N__35582),
            .I(N__35579));
    Odrv12 I__6830 (
            .O(N__35579),
            .I(RAM_ADD_c_13));
    InMux I__6829 (
            .O(N__35576),
            .I(N__35573));
    LocalMux I__6828 (
            .O(N__35573),
            .I(N__35570));
    Span4Mux_v I__6827 (
            .O(N__35570),
            .I(N__35567));
    Span4Mux_h I__6826 (
            .O(N__35567),
            .I(N__35564));
    Sp12to4 I__6825 (
            .O(N__35564),
            .I(N__35561));
    Span12Mux_h I__6824 (
            .O(N__35561),
            .I(N__35557));
    InMux I__6823 (
            .O(N__35560),
            .I(N__35554));
    Odrv12 I__6822 (
            .O(N__35557),
            .I(sRAM_pointer_writeZ0Z_14));
    LocalMux I__6821 (
            .O(N__35554),
            .I(sRAM_pointer_writeZ0Z_14));
    InMux I__6820 (
            .O(N__35549),
            .I(N__35546));
    LocalMux I__6819 (
            .O(N__35546),
            .I(N__35543));
    Span4Mux_h I__6818 (
            .O(N__35543),
            .I(N__35540));
    Span4Mux_h I__6817 (
            .O(N__35540),
            .I(N__35536));
    InMux I__6816 (
            .O(N__35539),
            .I(N__35533));
    Odrv4 I__6815 (
            .O(N__35536),
            .I(sRAM_pointer_readZ0Z_14));
    LocalMux I__6814 (
            .O(N__35533),
            .I(sRAM_pointer_readZ0Z_14));
    IoInMux I__6813 (
            .O(N__35528),
            .I(N__35525));
    LocalMux I__6812 (
            .O(N__35525),
            .I(N__35522));
    IoSpan4Mux I__6811 (
            .O(N__35522),
            .I(N__35519));
    Span4Mux_s1_h I__6810 (
            .O(N__35519),
            .I(N__35516));
    Sp12to4 I__6809 (
            .O(N__35516),
            .I(N__35513));
    Span12Mux_h I__6808 (
            .O(N__35513),
            .I(N__35510));
    Span12Mux_v I__6807 (
            .O(N__35510),
            .I(N__35507));
    Odrv12 I__6806 (
            .O(N__35507),
            .I(RAM_ADD_c_14));
    InMux I__6805 (
            .O(N__35504),
            .I(N__35501));
    LocalMux I__6804 (
            .O(N__35501),
            .I(N__35498));
    Span4Mux_h I__6803 (
            .O(N__35498),
            .I(N__35494));
    InMux I__6802 (
            .O(N__35497),
            .I(N__35491));
    Odrv4 I__6801 (
            .O(N__35494),
            .I(sRAM_pointer_readZ0Z_15));
    LocalMux I__6800 (
            .O(N__35491),
            .I(sRAM_pointer_readZ0Z_15));
    CascadeMux I__6799 (
            .O(N__35486),
            .I(N__35483));
    InMux I__6798 (
            .O(N__35483),
            .I(N__35480));
    LocalMux I__6797 (
            .O(N__35480),
            .I(N__35477));
    Span4Mux_v I__6796 (
            .O(N__35477),
            .I(N__35474));
    Span4Mux_h I__6795 (
            .O(N__35474),
            .I(N__35471));
    Span4Mux_h I__6794 (
            .O(N__35471),
            .I(N__35468));
    Sp12to4 I__6793 (
            .O(N__35468),
            .I(N__35465));
    Span12Mux_h I__6792 (
            .O(N__35465),
            .I(N__35461));
    InMux I__6791 (
            .O(N__35464),
            .I(N__35458));
    Odrv12 I__6790 (
            .O(N__35461),
            .I(sRAM_pointer_writeZ0Z_15));
    LocalMux I__6789 (
            .O(N__35458),
            .I(sRAM_pointer_writeZ0Z_15));
    IoInMux I__6788 (
            .O(N__35453),
            .I(N__35450));
    LocalMux I__6787 (
            .O(N__35450),
            .I(N__35447));
    IoSpan4Mux I__6786 (
            .O(N__35447),
            .I(N__35444));
    Span4Mux_s2_h I__6785 (
            .O(N__35444),
            .I(N__35441));
    Span4Mux_h I__6784 (
            .O(N__35441),
            .I(N__35438));
    Span4Mux_h I__6783 (
            .O(N__35438),
            .I(N__35435));
    Odrv4 I__6782 (
            .O(N__35435),
            .I(RAM_ADD_c_15));
    InMux I__6781 (
            .O(N__35432),
            .I(N__35429));
    LocalMux I__6780 (
            .O(N__35429),
            .I(N__35426));
    Span4Mux_h I__6779 (
            .O(N__35426),
            .I(N__35422));
    InMux I__6778 (
            .O(N__35425),
            .I(N__35419));
    Odrv4 I__6777 (
            .O(N__35422),
            .I(sRAM_pointer_readZ0Z_16));
    LocalMux I__6776 (
            .O(N__35419),
            .I(sRAM_pointer_readZ0Z_16));
    CascadeMux I__6775 (
            .O(N__35414),
            .I(N__35411));
    InMux I__6774 (
            .O(N__35411),
            .I(N__35408));
    LocalMux I__6773 (
            .O(N__35408),
            .I(N__35405));
    Span4Mux_v I__6772 (
            .O(N__35405),
            .I(N__35402));
    Span4Mux_h I__6771 (
            .O(N__35402),
            .I(N__35399));
    Span4Mux_h I__6770 (
            .O(N__35399),
            .I(N__35396));
    Span4Mux_h I__6769 (
            .O(N__35396),
            .I(N__35392));
    InMux I__6768 (
            .O(N__35395),
            .I(N__35389));
    Span4Mux_h I__6767 (
            .O(N__35392),
            .I(N__35386));
    LocalMux I__6766 (
            .O(N__35389),
            .I(sRAM_pointer_writeZ0Z_16));
    Odrv4 I__6765 (
            .O(N__35386),
            .I(sRAM_pointer_writeZ0Z_16));
    IoInMux I__6764 (
            .O(N__35381),
            .I(N__35378));
    LocalMux I__6763 (
            .O(N__35378),
            .I(N__35375));
    IoSpan4Mux I__6762 (
            .O(N__35375),
            .I(N__35372));
    Span4Mux_s1_h I__6761 (
            .O(N__35372),
            .I(N__35369));
    Span4Mux_h I__6760 (
            .O(N__35369),
            .I(N__35366));
    Span4Mux_h I__6759 (
            .O(N__35366),
            .I(N__35363));
    Odrv4 I__6758 (
            .O(N__35363),
            .I(RAM_ADD_c_16));
    InMux I__6757 (
            .O(N__35360),
            .I(N__35356));
    InMux I__6756 (
            .O(N__35359),
            .I(N__35353));
    LocalMux I__6755 (
            .O(N__35356),
            .I(button_debounce_counterZ0Z_19));
    LocalMux I__6754 (
            .O(N__35353),
            .I(button_debounce_counterZ0Z_19));
    InMux I__6753 (
            .O(N__35348),
            .I(un1_button_debounce_counter_cry_18));
    InMux I__6752 (
            .O(N__35345),
            .I(N__35341));
    InMux I__6751 (
            .O(N__35344),
            .I(N__35338));
    LocalMux I__6750 (
            .O(N__35341),
            .I(button_debounce_counterZ0Z_20));
    LocalMux I__6749 (
            .O(N__35338),
            .I(button_debounce_counterZ0Z_20));
    InMux I__6748 (
            .O(N__35333),
            .I(un1_button_debounce_counter_cry_19));
    CascadeMux I__6747 (
            .O(N__35330),
            .I(N__35326));
    InMux I__6746 (
            .O(N__35329),
            .I(N__35323));
    InMux I__6745 (
            .O(N__35326),
            .I(N__35320));
    LocalMux I__6744 (
            .O(N__35323),
            .I(button_debounce_counterZ0Z_21));
    LocalMux I__6743 (
            .O(N__35320),
            .I(button_debounce_counterZ0Z_21));
    InMux I__6742 (
            .O(N__35315),
            .I(un1_button_debounce_counter_cry_20));
    InMux I__6741 (
            .O(N__35312),
            .I(N__35309));
    LocalMux I__6740 (
            .O(N__35309),
            .I(N__35306));
    Span4Mux_v I__6739 (
            .O(N__35306),
            .I(N__35302));
    InMux I__6738 (
            .O(N__35305),
            .I(N__35299));
    Span4Mux_h I__6737 (
            .O(N__35302),
            .I(N__35296));
    LocalMux I__6736 (
            .O(N__35299),
            .I(button_debounce_counterZ0Z_22));
    Odrv4 I__6735 (
            .O(N__35296),
            .I(button_debounce_counterZ0Z_22));
    InMux I__6734 (
            .O(N__35291),
            .I(un1_button_debounce_counter_cry_21));
    InMux I__6733 (
            .O(N__35288),
            .I(bfn_16_16_0_));
    CascadeMux I__6732 (
            .O(N__35285),
            .I(N__35281));
    InMux I__6731 (
            .O(N__35284),
            .I(N__35278));
    InMux I__6730 (
            .O(N__35281),
            .I(N__35275));
    LocalMux I__6729 (
            .O(N__35278),
            .I(button_debounce_counterZ0Z_23));
    LocalMux I__6728 (
            .O(N__35275),
            .I(button_debounce_counterZ0Z_23));
    CEMux I__6727 (
            .O(N__35270),
            .I(N__35267));
    LocalMux I__6726 (
            .O(N__35267),
            .I(N__35264));
    Span4Mux_h I__6725 (
            .O(N__35264),
            .I(N__35261));
    Span4Mux_v I__6724 (
            .O(N__35261),
            .I(N__35258));
    Odrv4 I__6723 (
            .O(N__35258),
            .I(LED3_c_0));
    InMux I__6722 (
            .O(N__35255),
            .I(N__35252));
    LocalMux I__6721 (
            .O(N__35252),
            .I(N__35249));
    Span4Mux_h I__6720 (
            .O(N__35249),
            .I(N__35245));
    InMux I__6719 (
            .O(N__35248),
            .I(N__35242));
    Odrv4 I__6718 (
            .O(N__35245),
            .I(sRAM_pointer_readZ0Z_5));
    LocalMux I__6717 (
            .O(N__35242),
            .I(sRAM_pointer_readZ0Z_5));
    InMux I__6716 (
            .O(N__35237),
            .I(N__35234));
    LocalMux I__6715 (
            .O(N__35234),
            .I(N__35231));
    Span12Mux_v I__6714 (
            .O(N__35231),
            .I(N__35228));
    Span12Mux_h I__6713 (
            .O(N__35228),
            .I(N__35224));
    InMux I__6712 (
            .O(N__35227),
            .I(N__35221));
    Odrv12 I__6711 (
            .O(N__35224),
            .I(sRAM_pointer_writeZ0Z_5));
    LocalMux I__6710 (
            .O(N__35221),
            .I(sRAM_pointer_writeZ0Z_5));
    IoInMux I__6709 (
            .O(N__35216),
            .I(N__35213));
    LocalMux I__6708 (
            .O(N__35213),
            .I(N__35210));
    Span4Mux_s3_h I__6707 (
            .O(N__35210),
            .I(N__35207));
    Span4Mux_h I__6706 (
            .O(N__35207),
            .I(N__35204));
    Span4Mux_h I__6705 (
            .O(N__35204),
            .I(N__35201));
    Span4Mux_v I__6704 (
            .O(N__35201),
            .I(N__35198));
    Odrv4 I__6703 (
            .O(N__35198),
            .I(RAM_ADD_c_5));
    InMux I__6702 (
            .O(N__35195),
            .I(un1_button_debounce_counter_cry_9));
    InMux I__6701 (
            .O(N__35192),
            .I(un1_button_debounce_counter_cry_10));
    InMux I__6700 (
            .O(N__35189),
            .I(un1_button_debounce_counter_cry_11));
    InMux I__6699 (
            .O(N__35186),
            .I(un1_button_debounce_counter_cry_12));
    InMux I__6698 (
            .O(N__35183),
            .I(un1_button_debounce_counter_cry_13));
    InMux I__6697 (
            .O(N__35180),
            .I(N__35176));
    InMux I__6696 (
            .O(N__35179),
            .I(N__35173));
    LocalMux I__6695 (
            .O(N__35176),
            .I(N__35170));
    LocalMux I__6694 (
            .O(N__35173),
            .I(button_debounce_counterZ0Z_15));
    Odrv4 I__6693 (
            .O(N__35170),
            .I(button_debounce_counterZ0Z_15));
    InMux I__6692 (
            .O(N__35165),
            .I(un1_button_debounce_counter_cry_14));
    InMux I__6691 (
            .O(N__35162),
            .I(N__35159));
    LocalMux I__6690 (
            .O(N__35159),
            .I(N__35155));
    InMux I__6689 (
            .O(N__35158),
            .I(N__35152));
    Span4Mux_h I__6688 (
            .O(N__35155),
            .I(N__35149));
    LocalMux I__6687 (
            .O(N__35152),
            .I(button_debounce_counterZ0Z_16));
    Odrv4 I__6686 (
            .O(N__35149),
            .I(button_debounce_counterZ0Z_16));
    InMux I__6685 (
            .O(N__35144),
            .I(un1_button_debounce_counter_cry_15));
    InMux I__6684 (
            .O(N__35141),
            .I(N__35137));
    InMux I__6683 (
            .O(N__35140),
            .I(N__35134));
    LocalMux I__6682 (
            .O(N__35137),
            .I(N__35131));
    LocalMux I__6681 (
            .O(N__35134),
            .I(button_debounce_counterZ0Z_17));
    Odrv4 I__6680 (
            .O(N__35131),
            .I(button_debounce_counterZ0Z_17));
    InMux I__6679 (
            .O(N__35126),
            .I(bfn_16_15_0_));
    InMux I__6678 (
            .O(N__35123),
            .I(N__35119));
    InMux I__6677 (
            .O(N__35122),
            .I(N__35116));
    LocalMux I__6676 (
            .O(N__35119),
            .I(button_debounce_counterZ0Z_18));
    LocalMux I__6675 (
            .O(N__35116),
            .I(button_debounce_counterZ0Z_18));
    InMux I__6674 (
            .O(N__35111),
            .I(un1_button_debounce_counter_cry_17));
    CascadeMux I__6673 (
            .O(N__35108),
            .I(N__35105));
    InMux I__6672 (
            .O(N__35105),
            .I(N__35102));
    LocalMux I__6671 (
            .O(N__35102),
            .I(N__35098));
    InMux I__6670 (
            .O(N__35101),
            .I(N__35095));
    Odrv12 I__6669 (
            .O(N__35098),
            .I(button_debounce_counterZ0Z_2));
    LocalMux I__6668 (
            .O(N__35095),
            .I(button_debounce_counterZ0Z_2));
    InMux I__6667 (
            .O(N__35090),
            .I(un1_button_debounce_counter_cry_1));
    InMux I__6666 (
            .O(N__35087),
            .I(N__35083));
    InMux I__6665 (
            .O(N__35086),
            .I(N__35080));
    LocalMux I__6664 (
            .O(N__35083),
            .I(button_debounce_counterZ0Z_3));
    LocalMux I__6663 (
            .O(N__35080),
            .I(button_debounce_counterZ0Z_3));
    InMux I__6662 (
            .O(N__35075),
            .I(un1_button_debounce_counter_cry_2));
    InMux I__6661 (
            .O(N__35072),
            .I(N__35068));
    InMux I__6660 (
            .O(N__35071),
            .I(N__35065));
    LocalMux I__6659 (
            .O(N__35068),
            .I(button_debounce_counterZ0Z_4));
    LocalMux I__6658 (
            .O(N__35065),
            .I(button_debounce_counterZ0Z_4));
    InMux I__6657 (
            .O(N__35060),
            .I(un1_button_debounce_counter_cry_3));
    CascadeMux I__6656 (
            .O(N__35057),
            .I(N__35054));
    InMux I__6655 (
            .O(N__35054),
            .I(N__35050));
    InMux I__6654 (
            .O(N__35053),
            .I(N__35047));
    LocalMux I__6653 (
            .O(N__35050),
            .I(button_debounce_counterZ0Z_5));
    LocalMux I__6652 (
            .O(N__35047),
            .I(button_debounce_counterZ0Z_5));
    InMux I__6651 (
            .O(N__35042),
            .I(un1_button_debounce_counter_cry_4));
    InMux I__6650 (
            .O(N__35039),
            .I(N__35036));
    LocalMux I__6649 (
            .O(N__35036),
            .I(N__35032));
    InMux I__6648 (
            .O(N__35035),
            .I(N__35029));
    Odrv4 I__6647 (
            .O(N__35032),
            .I(button_debounce_counterZ0Z_6));
    LocalMux I__6646 (
            .O(N__35029),
            .I(button_debounce_counterZ0Z_6));
    InMux I__6645 (
            .O(N__35024),
            .I(un1_button_debounce_counter_cry_5));
    InMux I__6644 (
            .O(N__35021),
            .I(un1_button_debounce_counter_cry_6));
    InMux I__6643 (
            .O(N__35018),
            .I(un1_button_debounce_counter_cry_7));
    InMux I__6642 (
            .O(N__35015),
            .I(bfn_16_14_0_));
    InMux I__6641 (
            .O(N__35012),
            .I(N__35009));
    LocalMux I__6640 (
            .O(N__35009),
            .I(N__35006));
    Span4Mux_h I__6639 (
            .O(N__35006),
            .I(N__35003));
    Span4Mux_v I__6638 (
            .O(N__35003),
            .I(N__35000));
    Odrv4 I__6637 (
            .O(N__35000),
            .I(sDAC_mem_19Z0Z_3));
    CEMux I__6636 (
            .O(N__34997),
            .I(N__34994));
    LocalMux I__6635 (
            .O(N__34994),
            .I(N__34991));
    Span4Mux_v I__6634 (
            .O(N__34991),
            .I(N__34987));
    CEMux I__6633 (
            .O(N__34990),
            .I(N__34984));
    Span4Mux_v I__6632 (
            .O(N__34987),
            .I(N__34979));
    LocalMux I__6631 (
            .O(N__34984),
            .I(N__34979));
    Odrv4 I__6630 (
            .O(N__34979),
            .I(sDAC_mem_19_1_sqmuxa));
    InMux I__6629 (
            .O(N__34976),
            .I(N__34973));
    LocalMux I__6628 (
            .O(N__34973),
            .I(N__34970));
    Span12Mux_v I__6627 (
            .O(N__34970),
            .I(N__34967));
    Odrv12 I__6626 (
            .O(N__34967),
            .I(sDAC_mem_35Z0Z_7));
    InMux I__6625 (
            .O(N__34964),
            .I(N__34961));
    LocalMux I__6624 (
            .O(N__34961),
            .I(sDAC_data_2_6_bm_1_10));
    CascadeMux I__6623 (
            .O(N__34958),
            .I(sDAC_data_RNO_15Z0Z_10_cascade_));
    InMux I__6622 (
            .O(N__34955),
            .I(N__34952));
    LocalMux I__6621 (
            .O(N__34952),
            .I(N__34949));
    Odrv4 I__6620 (
            .O(N__34949),
            .I(sDAC_data_RNO_5Z0Z_10));
    CascadeMux I__6619 (
            .O(N__34946),
            .I(sDAC_data_2_14_ns_1_10_cascade_));
    InMux I__6618 (
            .O(N__34943),
            .I(N__34940));
    LocalMux I__6617 (
            .O(N__34940),
            .I(sDAC_data_RNO_1Z0Z_10));
    InMux I__6616 (
            .O(N__34937),
            .I(N__34934));
    LocalMux I__6615 (
            .O(N__34934),
            .I(N__34931));
    Span4Mux_h I__6614 (
            .O(N__34931),
            .I(N__34928));
    Span4Mux_v I__6613 (
            .O(N__34928),
            .I(N__34925));
    Span4Mux_v I__6612 (
            .O(N__34925),
            .I(N__34922));
    Odrv4 I__6611 (
            .O(N__34922),
            .I(sDAC_mem_36Z0Z_7));
    CascadeMux I__6610 (
            .O(N__34919),
            .I(sDAC_data_2_13_am_1_10_cascade_));
    InMux I__6609 (
            .O(N__34916),
            .I(N__34913));
    LocalMux I__6608 (
            .O(N__34913),
            .I(sDAC_data_RNO_4Z0Z_10));
    InMux I__6607 (
            .O(N__34910),
            .I(N__34907));
    LocalMux I__6606 (
            .O(N__34907),
            .I(sDAC_data_RNO_26Z0Z_10));
    InMux I__6605 (
            .O(N__34904),
            .I(N__34901));
    LocalMux I__6604 (
            .O(N__34901),
            .I(sDAC_data_RNO_14Z0Z_10));
    CascadeMux I__6603 (
            .O(N__34898),
            .I(sDAC_data_2_20_am_1_3_cascade_));
    InMux I__6602 (
            .O(N__34895),
            .I(N__34892));
    LocalMux I__6601 (
            .O(N__34892),
            .I(N__34889));
    Span4Mux_h I__6600 (
            .O(N__34889),
            .I(N__34886));
    Odrv4 I__6599 (
            .O(N__34886),
            .I(sDAC_data_2_24_ns_1_3));
    CascadeMux I__6598 (
            .O(N__34883),
            .I(sDAC_data_RNO_7Z0Z_3_cascade_));
    InMux I__6597 (
            .O(N__34880),
            .I(N__34877));
    LocalMux I__6596 (
            .O(N__34877),
            .I(sDAC_data_RNO_8Z0Z_3));
    InMux I__6595 (
            .O(N__34874),
            .I(N__34871));
    LocalMux I__6594 (
            .O(N__34871),
            .I(N__34868));
    Span4Mux_v I__6593 (
            .O(N__34868),
            .I(N__34863));
    InMux I__6592 (
            .O(N__34867),
            .I(N__34860));
    CascadeMux I__6591 (
            .O(N__34866),
            .I(N__34854));
    Span4Mux_h I__6590 (
            .O(N__34863),
            .I(N__34850));
    LocalMux I__6589 (
            .O(N__34860),
            .I(N__34847));
    InMux I__6588 (
            .O(N__34859),
            .I(N__34836));
    InMux I__6587 (
            .O(N__34858),
            .I(N__34836));
    InMux I__6586 (
            .O(N__34857),
            .I(N__34836));
    InMux I__6585 (
            .O(N__34854),
            .I(N__34836));
    InMux I__6584 (
            .O(N__34853),
            .I(N__34836));
    Odrv4 I__6583 (
            .O(N__34850),
            .I(N_333));
    Odrv12 I__6582 (
            .O(N__34847),
            .I(N_333));
    LocalMux I__6581 (
            .O(N__34836),
            .I(N_333));
    InMux I__6580 (
            .O(N__34829),
            .I(N__34826));
    LocalMux I__6579 (
            .O(N__34826),
            .I(sDAC_mem_19Z0Z_0));
    InMux I__6578 (
            .O(N__34823),
            .I(N__34820));
    LocalMux I__6577 (
            .O(N__34820),
            .I(N__34817));
    Span4Mux_h I__6576 (
            .O(N__34817),
            .I(N__34814));
    Span4Mux_h I__6575 (
            .O(N__34814),
            .I(N__34811));
    Odrv4 I__6574 (
            .O(N__34811),
            .I(sDAC_mem_18Z0Z_0));
    InMux I__6573 (
            .O(N__34808),
            .I(N__34805));
    LocalMux I__6572 (
            .O(N__34805),
            .I(sDAC_mem_19Z0Z_1));
    InMux I__6571 (
            .O(N__34802),
            .I(N__34799));
    LocalMux I__6570 (
            .O(N__34799),
            .I(N__34796));
    Span4Mux_h I__6569 (
            .O(N__34796),
            .I(N__34793));
    Span4Mux_h I__6568 (
            .O(N__34793),
            .I(N__34790));
    Odrv4 I__6567 (
            .O(N__34790),
            .I(sDAC_mem_18Z0Z_1));
    InMux I__6566 (
            .O(N__34787),
            .I(N__34784));
    LocalMux I__6565 (
            .O(N__34784),
            .I(N__34781));
    Span4Mux_v I__6564 (
            .O(N__34781),
            .I(N__34778));
    Odrv4 I__6563 (
            .O(N__34778),
            .I(sDAC_data_RNO_29Z0Z_4));
    InMux I__6562 (
            .O(N__34775),
            .I(N__34772));
    LocalMux I__6561 (
            .O(N__34772),
            .I(sDAC_mem_19Z0Z_2));
    InMux I__6560 (
            .O(N__34769),
            .I(N__34766));
    LocalMux I__6559 (
            .O(N__34766),
            .I(N__34763));
    Span12Mux_v I__6558 (
            .O(N__34763),
            .I(N__34760));
    Odrv12 I__6557 (
            .O(N__34760),
            .I(sDAC_mem_18Z0Z_2));
    InMux I__6556 (
            .O(N__34757),
            .I(N__34754));
    LocalMux I__6555 (
            .O(N__34754),
            .I(N__34751));
    Span4Mux_v I__6554 (
            .O(N__34751),
            .I(N__34748));
    Span4Mux_v I__6553 (
            .O(N__34748),
            .I(N__34745));
    Odrv4 I__6552 (
            .O(N__34745),
            .I(sDAC_mem_40Z0Z_2));
    InMux I__6551 (
            .O(N__34742),
            .I(N__34739));
    LocalMux I__6550 (
            .O(N__34739),
            .I(N__34736));
    Span4Mux_v I__6549 (
            .O(N__34736),
            .I(N__34733));
    Span4Mux_h I__6548 (
            .O(N__34733),
            .I(N__34730));
    Odrv4 I__6547 (
            .O(N__34730),
            .I(sDAC_mem_8Z0Z_2));
    CascadeMux I__6546 (
            .O(N__34727),
            .I(sDAC_data_2_20_am_1_5_cascade_));
    InMux I__6545 (
            .O(N__34724),
            .I(N__34721));
    LocalMux I__6544 (
            .O(N__34721),
            .I(N__34718));
    Odrv4 I__6543 (
            .O(N__34718),
            .I(sDAC_data_2_24_ns_1_5));
    CascadeMux I__6542 (
            .O(N__34715),
            .I(sDAC_data_RNO_7Z0Z_5_cascade_));
    InMux I__6541 (
            .O(N__34712),
            .I(N__34709));
    LocalMux I__6540 (
            .O(N__34709),
            .I(sDAC_data_RNO_8Z0Z_5));
    InMux I__6539 (
            .O(N__34706),
            .I(N__34703));
    LocalMux I__6538 (
            .O(N__34703),
            .I(N__34700));
    Span4Mux_h I__6537 (
            .O(N__34700),
            .I(N__34697));
    Odrv4 I__6536 (
            .O(N__34697),
            .I(sDAC_mem_34Z0Z_0));
    InMux I__6535 (
            .O(N__34694),
            .I(N__34691));
    LocalMux I__6534 (
            .O(N__34691),
            .I(N__34688));
    Span4Mux_v I__6533 (
            .O(N__34688),
            .I(N__34685));
    Odrv4 I__6532 (
            .O(N__34685),
            .I(sDAC_mem_2Z0Z_0));
    InMux I__6531 (
            .O(N__34682),
            .I(N__34679));
    LocalMux I__6530 (
            .O(N__34679),
            .I(N__34676));
    Span4Mux_h I__6529 (
            .O(N__34676),
            .I(N__34673));
    Span4Mux_v I__6528 (
            .O(N__34673),
            .I(N__34670));
    Span4Mux_h I__6527 (
            .O(N__34670),
            .I(N__34667));
    Odrv4 I__6526 (
            .O(N__34667),
            .I(sDAC_mem_35Z0Z_0));
    CascadeMux I__6525 (
            .O(N__34664),
            .I(sDAC_data_2_6_bm_1_3_cascade_));
    InMux I__6524 (
            .O(N__34661),
            .I(N__34658));
    LocalMux I__6523 (
            .O(N__34658),
            .I(sDAC_mem_3Z0Z_0));
    InMux I__6522 (
            .O(N__34655),
            .I(N__34652));
    LocalMux I__6521 (
            .O(N__34652),
            .I(N__34649));
    Span4Mux_h I__6520 (
            .O(N__34649),
            .I(N__34646));
    Span4Mux_h I__6519 (
            .O(N__34646),
            .I(N__34643));
    Span4Mux_v I__6518 (
            .O(N__34643),
            .I(N__34640));
    Odrv4 I__6517 (
            .O(N__34640),
            .I(sDAC_mem_42Z0Z_0));
    InMux I__6516 (
            .O(N__34637),
            .I(N__34634));
    LocalMux I__6515 (
            .O(N__34634),
            .I(N__34631));
    Sp12to4 I__6514 (
            .O(N__34631),
            .I(N__34628));
    Span12Mux_v I__6513 (
            .O(N__34628),
            .I(N__34625));
    Odrv12 I__6512 (
            .O(N__34625),
            .I(sDAC_mem_10Z0Z_0));
    CascadeMux I__6511 (
            .O(N__34622),
            .I(sDAC_data_RNO_17Z0Z_3_cascade_));
    InMux I__6510 (
            .O(N__34619),
            .I(N__34616));
    LocalMux I__6509 (
            .O(N__34616),
            .I(N__34613));
    Span12Mux_v I__6508 (
            .O(N__34613),
            .I(N__34610));
    Odrv12 I__6507 (
            .O(N__34610),
            .I(sDAC_mem_11Z0Z_0));
    InMux I__6506 (
            .O(N__34607),
            .I(N__34604));
    LocalMux I__6505 (
            .O(N__34604),
            .I(N__34601));
    Span4Mux_v I__6504 (
            .O(N__34601),
            .I(N__34598));
    Span4Mux_v I__6503 (
            .O(N__34598),
            .I(N__34595));
    Odrv4 I__6502 (
            .O(N__34595),
            .I(sDAC_mem_40Z0Z_0));
    InMux I__6501 (
            .O(N__34592),
            .I(N__34589));
    LocalMux I__6500 (
            .O(N__34589),
            .I(N__34586));
    Span4Mux_v I__6499 (
            .O(N__34586),
            .I(N__34583));
    Span4Mux_h I__6498 (
            .O(N__34583),
            .I(N__34580));
    Odrv4 I__6497 (
            .O(N__34580),
            .I(sDAC_mem_8Z0Z_0));
    InMux I__6496 (
            .O(N__34577),
            .I(sDAC_mem_pointer_0_cry_1));
    InMux I__6495 (
            .O(N__34574),
            .I(sDAC_mem_pointer_0_cry_2));
    InMux I__6494 (
            .O(N__34571),
            .I(sDAC_mem_pointer_0_cry_3));
    InMux I__6493 (
            .O(N__34568),
            .I(sDAC_mem_pointer_0_cry_4));
    InMux I__6492 (
            .O(N__34565),
            .I(N__34562));
    LocalMux I__6491 (
            .O(N__34562),
            .I(N__34559));
    Span4Mux_h I__6490 (
            .O(N__34559),
            .I(N__34556));
    Odrv4 I__6489 (
            .O(N__34556),
            .I(sDAC_mem_34Z0Z_2));
    InMux I__6488 (
            .O(N__34553),
            .I(N__34550));
    LocalMux I__6487 (
            .O(N__34550),
            .I(N__34547));
    Span4Mux_h I__6486 (
            .O(N__34547),
            .I(N__34544));
    Odrv4 I__6485 (
            .O(N__34544),
            .I(sDAC_mem_2Z0Z_2));
    InMux I__6484 (
            .O(N__34541),
            .I(N__34538));
    LocalMux I__6483 (
            .O(N__34538),
            .I(N__34535));
    Span4Mux_h I__6482 (
            .O(N__34535),
            .I(N__34532));
    Span4Mux_h I__6481 (
            .O(N__34532),
            .I(N__34529));
    Span4Mux_h I__6480 (
            .O(N__34529),
            .I(N__34526));
    Odrv4 I__6479 (
            .O(N__34526),
            .I(sDAC_mem_35Z0Z_2));
    CascadeMux I__6478 (
            .O(N__34523),
            .I(sDAC_data_2_6_bm_1_5_cascade_));
    InMux I__6477 (
            .O(N__34520),
            .I(N__34517));
    LocalMux I__6476 (
            .O(N__34517),
            .I(sDAC_mem_3Z0Z_2));
    InMux I__6475 (
            .O(N__34514),
            .I(N__34511));
    LocalMux I__6474 (
            .O(N__34511),
            .I(N__34508));
    Span12Mux_v I__6473 (
            .O(N__34508),
            .I(N__34505));
    Odrv12 I__6472 (
            .O(N__34505),
            .I(sDAC_mem_42Z0Z_2));
    InMux I__6471 (
            .O(N__34502),
            .I(N__34499));
    LocalMux I__6470 (
            .O(N__34499),
            .I(N__34496));
    Span4Mux_v I__6469 (
            .O(N__34496),
            .I(N__34493));
    Span4Mux_h I__6468 (
            .O(N__34493),
            .I(N__34490));
    Odrv4 I__6467 (
            .O(N__34490),
            .I(sDAC_mem_10Z0Z_2));
    CascadeMux I__6466 (
            .O(N__34487),
            .I(sDAC_data_RNO_17Z0Z_5_cascade_));
    InMux I__6465 (
            .O(N__34484),
            .I(N__34481));
    LocalMux I__6464 (
            .O(N__34481),
            .I(N__34478));
    Span4Mux_h I__6463 (
            .O(N__34478),
            .I(N__34475));
    Span4Mux_h I__6462 (
            .O(N__34475),
            .I(N__34472));
    Odrv4 I__6461 (
            .O(N__34472),
            .I(sDAC_mem_11Z0Z_2));
    CascadeMux I__6460 (
            .O(N__34469),
            .I(sDAC_data_RNO_26Z0Z_9_cascade_));
    InMux I__6459 (
            .O(N__34466),
            .I(N__34463));
    LocalMux I__6458 (
            .O(N__34463),
            .I(sDAC_mem_32Z0Z_6));
    InMux I__6457 (
            .O(N__34460),
            .I(N__34457));
    LocalMux I__6456 (
            .O(N__34457),
            .I(sDAC_data_RNO_14Z0Z_9));
    InMux I__6455 (
            .O(N__34454),
            .I(N__34451));
    LocalMux I__6454 (
            .O(N__34451),
            .I(N__34448));
    Odrv12 I__6453 (
            .O(N__34448),
            .I(sDAC_mem_21Z0Z_0));
    InMux I__6452 (
            .O(N__34445),
            .I(N__34442));
    LocalMux I__6451 (
            .O(N__34442),
            .I(N__34439));
    Odrv12 I__6450 (
            .O(N__34439),
            .I(sDAC_mem_21Z0Z_1));
    InMux I__6449 (
            .O(N__34436),
            .I(N__34433));
    LocalMux I__6448 (
            .O(N__34433),
            .I(N__34430));
    Span4Mux_v I__6447 (
            .O(N__34430),
            .I(N__34427));
    Odrv4 I__6446 (
            .O(N__34427),
            .I(sDAC_data_RNO_20Z0Z_4));
    InMux I__6445 (
            .O(N__34424),
            .I(N__34421));
    LocalMux I__6444 (
            .O(N__34421),
            .I(N__34418));
    Odrv4 I__6443 (
            .O(N__34418),
            .I(sDAC_mem_21Z0Z_2));
    InMux I__6442 (
            .O(N__34415),
            .I(N__34412));
    LocalMux I__6441 (
            .O(N__34412),
            .I(N__34409));
    Odrv4 I__6440 (
            .O(N__34409),
            .I(sDAC_mem_21Z0Z_3));
    InMux I__6439 (
            .O(N__34406),
            .I(N__34403));
    LocalMux I__6438 (
            .O(N__34403),
            .I(N__34400));
    Span4Mux_h I__6437 (
            .O(N__34400),
            .I(N__34397));
    Odrv4 I__6436 (
            .O(N__34397),
            .I(sDAC_data_RNO_20Z0Z_6));
    InMux I__6435 (
            .O(N__34394),
            .I(N__34391));
    LocalMux I__6434 (
            .O(N__34391),
            .I(N__34388));
    Odrv4 I__6433 (
            .O(N__34388),
            .I(sDAC_mem_21Z0Z_4));
    InMux I__6432 (
            .O(N__34385),
            .I(N__34382));
    LocalMux I__6431 (
            .O(N__34382),
            .I(N__34379));
    Odrv4 I__6430 (
            .O(N__34379),
            .I(sDAC_data_RNO_20Z0Z_7));
    InMux I__6429 (
            .O(N__34376),
            .I(N__34373));
    LocalMux I__6428 (
            .O(N__34373),
            .I(N__34370));
    Span4Mux_h I__6427 (
            .O(N__34370),
            .I(N__34367));
    Odrv4 I__6426 (
            .O(N__34367),
            .I(sDAC_mem_34Z0Z_6));
    InMux I__6425 (
            .O(N__34364),
            .I(N__34361));
    LocalMux I__6424 (
            .O(N__34361),
            .I(N__34358));
    Odrv12 I__6423 (
            .O(N__34358),
            .I(sDAC_mem_2Z0Z_6));
    InMux I__6422 (
            .O(N__34355),
            .I(N__34352));
    LocalMux I__6421 (
            .O(N__34352),
            .I(N__34349));
    Odrv12 I__6420 (
            .O(N__34349),
            .I(sDAC_mem_35Z0Z_6));
    CascadeMux I__6419 (
            .O(N__34346),
            .I(sDAC_data_2_6_bm_1_9_cascade_));
    InMux I__6418 (
            .O(N__34343),
            .I(N__34340));
    LocalMux I__6417 (
            .O(N__34340),
            .I(sDAC_mem_3Z0Z_6));
    InMux I__6416 (
            .O(N__34337),
            .I(N__34334));
    LocalMux I__6415 (
            .O(N__34334),
            .I(sDAC_data_RNO_15Z0Z_9));
    InMux I__6414 (
            .O(N__34331),
            .I(N__34328));
    LocalMux I__6413 (
            .O(N__34328),
            .I(N__34325));
    Span4Mux_h I__6412 (
            .O(N__34325),
            .I(N__34322));
    Span4Mux_h I__6411 (
            .O(N__34322),
            .I(N__34319));
    Odrv4 I__6410 (
            .O(N__34319),
            .I(sDAC_mem_42Z0Z_6));
    InMux I__6409 (
            .O(N__34316),
            .I(N__34313));
    LocalMux I__6408 (
            .O(N__34313),
            .I(N__34310));
    Span4Mux_h I__6407 (
            .O(N__34310),
            .I(N__34307));
    Span4Mux_h I__6406 (
            .O(N__34307),
            .I(N__34304));
    Odrv4 I__6405 (
            .O(N__34304),
            .I(sDAC_mem_10Z0Z_6));
    CascadeMux I__6404 (
            .O(N__34301),
            .I(sDAC_data_RNO_17Z0Z_9_cascade_));
    InMux I__6403 (
            .O(N__34298),
            .I(N__34295));
    LocalMux I__6402 (
            .O(N__34295),
            .I(N__34292));
    Odrv12 I__6401 (
            .O(N__34292),
            .I(sDAC_mem_11Z0Z_6));
    InMux I__6400 (
            .O(N__34289),
            .I(N__34286));
    LocalMux I__6399 (
            .O(N__34286),
            .I(N__34283));
    Span4Mux_h I__6398 (
            .O(N__34283),
            .I(N__34280));
    Odrv4 I__6397 (
            .O(N__34280),
            .I(sDAC_mem_40Z0Z_6));
    InMux I__6396 (
            .O(N__34277),
            .I(N__34274));
    LocalMux I__6395 (
            .O(N__34274),
            .I(N__34271));
    Span4Mux_h I__6394 (
            .O(N__34271),
            .I(N__34268));
    Odrv4 I__6393 (
            .O(N__34268),
            .I(sDAC_mem_8Z0Z_6));
    CascadeMux I__6392 (
            .O(N__34265),
            .I(sDAC_data_2_20_am_1_9_cascade_));
    CascadeMux I__6391 (
            .O(N__34262),
            .I(sDAC_data_RNO_7Z0Z_9_cascade_));
    InMux I__6390 (
            .O(N__34259),
            .I(N__34256));
    LocalMux I__6389 (
            .O(N__34256),
            .I(sDAC_data_RNO_8Z0Z_9));
    InMux I__6388 (
            .O(N__34253),
            .I(N__34250));
    LocalMux I__6387 (
            .O(N__34250),
            .I(sDAC_data_RNO_2Z0Z_9));
    CEMux I__6386 (
            .O(N__34247),
            .I(N__34244));
    LocalMux I__6385 (
            .O(N__34244),
            .I(N__34241));
    Span4Mux_h I__6384 (
            .O(N__34241),
            .I(N__34238));
    Odrv4 I__6383 (
            .O(N__34238),
            .I(sDAC_mem_21_1_sqmuxa));
    InMux I__6382 (
            .O(N__34235),
            .I(N__34232));
    LocalMux I__6381 (
            .O(N__34232),
            .I(N__34229));
    Span4Mux_v I__6380 (
            .O(N__34229),
            .I(N__34226));
    Odrv4 I__6379 (
            .O(N__34226),
            .I(sDAC_mem_34Z0Z_4));
    InMux I__6378 (
            .O(N__34223),
            .I(N__34220));
    LocalMux I__6377 (
            .O(N__34220),
            .I(N__34217));
    Span4Mux_h I__6376 (
            .O(N__34217),
            .I(N__34214));
    Odrv4 I__6375 (
            .O(N__34214),
            .I(sDAC_mem_2Z0Z_4));
    InMux I__6374 (
            .O(N__34211),
            .I(N__34208));
    LocalMux I__6373 (
            .O(N__34208),
            .I(N__34205));
    Span4Mux_v I__6372 (
            .O(N__34205),
            .I(N__34202));
    Sp12to4 I__6371 (
            .O(N__34202),
            .I(N__34199));
    Odrv12 I__6370 (
            .O(N__34199),
            .I(sDAC_mem_35Z0Z_4));
    CascadeMux I__6369 (
            .O(N__34196),
            .I(sDAC_data_2_6_bm_1_7_cascade_));
    InMux I__6368 (
            .O(N__34193),
            .I(N__34190));
    LocalMux I__6367 (
            .O(N__34190),
            .I(sDAC_mem_3Z0Z_4));
    InMux I__6366 (
            .O(N__34187),
            .I(N__34184));
    LocalMux I__6365 (
            .O(N__34184),
            .I(sDAC_data_RNO_15Z0Z_7));
    InMux I__6364 (
            .O(N__34181),
            .I(N__34178));
    LocalMux I__6363 (
            .O(N__34178),
            .I(N__34175));
    Span4Mux_h I__6362 (
            .O(N__34175),
            .I(N__34172));
    Odrv4 I__6361 (
            .O(N__34172),
            .I(sDAC_mem_40Z0Z_4));
    InMux I__6360 (
            .O(N__34169),
            .I(N__34166));
    LocalMux I__6359 (
            .O(N__34166),
            .I(N__34163));
    Span12Mux_v I__6358 (
            .O(N__34163),
            .I(N__34160));
    Odrv12 I__6357 (
            .O(N__34160),
            .I(sDAC_mem_8Z0Z_4));
    CascadeMux I__6356 (
            .O(N__34157),
            .I(sDAC_data_2_20_am_1_7_cascade_));
    InMux I__6355 (
            .O(N__34154),
            .I(N__34151));
    LocalMux I__6354 (
            .O(N__34151),
            .I(N__34148));
    Odrv4 I__6353 (
            .O(N__34148),
            .I(sDAC_data_2_24_ns_1_7));
    CascadeMux I__6352 (
            .O(N__34145),
            .I(sDAC_data_RNO_7Z0Z_7_cascade_));
    InMux I__6351 (
            .O(N__34142),
            .I(N__34139));
    LocalMux I__6350 (
            .O(N__34139),
            .I(sDAC_data_RNO_2Z0Z_7));
    InMux I__6349 (
            .O(N__34136),
            .I(N__34133));
    LocalMux I__6348 (
            .O(N__34133),
            .I(N__34130));
    Span4Mux_h I__6347 (
            .O(N__34130),
            .I(N__34127));
    Span4Mux_h I__6346 (
            .O(N__34127),
            .I(N__34124));
    Odrv4 I__6345 (
            .O(N__34124),
            .I(sDAC_mem_11Z0Z_4));
    InMux I__6344 (
            .O(N__34121),
            .I(N__34118));
    LocalMux I__6343 (
            .O(N__34118),
            .I(sDAC_data_RNO_8Z0Z_7));
    InMux I__6342 (
            .O(N__34115),
            .I(N__34112));
    LocalMux I__6341 (
            .O(N__34112),
            .I(N__34109));
    Odrv12 I__6340 (
            .O(N__34109),
            .I(sDAC_mem_42Z0Z_4));
    InMux I__6339 (
            .O(N__34106),
            .I(N__34103));
    LocalMux I__6338 (
            .O(N__34103),
            .I(N__34100));
    Odrv12 I__6337 (
            .O(N__34100),
            .I(sDAC_mem_10Z0Z_4));
    InMux I__6336 (
            .O(N__34097),
            .I(N__34094));
    LocalMux I__6335 (
            .O(N__34094),
            .I(sDAC_data_RNO_17Z0Z_7));
    InMux I__6334 (
            .O(N__34091),
            .I(N__34088));
    LocalMux I__6333 (
            .O(N__34088),
            .I(N__34085));
    Span4Mux_h I__6332 (
            .O(N__34085),
            .I(N__34082));
    Odrv4 I__6331 (
            .O(N__34082),
            .I(sDAC_mem_19Z0Z_6));
    InMux I__6330 (
            .O(N__34079),
            .I(N__34076));
    LocalMux I__6329 (
            .O(N__34076),
            .I(N__34073));
    Sp12to4 I__6328 (
            .O(N__34073),
            .I(N__34070));
    Odrv12 I__6327 (
            .O(N__34070),
            .I(sDAC_mem_19Z0Z_7));
    InMux I__6326 (
            .O(N__34067),
            .I(N__34064));
    LocalMux I__6325 (
            .O(N__34064),
            .I(N__34061));
    Odrv4 I__6324 (
            .O(N__34061),
            .I(sDAC_mem_21Z0Z_5));
    InMux I__6323 (
            .O(N__34058),
            .I(N__34055));
    LocalMux I__6322 (
            .O(N__34055),
            .I(N__34052));
    Span4Mux_h I__6321 (
            .O(N__34052),
            .I(N__34049));
    Odrv4 I__6320 (
            .O(N__34049),
            .I(sDAC_mem_21Z0Z_6));
    InMux I__6319 (
            .O(N__34046),
            .I(N__34043));
    LocalMux I__6318 (
            .O(N__34043),
            .I(N__34040));
    Span4Mux_v I__6317 (
            .O(N__34040),
            .I(N__34037));
    Span4Mux_v I__6316 (
            .O(N__34037),
            .I(N__34034));
    Odrv4 I__6315 (
            .O(N__34034),
            .I(sDAC_mem_21Z0Z_7));
    CascadeMux I__6314 (
            .O(N__34031),
            .I(sRead_data_RNOZ0Z_0_cascade_));
    IoInMux I__6313 (
            .O(N__34028),
            .I(N__34025));
    LocalMux I__6312 (
            .O(N__34025),
            .I(N__34022));
    IoSpan4Mux I__6311 (
            .O(N__34022),
            .I(N__34019));
    IoSpan4Mux I__6310 (
            .O(N__34019),
            .I(N__34016));
    Span4Mux_s3_v I__6309 (
            .O(N__34016),
            .I(N__34010));
    InMux I__6308 (
            .O(N__34015),
            .I(N__34007));
    InMux I__6307 (
            .O(N__34014),
            .I(N__34001));
    InMux I__6306 (
            .O(N__34013),
            .I(N__34001));
    Span4Mux_v I__6305 (
            .O(N__34010),
            .I(N__33996));
    LocalMux I__6304 (
            .O(N__34007),
            .I(N__33996));
    InMux I__6303 (
            .O(N__34006),
            .I(N__33993));
    LocalMux I__6302 (
            .O(N__34001),
            .I(N__33990));
    Odrv4 I__6301 (
            .O(N__33996),
            .I(ADC_clk_c));
    LocalMux I__6300 (
            .O(N__33993),
            .I(ADC_clk_c));
    Odrv4 I__6299 (
            .O(N__33990),
            .I(ADC_clk_c));
    InMux I__6298 (
            .O(N__33983),
            .I(N__33979));
    InMux I__6297 (
            .O(N__33982),
            .I(N__33976));
    LocalMux I__6296 (
            .O(N__33979),
            .I(sRead_dataZ0));
    LocalMux I__6295 (
            .O(N__33976),
            .I(sRead_dataZ0));
    InMux I__6294 (
            .O(N__33971),
            .I(N__33968));
    LocalMux I__6293 (
            .O(N__33968),
            .I(spi_data_miso_0_sqmuxa_2_i_o2_4));
    InMux I__6292 (
            .O(N__33965),
            .I(N__33962));
    LocalMux I__6291 (
            .O(N__33962),
            .I(spi_data_miso_0_sqmuxa_2_i_o2_5));
    InMux I__6290 (
            .O(N__33959),
            .I(N__33956));
    LocalMux I__6289 (
            .O(N__33956),
            .I(N__33953));
    Span12Mux_v I__6288 (
            .O(N__33953),
            .I(N__33950));
    Span12Mux_h I__6287 (
            .O(N__33950),
            .I(N__33947));
    Odrv12 I__6286 (
            .O(N__33947),
            .I(ADC3_c));
    IoInMux I__6285 (
            .O(N__33944),
            .I(N__33941));
    LocalMux I__6284 (
            .O(N__33941),
            .I(N__33938));
    Span4Mux_s2_v I__6283 (
            .O(N__33938),
            .I(N__33935));
    Span4Mux_h I__6282 (
            .O(N__33935),
            .I(N__33932));
    Span4Mux_h I__6281 (
            .O(N__33932),
            .I(N__33929));
    Span4Mux_v I__6280 (
            .O(N__33929),
            .I(N__33926));
    Odrv4 I__6279 (
            .O(N__33926),
            .I(RAM_DATA_1Z0Z_3));
    InMux I__6278 (
            .O(N__33923),
            .I(N__33920));
    LocalMux I__6277 (
            .O(N__33920),
            .I(N__33917));
    Span4Mux_h I__6276 (
            .O(N__33917),
            .I(N__33914));
    Odrv4 I__6275 (
            .O(N__33914),
            .I(sDAC_mem_19Z0Z_4));
    InMux I__6274 (
            .O(N__33911),
            .I(N__33908));
    LocalMux I__6273 (
            .O(N__33908),
            .I(N__33905));
    Span4Mux_h I__6272 (
            .O(N__33905),
            .I(N__33902));
    Odrv4 I__6271 (
            .O(N__33902),
            .I(sDAC_mem_19Z0Z_5));
    InMux I__6270 (
            .O(N__33899),
            .I(N__33896));
    LocalMux I__6269 (
            .O(N__33896),
            .I(sDAC_mem_22Z0Z_6));
    CEMux I__6268 (
            .O(N__33893),
            .I(N__33890));
    LocalMux I__6267 (
            .O(N__33890),
            .I(N__33887));
    Span4Mux_v I__6266 (
            .O(N__33887),
            .I(N__33884));
    Span4Mux_v I__6265 (
            .O(N__33884),
            .I(N__33880));
    CEMux I__6264 (
            .O(N__33883),
            .I(N__33877));
    Span4Mux_h I__6263 (
            .O(N__33880),
            .I(N__33872));
    LocalMux I__6262 (
            .O(N__33877),
            .I(N__33872));
    Odrv4 I__6261 (
            .O(N__33872),
            .I(sDAC_mem_22_1_sqmuxa));
    InMux I__6260 (
            .O(N__33869),
            .I(N__33866));
    LocalMux I__6259 (
            .O(N__33866),
            .I(N__33863));
    Odrv12 I__6258 (
            .O(N__33863),
            .I(sDAC_mem_29Z0Z_0));
    InMux I__6257 (
            .O(N__33860),
            .I(N__33857));
    LocalMux I__6256 (
            .O(N__33857),
            .I(N__33854));
    Span4Mux_v I__6255 (
            .O(N__33854),
            .I(N__33851));
    Span4Mux_h I__6254 (
            .O(N__33851),
            .I(N__33848));
    Odrv4 I__6253 (
            .O(N__33848),
            .I(sDAC_mem_28Z0Z_0));
    InMux I__6252 (
            .O(N__33845),
            .I(N__33842));
    LocalMux I__6251 (
            .O(N__33842),
            .I(sDAC_data_RNO_23Z0Z_3));
    InMux I__6250 (
            .O(N__33839),
            .I(N__33836));
    LocalMux I__6249 (
            .O(N__33836),
            .I(N__33833));
    Span4Mux_h I__6248 (
            .O(N__33833),
            .I(N__33830));
    Odrv4 I__6247 (
            .O(N__33830),
            .I(sDAC_mem_29Z0Z_3));
    InMux I__6246 (
            .O(N__33827),
            .I(N__33824));
    LocalMux I__6245 (
            .O(N__33824),
            .I(N__33821));
    Span4Mux_h I__6244 (
            .O(N__33821),
            .I(N__33818));
    Span4Mux_h I__6243 (
            .O(N__33818),
            .I(N__33815));
    Odrv4 I__6242 (
            .O(N__33815),
            .I(sDAC_mem_28Z0Z_3));
    CascadeMux I__6241 (
            .O(N__33812),
            .I(sbuttonModeStatus_0_sqmuxa_14_cascade_));
    InMux I__6240 (
            .O(N__33809),
            .I(N__33806));
    LocalMux I__6239 (
            .O(N__33806),
            .I(sbuttonModeStatus_0_sqmuxa_13));
    InMux I__6238 (
            .O(N__33803),
            .I(N__33800));
    LocalMux I__6237 (
            .O(N__33800),
            .I(N__33797));
    Span4Mux_h I__6236 (
            .O(N__33797),
            .I(N__33794));
    Odrv4 I__6235 (
            .O(N__33794),
            .I(sbuttonModeStatus_0_sqmuxa_22));
    InMux I__6234 (
            .O(N__33791),
            .I(N__33788));
    LocalMux I__6233 (
            .O(N__33788),
            .I(N__33785));
    Span4Mux_h I__6232 (
            .O(N__33785),
            .I(N__33782));
    Span4Mux_h I__6231 (
            .O(N__33782),
            .I(N__33779));
    Span4Mux_v I__6230 (
            .O(N__33779),
            .I(N__33776));
    Odrv4 I__6229 (
            .O(N__33776),
            .I(sEEPonPoff_1_sqmuxa_0_a3_0_a2_1));
    InMux I__6228 (
            .O(N__33773),
            .I(N__33770));
    LocalMux I__6227 (
            .O(N__33770),
            .I(N__33765));
    InMux I__6226 (
            .O(N__33769),
            .I(N__33762));
    InMux I__6225 (
            .O(N__33768),
            .I(N__33759));
    Span4Mux_v I__6224 (
            .O(N__33765),
            .I(N__33756));
    LocalMux I__6223 (
            .O(N__33762),
            .I(N__33751));
    LocalMux I__6222 (
            .O(N__33759),
            .I(N__33748));
    Span4Mux_h I__6221 (
            .O(N__33756),
            .I(N__33740));
    InMux I__6220 (
            .O(N__33755),
            .I(N__33734));
    InMux I__6219 (
            .O(N__33754),
            .I(N__33734));
    Span12Mux_v I__6218 (
            .O(N__33751),
            .I(N__33729));
    Span4Mux_v I__6217 (
            .O(N__33748),
            .I(N__33726));
    InMux I__6216 (
            .O(N__33747),
            .I(N__33723));
    InMux I__6215 (
            .O(N__33746),
            .I(N__33718));
    InMux I__6214 (
            .O(N__33745),
            .I(N__33718));
    InMux I__6213 (
            .O(N__33744),
            .I(N__33715));
    InMux I__6212 (
            .O(N__33743),
            .I(N__33712));
    Span4Mux_h I__6211 (
            .O(N__33740),
            .I(N__33709));
    InMux I__6210 (
            .O(N__33739),
            .I(N__33706));
    LocalMux I__6209 (
            .O(N__33734),
            .I(N__33703));
    InMux I__6208 (
            .O(N__33733),
            .I(N__33698));
    InMux I__6207 (
            .O(N__33732),
            .I(N__33698));
    Odrv12 I__6206 (
            .O(N__33729),
            .I(sPointer_RNI5LBD1Z0Z_0));
    Odrv4 I__6205 (
            .O(N__33726),
            .I(sPointer_RNI5LBD1Z0Z_0));
    LocalMux I__6204 (
            .O(N__33723),
            .I(sPointer_RNI5LBD1Z0Z_0));
    LocalMux I__6203 (
            .O(N__33718),
            .I(sPointer_RNI5LBD1Z0Z_0));
    LocalMux I__6202 (
            .O(N__33715),
            .I(sPointer_RNI5LBD1Z0Z_0));
    LocalMux I__6201 (
            .O(N__33712),
            .I(sPointer_RNI5LBD1Z0Z_0));
    Odrv4 I__6200 (
            .O(N__33709),
            .I(sPointer_RNI5LBD1Z0Z_0));
    LocalMux I__6199 (
            .O(N__33706),
            .I(sPointer_RNI5LBD1Z0Z_0));
    Odrv4 I__6198 (
            .O(N__33703),
            .I(sPointer_RNI5LBD1Z0Z_0));
    LocalMux I__6197 (
            .O(N__33698),
            .I(sPointer_RNI5LBD1Z0Z_0));
    CEMux I__6196 (
            .O(N__33677),
            .I(N__33674));
    LocalMux I__6195 (
            .O(N__33674),
            .I(sEEPonPoff_1_sqmuxa));
    IoInMux I__6194 (
            .O(N__33671),
            .I(N__33668));
    LocalMux I__6193 (
            .O(N__33668),
            .I(N__33665));
    IoSpan4Mux I__6192 (
            .O(N__33665),
            .I(N__33662));
    IoSpan4Mux I__6191 (
            .O(N__33662),
            .I(N__33659));
    Span4Mux_s2_h I__6190 (
            .O(N__33659),
            .I(N__33656));
    Sp12to4 I__6189 (
            .O(N__33656),
            .I(N__33653));
    Odrv12 I__6188 (
            .O(N__33653),
            .I(RAM_nWE_0_i));
    InMux I__6187 (
            .O(N__33650),
            .I(N__33647));
    LocalMux I__6186 (
            .O(N__33647),
            .I(sDAC_mem_27Z0Z_0));
    InMux I__6185 (
            .O(N__33644),
            .I(N__33641));
    LocalMux I__6184 (
            .O(N__33641),
            .I(N__33638));
    Odrv12 I__6183 (
            .O(N__33638),
            .I(sDAC_mem_26Z0Z_0));
    InMux I__6182 (
            .O(N__33635),
            .I(N__33632));
    LocalMux I__6181 (
            .O(N__33632),
            .I(N__33629));
    Span4Mux_v I__6180 (
            .O(N__33629),
            .I(N__33626));
    Span4Mux_h I__6179 (
            .O(N__33626),
            .I(N__33623));
    Odrv4 I__6178 (
            .O(N__33623),
            .I(sDAC_mem_24Z0Z_0));
    CascadeMux I__6177 (
            .O(N__33620),
            .I(sDAC_data_RNO_30Z0Z_3_cascade_));
    InMux I__6176 (
            .O(N__33617),
            .I(N__33614));
    LocalMux I__6175 (
            .O(N__33614),
            .I(sDAC_data_RNO_31Z0Z_3));
    InMux I__6174 (
            .O(N__33611),
            .I(N__33608));
    LocalMux I__6173 (
            .O(N__33608),
            .I(sDAC_data_RNO_24Z0Z_3));
    CascadeMux I__6172 (
            .O(N__33605),
            .I(sDAC_data_2_39_ns_1_3_cascade_));
    InMux I__6171 (
            .O(N__33602),
            .I(N__33599));
    LocalMux I__6170 (
            .O(N__33599),
            .I(N__33596));
    Span4Mux_v I__6169 (
            .O(N__33596),
            .I(N__33593));
    Span4Mux_v I__6168 (
            .O(N__33593),
            .I(N__33590));
    Odrv4 I__6167 (
            .O(N__33590),
            .I(sDAC_data_RNO_21Z0Z_7));
    InMux I__6166 (
            .O(N__33587),
            .I(N__33584));
    LocalMux I__6165 (
            .O(N__33584),
            .I(sDAC_mem_22Z0Z_4));
    InMux I__6164 (
            .O(N__33581),
            .I(N__33578));
    LocalMux I__6163 (
            .O(N__33578),
            .I(N__33575));
    Span4Mux_h I__6162 (
            .O(N__33575),
            .I(N__33572));
    Span4Mux_v I__6161 (
            .O(N__33572),
            .I(N__33569));
    Odrv4 I__6160 (
            .O(N__33569),
            .I(sDAC_data_RNO_21Z0Z_8));
    InMux I__6159 (
            .O(N__33566),
            .I(N__33563));
    LocalMux I__6158 (
            .O(N__33563),
            .I(sDAC_mem_22Z0Z_5));
    InMux I__6157 (
            .O(N__33560),
            .I(N__33557));
    LocalMux I__6156 (
            .O(N__33557),
            .I(N__33554));
    Span12Mux_v I__6155 (
            .O(N__33554),
            .I(N__33551));
    Odrv12 I__6154 (
            .O(N__33551),
            .I(sDAC_data_RNO_21Z0Z_9));
    InMux I__6153 (
            .O(N__33548),
            .I(N__33545));
    LocalMux I__6152 (
            .O(N__33545),
            .I(sDAC_data_RNO_20Z0Z_10));
    CascadeMux I__6151 (
            .O(N__33542),
            .I(N__33539));
    InMux I__6150 (
            .O(N__33539),
            .I(N__33536));
    LocalMux I__6149 (
            .O(N__33536),
            .I(N__33533));
    Span4Mux_v I__6148 (
            .O(N__33533),
            .I(N__33530));
    Span4Mux_h I__6147 (
            .O(N__33530),
            .I(N__33527));
    Odrv4 I__6146 (
            .O(N__33527),
            .I(sDAC_mem_18Z0Z_7));
    InMux I__6145 (
            .O(N__33524),
            .I(N__33521));
    LocalMux I__6144 (
            .O(N__33521),
            .I(sDAC_data_RNO_29Z0Z_10));
    InMux I__6143 (
            .O(N__33518),
            .I(N__33515));
    LocalMux I__6142 (
            .O(N__33515),
            .I(sDAC_mem_16Z0Z_7));
    CEMux I__6141 (
            .O(N__33512),
            .I(N__33509));
    LocalMux I__6140 (
            .O(N__33509),
            .I(N__33505));
    CEMux I__6139 (
            .O(N__33508),
            .I(N__33501));
    Span4Mux_h I__6138 (
            .O(N__33505),
            .I(N__33498));
    CEMux I__6137 (
            .O(N__33504),
            .I(N__33495));
    LocalMux I__6136 (
            .O(N__33501),
            .I(N__33492));
    Span4Mux_h I__6135 (
            .O(N__33498),
            .I(N__33487));
    LocalMux I__6134 (
            .O(N__33495),
            .I(N__33487));
    Span4Mux_v I__6133 (
            .O(N__33492),
            .I(N__33484));
    Span4Mux_v I__6132 (
            .O(N__33487),
            .I(N__33481));
    Span4Mux_h I__6131 (
            .O(N__33484),
            .I(N__33478));
    Span4Mux_h I__6130 (
            .O(N__33481),
            .I(N__33475));
    Odrv4 I__6129 (
            .O(N__33478),
            .I(sDAC_mem_16_1_sqmuxa));
    Odrv4 I__6128 (
            .O(N__33475),
            .I(sDAC_mem_16_1_sqmuxa));
    InMux I__6127 (
            .O(N__33470),
            .I(N__33467));
    LocalMux I__6126 (
            .O(N__33467),
            .I(sDAC_data_RNO_31Z0Z_10));
    InMux I__6125 (
            .O(N__33464),
            .I(N__33461));
    LocalMux I__6124 (
            .O(N__33461),
            .I(sDAC_data_RNO_30Z0Z_10));
    InMux I__6123 (
            .O(N__33458),
            .I(N__33455));
    LocalMux I__6122 (
            .O(N__33455),
            .I(N__33452));
    Odrv12 I__6121 (
            .O(N__33452),
            .I(sDAC_mem_31Z0Z_7));
    InMux I__6120 (
            .O(N__33449),
            .I(N__33446));
    LocalMux I__6119 (
            .O(N__33446),
            .I(N__33443));
    Span4Mux_h I__6118 (
            .O(N__33443),
            .I(N__33440));
    Span4Mux_h I__6117 (
            .O(N__33440),
            .I(N__33437));
    Odrv4 I__6116 (
            .O(N__33437),
            .I(sDAC_mem_30Z0Z_7));
    InMux I__6115 (
            .O(N__33434),
            .I(N__33431));
    LocalMux I__6114 (
            .O(N__33431),
            .I(N__33428));
    Span4Mux_h I__6113 (
            .O(N__33428),
            .I(N__33425));
    Span4Mux_h I__6112 (
            .O(N__33425),
            .I(N__33422));
    Odrv4 I__6111 (
            .O(N__33422),
            .I(sDAC_mem_29Z0Z_7));
    InMux I__6110 (
            .O(N__33419),
            .I(N__33416));
    LocalMux I__6109 (
            .O(N__33416),
            .I(sDAC_data_RNO_24Z0Z_10));
    CascadeMux I__6108 (
            .O(N__33413),
            .I(sDAC_data_RNO_23Z0Z_10_cascade_));
    InMux I__6107 (
            .O(N__33410),
            .I(N__33407));
    LocalMux I__6106 (
            .O(N__33407),
            .I(sDAC_data_2_39_ns_1_10));
    InMux I__6105 (
            .O(N__33404),
            .I(N__33401));
    LocalMux I__6104 (
            .O(N__33401),
            .I(N__33398));
    Odrv4 I__6103 (
            .O(N__33398),
            .I(sDAC_data_RNO_11Z0Z_10));
    InMux I__6102 (
            .O(N__33395),
            .I(N__33392));
    LocalMux I__6101 (
            .O(N__33392),
            .I(sDAC_mem_28Z0Z_7));
    CascadeMux I__6100 (
            .O(N__33389),
            .I(N__33385));
    CascadeMux I__6099 (
            .O(N__33388),
            .I(N__33382));
    InMux I__6098 (
            .O(N__33385),
            .I(N__33377));
    InMux I__6097 (
            .O(N__33382),
            .I(N__33370));
    CascadeMux I__6096 (
            .O(N__33381),
            .I(N__33367));
    CascadeMux I__6095 (
            .O(N__33380),
            .I(N__33363));
    LocalMux I__6094 (
            .O(N__33377),
            .I(N__33359));
    InMux I__6093 (
            .O(N__33376),
            .I(N__33356));
    InMux I__6092 (
            .O(N__33375),
            .I(N__33353));
    InMux I__6091 (
            .O(N__33374),
            .I(N__33350));
    InMux I__6090 (
            .O(N__33373),
            .I(N__33347));
    LocalMux I__6089 (
            .O(N__33370),
            .I(N__33344));
    InMux I__6088 (
            .O(N__33367),
            .I(N__33339));
    InMux I__6087 (
            .O(N__33366),
            .I(N__33339));
    InMux I__6086 (
            .O(N__33363),
            .I(N__33336));
    InMux I__6085 (
            .O(N__33362),
            .I(N__33333));
    Span4Mux_v I__6084 (
            .O(N__33359),
            .I(N__33326));
    LocalMux I__6083 (
            .O(N__33356),
            .I(N__33326));
    LocalMux I__6082 (
            .O(N__33353),
            .I(N__33321));
    LocalMux I__6081 (
            .O(N__33350),
            .I(N__33321));
    LocalMux I__6080 (
            .O(N__33347),
            .I(N__33318));
    Span4Mux_h I__6079 (
            .O(N__33344),
            .I(N__33313));
    LocalMux I__6078 (
            .O(N__33339),
            .I(N__33313));
    LocalMux I__6077 (
            .O(N__33336),
            .I(N__33310));
    LocalMux I__6076 (
            .O(N__33333),
            .I(N__33307));
    InMux I__6075 (
            .O(N__33332),
            .I(N__33304));
    InMux I__6074 (
            .O(N__33331),
            .I(N__33301));
    Span4Mux_v I__6073 (
            .O(N__33326),
            .I(N__33294));
    Span4Mux_h I__6072 (
            .O(N__33321),
            .I(N__33294));
    Span4Mux_v I__6071 (
            .O(N__33318),
            .I(N__33294));
    Span4Mux_v I__6070 (
            .O(N__33313),
            .I(N__33287));
    Span4Mux_v I__6069 (
            .O(N__33310),
            .I(N__33287));
    Span4Mux_h I__6068 (
            .O(N__33307),
            .I(N__33287));
    LocalMux I__6067 (
            .O(N__33304),
            .I(un7_spon_20));
    LocalMux I__6066 (
            .O(N__33301),
            .I(un7_spon_20));
    Odrv4 I__6065 (
            .O(N__33294),
            .I(un7_spon_20));
    Odrv4 I__6064 (
            .O(N__33287),
            .I(un7_spon_20));
    CascadeMux I__6063 (
            .O(N__33278),
            .I(N__33270));
    InMux I__6062 (
            .O(N__33277),
            .I(N__33267));
    CascadeMux I__6061 (
            .O(N__33276),
            .I(N__33264));
    CascadeMux I__6060 (
            .O(N__33275),
            .I(N__33261));
    CascadeMux I__6059 (
            .O(N__33274),
            .I(N__33258));
    InMux I__6058 (
            .O(N__33273),
            .I(N__33254));
    InMux I__6057 (
            .O(N__33270),
            .I(N__33250));
    LocalMux I__6056 (
            .O(N__33267),
            .I(N__33246));
    InMux I__6055 (
            .O(N__33264),
            .I(N__33241));
    InMux I__6054 (
            .O(N__33261),
            .I(N__33241));
    InMux I__6053 (
            .O(N__33258),
            .I(N__33238));
    InMux I__6052 (
            .O(N__33257),
            .I(N__33235));
    LocalMux I__6051 (
            .O(N__33254),
            .I(N__33232));
    InMux I__6050 (
            .O(N__33253),
            .I(N__33229));
    LocalMux I__6049 (
            .O(N__33250),
            .I(N__33226));
    InMux I__6048 (
            .O(N__33249),
            .I(N__33220));
    Span4Mux_v I__6047 (
            .O(N__33246),
            .I(N__33215));
    LocalMux I__6046 (
            .O(N__33241),
            .I(N__33215));
    LocalMux I__6045 (
            .O(N__33238),
            .I(N__33210));
    LocalMux I__6044 (
            .O(N__33235),
            .I(N__33210));
    Span4Mux_v I__6043 (
            .O(N__33232),
            .I(N__33205));
    LocalMux I__6042 (
            .O(N__33229),
            .I(N__33205));
    Span4Mux_h I__6041 (
            .O(N__33226),
            .I(N__33202));
    InMux I__6040 (
            .O(N__33225),
            .I(N__33199));
    InMux I__6039 (
            .O(N__33224),
            .I(N__33196));
    InMux I__6038 (
            .O(N__33223),
            .I(N__33193));
    LocalMux I__6037 (
            .O(N__33220),
            .I(N__33190));
    Span4Mux_v I__6036 (
            .O(N__33215),
            .I(N__33181));
    Span4Mux_h I__6035 (
            .O(N__33210),
            .I(N__33181));
    Span4Mux_v I__6034 (
            .O(N__33205),
            .I(N__33181));
    Span4Mux_v I__6033 (
            .O(N__33202),
            .I(N__33181));
    LocalMux I__6032 (
            .O(N__33199),
            .I(un7_spon_19));
    LocalMux I__6031 (
            .O(N__33196),
            .I(un7_spon_19));
    LocalMux I__6030 (
            .O(N__33193),
            .I(un7_spon_19));
    Odrv12 I__6029 (
            .O(N__33190),
            .I(un7_spon_19));
    Odrv4 I__6028 (
            .O(N__33181),
            .I(un7_spon_19));
    InMux I__6027 (
            .O(N__33170),
            .I(N__33162));
    CascadeMux I__6026 (
            .O(N__33169),
            .I(N__33158));
    CascadeMux I__6025 (
            .O(N__33168),
            .I(N__33155));
    InMux I__6024 (
            .O(N__33167),
            .I(N__33151));
    CascadeMux I__6023 (
            .O(N__33166),
            .I(N__33147));
    CascadeMux I__6022 (
            .O(N__33165),
            .I(N__33144));
    LocalMux I__6021 (
            .O(N__33162),
            .I(N__33141));
    InMux I__6020 (
            .O(N__33161),
            .I(N__33138));
    InMux I__6019 (
            .O(N__33158),
            .I(N__33135));
    InMux I__6018 (
            .O(N__33155),
            .I(N__33132));
    InMux I__6017 (
            .O(N__33154),
            .I(N__33129));
    LocalMux I__6016 (
            .O(N__33151),
            .I(N__33126));
    InMux I__6015 (
            .O(N__33150),
            .I(N__33123));
    InMux I__6014 (
            .O(N__33147),
            .I(N__33120));
    InMux I__6013 (
            .O(N__33144),
            .I(N__33117));
    Span4Mux_v I__6012 (
            .O(N__33141),
            .I(N__33110));
    LocalMux I__6011 (
            .O(N__33138),
            .I(N__33110));
    LocalMux I__6010 (
            .O(N__33135),
            .I(N__33105));
    LocalMux I__6009 (
            .O(N__33132),
            .I(N__33105));
    LocalMux I__6008 (
            .O(N__33129),
            .I(N__33102));
    Span4Mux_h I__6007 (
            .O(N__33126),
            .I(N__33097));
    LocalMux I__6006 (
            .O(N__33123),
            .I(N__33097));
    LocalMux I__6005 (
            .O(N__33120),
            .I(N__33094));
    LocalMux I__6004 (
            .O(N__33117),
            .I(N__33091));
    InMux I__6003 (
            .O(N__33116),
            .I(N__33088));
    InMux I__6002 (
            .O(N__33115),
            .I(N__33085));
    Span4Mux_v I__6001 (
            .O(N__33110),
            .I(N__33078));
    Span4Mux_h I__6000 (
            .O(N__33105),
            .I(N__33078));
    Span4Mux_v I__5999 (
            .O(N__33102),
            .I(N__33078));
    Span4Mux_v I__5998 (
            .O(N__33097),
            .I(N__33071));
    Span4Mux_v I__5997 (
            .O(N__33094),
            .I(N__33071));
    Span4Mux_h I__5996 (
            .O(N__33091),
            .I(N__33071));
    LocalMux I__5995 (
            .O(N__33088),
            .I(un7_spon_21));
    LocalMux I__5994 (
            .O(N__33085),
            .I(un7_spon_21));
    Odrv4 I__5993 (
            .O(N__33078),
            .I(un7_spon_21));
    Odrv4 I__5992 (
            .O(N__33071),
            .I(un7_spon_21));
    CascadeMux I__5991 (
            .O(N__33062),
            .I(N__33059));
    InMux I__5990 (
            .O(N__33059),
            .I(N__33054));
    InMux I__5989 (
            .O(N__33058),
            .I(N__33049));
    CascadeMux I__5988 (
            .O(N__33057),
            .I(N__33043));
    LocalMux I__5987 (
            .O(N__33054),
            .I(N__33040));
    InMux I__5986 (
            .O(N__33053),
            .I(N__33036));
    InMux I__5985 (
            .O(N__33052),
            .I(N__33033));
    LocalMux I__5984 (
            .O(N__33049),
            .I(N__33030));
    InMux I__5983 (
            .O(N__33048),
            .I(N__33027));
    InMux I__5982 (
            .O(N__33047),
            .I(N__33024));
    CascadeMux I__5981 (
            .O(N__33046),
            .I(N__33021));
    InMux I__5980 (
            .O(N__33043),
            .I(N__33018));
    Span4Mux_v I__5979 (
            .O(N__33040),
            .I(N__33014));
    InMux I__5978 (
            .O(N__33039),
            .I(N__33011));
    LocalMux I__5977 (
            .O(N__33036),
            .I(N__33008));
    LocalMux I__5976 (
            .O(N__33033),
            .I(N__33005));
    Span4Mux_v I__5975 (
            .O(N__33030),
            .I(N__33000));
    LocalMux I__5974 (
            .O(N__33027),
            .I(N__33000));
    LocalMux I__5973 (
            .O(N__33024),
            .I(N__32997));
    InMux I__5972 (
            .O(N__33021),
            .I(N__32994));
    LocalMux I__5971 (
            .O(N__33018),
            .I(N__32991));
    InMux I__5970 (
            .O(N__33017),
            .I(N__32987));
    Span4Mux_v I__5969 (
            .O(N__33014),
            .I(N__32976));
    LocalMux I__5968 (
            .O(N__33011),
            .I(N__32976));
    Span4Mux_h I__5967 (
            .O(N__33008),
            .I(N__32976));
    Span4Mux_h I__5966 (
            .O(N__33005),
            .I(N__32976));
    Span4Mux_v I__5965 (
            .O(N__33000),
            .I(N__32976));
    Span4Mux_h I__5964 (
            .O(N__32997),
            .I(N__32973));
    LocalMux I__5963 (
            .O(N__32994),
            .I(N__32970));
    Span4Mux_h I__5962 (
            .O(N__32991),
            .I(N__32967));
    InMux I__5961 (
            .O(N__32990),
            .I(N__32964));
    LocalMux I__5960 (
            .O(N__32987),
            .I(un7_spon_11));
    Odrv4 I__5959 (
            .O(N__32976),
            .I(un7_spon_11));
    Odrv4 I__5958 (
            .O(N__32973),
            .I(un7_spon_11));
    Odrv12 I__5957 (
            .O(N__32970),
            .I(un7_spon_11));
    Odrv4 I__5956 (
            .O(N__32967),
            .I(un7_spon_11));
    LocalMux I__5955 (
            .O(N__32964),
            .I(un7_spon_11));
    CascadeMux I__5954 (
            .O(N__32951),
            .I(N__32948));
    InMux I__5953 (
            .O(N__32948),
            .I(N__32945));
    LocalMux I__5952 (
            .O(N__32945),
            .I(N__32942));
    Span4Mux_h I__5951 (
            .O(N__32942),
            .I(N__32939));
    Odrv4 I__5950 (
            .O(N__32939),
            .I(g0_12));
    InMux I__5949 (
            .O(N__32936),
            .I(N__32933));
    LocalMux I__5948 (
            .O(N__32933),
            .I(sDAC_data_RNO_2Z0Z_10));
    CascadeMux I__5947 (
            .O(N__32930),
            .I(sDAC_data_2_41_ns_1_10_cascade_));
    InMux I__5946 (
            .O(N__32927),
            .I(N__32924));
    LocalMux I__5945 (
            .O(N__32924),
            .I(sDAC_data_2_10));
    InMux I__5944 (
            .O(N__32921),
            .I(N__32918));
    LocalMux I__5943 (
            .O(N__32918),
            .I(N__32915));
    Span4Mux_v I__5942 (
            .O(N__32915),
            .I(N__32912));
    Odrv4 I__5941 (
            .O(N__32912),
            .I(sbuttonModeStatus_0_sqmuxa_17));
    InMux I__5940 (
            .O(N__32909),
            .I(N__32906));
    LocalMux I__5939 (
            .O(N__32906),
            .I(N__32903));
    Span4Mux_v I__5938 (
            .O(N__32903),
            .I(N__32900));
    Span4Mux_h I__5937 (
            .O(N__32900),
            .I(N__32897));
    Span4Mux_h I__5936 (
            .O(N__32897),
            .I(N__32894));
    Odrv4 I__5935 (
            .O(N__32894),
            .I(sDAC_mem_22Z0Z_7));
    CascadeMux I__5934 (
            .O(N__32891),
            .I(sDAC_data_RNO_28Z0Z_10_cascade_));
    InMux I__5933 (
            .O(N__32888),
            .I(N__32885));
    LocalMux I__5932 (
            .O(N__32885),
            .I(sDAC_data_RNO_21Z0Z_10));
    CascadeMux I__5931 (
            .O(N__32882),
            .I(sDAC_data_2_32_ns_1_10_cascade_));
    InMux I__5930 (
            .O(N__32879),
            .I(N__32876));
    LocalMux I__5929 (
            .O(N__32876),
            .I(sDAC_data_RNO_10Z0Z_10));
    InMux I__5928 (
            .O(N__32873),
            .I(N__32870));
    LocalMux I__5927 (
            .O(N__32870),
            .I(N__32867));
    Span4Mux_h I__5926 (
            .O(N__32867),
            .I(N__32864));
    Odrv4 I__5925 (
            .O(N__32864),
            .I(sDAC_mem_34Z0Z_7));
    InMux I__5924 (
            .O(N__32861),
            .I(N__32858));
    LocalMux I__5923 (
            .O(N__32858),
            .I(sDAC_mem_2Z0Z_7));
    CEMux I__5922 (
            .O(N__32855),
            .I(N__32852));
    LocalMux I__5921 (
            .O(N__32852),
            .I(N__32848));
    CEMux I__5920 (
            .O(N__32851),
            .I(N__32845));
    Span4Mux_v I__5919 (
            .O(N__32848),
            .I(N__32842));
    LocalMux I__5918 (
            .O(N__32845),
            .I(N__32839));
    Span4Mux_h I__5917 (
            .O(N__32842),
            .I(N__32836));
    Span4Mux_h I__5916 (
            .O(N__32839),
            .I(N__32833));
    Odrv4 I__5915 (
            .O(N__32836),
            .I(sDAC_mem_2_1_sqmuxa));
    Odrv4 I__5914 (
            .O(N__32833),
            .I(sDAC_mem_2_1_sqmuxa));
    InMux I__5913 (
            .O(N__32828),
            .I(N__32825));
    LocalMux I__5912 (
            .O(N__32825),
            .I(N__32822));
    Sp12to4 I__5911 (
            .O(N__32822),
            .I(N__32819));
    Span12Mux_h I__5910 (
            .O(N__32819),
            .I(N__32816));
    Odrv12 I__5909 (
            .O(N__32816),
            .I(sDAC_mem_12Z0Z_7));
    CascadeMux I__5908 (
            .O(N__32813),
            .I(sDAC_data_RNO_18Z0Z_10_cascade_));
    InMux I__5907 (
            .O(N__32810),
            .I(N__32807));
    LocalMux I__5906 (
            .O(N__32807),
            .I(N__32804));
    Span4Mux_v I__5905 (
            .O(N__32804),
            .I(N__32801));
    Span4Mux_h I__5904 (
            .O(N__32801),
            .I(N__32798));
    Odrv4 I__5903 (
            .O(N__32798),
            .I(sDAC_mem_15Z0Z_7));
    InMux I__5902 (
            .O(N__32795),
            .I(N__32792));
    LocalMux I__5901 (
            .O(N__32792),
            .I(N__32789));
    Span4Mux_v I__5900 (
            .O(N__32789),
            .I(N__32786));
    Span4Mux_h I__5899 (
            .O(N__32786),
            .I(N__32783));
    Odrv4 I__5898 (
            .O(N__32783),
            .I(sDAC_mem_14Z0Z_7));
    InMux I__5897 (
            .O(N__32780),
            .I(N__32777));
    LocalMux I__5896 (
            .O(N__32777),
            .I(sDAC_data_RNO_19Z0Z_10));
    InMux I__5895 (
            .O(N__32774),
            .I(N__32771));
    LocalMux I__5894 (
            .O(N__32771),
            .I(N__32768));
    Span4Mux_v I__5893 (
            .O(N__32768),
            .I(N__32765));
    Span4Mux_h I__5892 (
            .O(N__32765),
            .I(N__32762));
    Odrv4 I__5891 (
            .O(N__32762),
            .I(sDAC_mem_42Z0Z_7));
    InMux I__5890 (
            .O(N__32759),
            .I(N__32756));
    LocalMux I__5889 (
            .O(N__32756),
            .I(N__32753));
    Span4Mux_h I__5888 (
            .O(N__32753),
            .I(N__32750));
    Span4Mux_h I__5887 (
            .O(N__32750),
            .I(N__32747));
    Span4Mux_v I__5886 (
            .O(N__32747),
            .I(N__32744));
    Odrv4 I__5885 (
            .O(N__32744),
            .I(sDAC_mem_10Z0Z_7));
    CascadeMux I__5884 (
            .O(N__32741),
            .I(sDAC_data_RNO_17Z0Z_10_cascade_));
    InMux I__5883 (
            .O(N__32738),
            .I(N__32735));
    LocalMux I__5882 (
            .O(N__32735),
            .I(N__32732));
    Span4Mux_v I__5881 (
            .O(N__32732),
            .I(N__32729));
    Span4Mux_h I__5880 (
            .O(N__32729),
            .I(N__32726));
    Span4Mux_h I__5879 (
            .O(N__32726),
            .I(N__32723));
    Odrv4 I__5878 (
            .O(N__32723),
            .I(sDAC_mem_11Z0Z_7));
    InMux I__5877 (
            .O(N__32720),
            .I(N__32717));
    LocalMux I__5876 (
            .O(N__32717),
            .I(sDAC_data_2_24_ns_1_10));
    CascadeMux I__5875 (
            .O(N__32714),
            .I(sDAC_data_RNO_8Z0Z_10_cascade_));
    InMux I__5874 (
            .O(N__32711),
            .I(N__32708));
    LocalMux I__5873 (
            .O(N__32708),
            .I(N__32705));
    Odrv4 I__5872 (
            .O(N__32705),
            .I(sDAC_data_RNO_7Z0Z_10));
    CascadeMux I__5871 (
            .O(N__32702),
            .I(sDAC_data_2_20_am_1_10_cascade_));
    InMux I__5870 (
            .O(N__32699),
            .I(N__32696));
    LocalMux I__5869 (
            .O(N__32696),
            .I(N__32693));
    Span4Mux_v I__5868 (
            .O(N__32693),
            .I(N__32690));
    Odrv4 I__5867 (
            .O(N__32690),
            .I(sDAC_mem_36Z0Z_6));
    CascadeMux I__5866 (
            .O(N__32687),
            .I(sDAC_data_2_13_am_1_9_cascade_));
    InMux I__5865 (
            .O(N__32684),
            .I(N__32681));
    LocalMux I__5864 (
            .O(N__32681),
            .I(N__32678));
    Span4Mux_h I__5863 (
            .O(N__32678),
            .I(N__32675));
    Odrv4 I__5862 (
            .O(N__32675),
            .I(sDAC_data_RNO_4Z0Z_9));
    CascadeMux I__5861 (
            .O(N__32672),
            .I(N__32669));
    InMux I__5860 (
            .O(N__32669),
            .I(N__32666));
    LocalMux I__5859 (
            .O(N__32666),
            .I(sDAC_mem_4Z0Z_6));
    InMux I__5858 (
            .O(N__32663),
            .I(N__32660));
    LocalMux I__5857 (
            .O(N__32660),
            .I(N__32657));
    Span4Mux_h I__5856 (
            .O(N__32657),
            .I(N__32654));
    Span4Mux_v I__5855 (
            .O(N__32654),
            .I(N__32651));
    Odrv4 I__5854 (
            .O(N__32651),
            .I(sDAC_mem_38Z0Z_7));
    InMux I__5853 (
            .O(N__32648),
            .I(N__32645));
    LocalMux I__5852 (
            .O(N__32645),
            .I(N__32642));
    Span4Mux_v I__5851 (
            .O(N__32642),
            .I(N__32639));
    Odrv4 I__5850 (
            .O(N__32639),
            .I(sDAC_mem_39Z0Z_7));
    CascadeMux I__5849 (
            .O(N__32636),
            .I(sDAC_data_2_13_bm_1_10_cascade_));
    InMux I__5848 (
            .O(N__32633),
            .I(N__32630));
    LocalMux I__5847 (
            .O(N__32630),
            .I(N__32627));
    Span4Mux_h I__5846 (
            .O(N__32627),
            .I(N__32624));
    Odrv4 I__5845 (
            .O(N__32624),
            .I(sDAC_mem_7Z0Z_7));
    InMux I__5844 (
            .O(N__32621),
            .I(N__32618));
    LocalMux I__5843 (
            .O(N__32618),
            .I(N__32615));
    Span4Mux_h I__5842 (
            .O(N__32615),
            .I(N__32612));
    Span4Mux_v I__5841 (
            .O(N__32612),
            .I(N__32609));
    Odrv4 I__5840 (
            .O(N__32609),
            .I(sDAC_mem_38Z0Z_0));
    InMux I__5839 (
            .O(N__32606),
            .I(N__32603));
    LocalMux I__5838 (
            .O(N__32603),
            .I(N__32600));
    Span4Mux_v I__5837 (
            .O(N__32600),
            .I(N__32597));
    Odrv4 I__5836 (
            .O(N__32597),
            .I(sDAC_mem_39Z0Z_0));
    CascadeMux I__5835 (
            .O(N__32594),
            .I(sDAC_data_2_13_bm_1_3_cascade_));
    InMux I__5834 (
            .O(N__32591),
            .I(N__32588));
    LocalMux I__5833 (
            .O(N__32588),
            .I(N__32585));
    Span12Mux_h I__5832 (
            .O(N__32585),
            .I(N__32582));
    Odrv12 I__5831 (
            .O(N__32582),
            .I(sDAC_mem_7Z0Z_0));
    InMux I__5830 (
            .O(N__32579),
            .I(N__32576));
    LocalMux I__5829 (
            .O(N__32576),
            .I(N__32573));
    Span4Mux_h I__5828 (
            .O(N__32573),
            .I(N__32570));
    Span4Mux_v I__5827 (
            .O(N__32570),
            .I(N__32567));
    Odrv4 I__5826 (
            .O(N__32567),
            .I(sDAC_mem_38Z0Z_1));
    InMux I__5825 (
            .O(N__32564),
            .I(N__32561));
    LocalMux I__5824 (
            .O(N__32561),
            .I(N__32558));
    Span4Mux_h I__5823 (
            .O(N__32558),
            .I(N__32555));
    Odrv4 I__5822 (
            .O(N__32555),
            .I(sDAC_data_2_13_bm_1_4));
    CascadeMux I__5821 (
            .O(N__32552),
            .I(sDAC_data_2_13_am_1_8_cascade_));
    InMux I__5820 (
            .O(N__32549),
            .I(N__32546));
    LocalMux I__5819 (
            .O(N__32546),
            .I(N__32543));
    Span4Mux_h I__5818 (
            .O(N__32543),
            .I(N__32540));
    Odrv4 I__5817 (
            .O(N__32540),
            .I(sDAC_data_RNO_4Z0Z_8));
    InMux I__5816 (
            .O(N__32537),
            .I(N__32534));
    LocalMux I__5815 (
            .O(N__32534),
            .I(N__32531));
    Span4Mux_h I__5814 (
            .O(N__32531),
            .I(N__32528));
    Span4Mux_h I__5813 (
            .O(N__32528),
            .I(N__32525));
    Odrv4 I__5812 (
            .O(N__32525),
            .I(sDAC_mem_38Z0Z_5));
    InMux I__5811 (
            .O(N__32522),
            .I(N__32519));
    LocalMux I__5810 (
            .O(N__32519),
            .I(N__32516));
    Odrv4 I__5809 (
            .O(N__32516),
            .I(sDAC_mem_39Z0Z_5));
    CascadeMux I__5808 (
            .O(N__32513),
            .I(sDAC_data_2_13_bm_1_8_cascade_));
    InMux I__5807 (
            .O(N__32510),
            .I(N__32507));
    LocalMux I__5806 (
            .O(N__32507),
            .I(N__32504));
    Span4Mux_h I__5805 (
            .O(N__32504),
            .I(N__32501));
    Odrv4 I__5804 (
            .O(N__32501),
            .I(sDAC_mem_7Z0Z_5));
    InMux I__5803 (
            .O(N__32498),
            .I(N__32495));
    LocalMux I__5802 (
            .O(N__32495),
            .I(N__32492));
    Span4Mux_v I__5801 (
            .O(N__32492),
            .I(N__32489));
    Odrv4 I__5800 (
            .O(N__32489),
            .I(sDAC_data_RNO_5Z0Z_8));
    InMux I__5799 (
            .O(N__32486),
            .I(N__32483));
    LocalMux I__5798 (
            .O(N__32483),
            .I(sDAC_mem_6Z0Z_5));
    InMux I__5797 (
            .O(N__32480),
            .I(N__32477));
    LocalMux I__5796 (
            .O(N__32477),
            .I(N__32474));
    Span4Mux_h I__5795 (
            .O(N__32474),
            .I(N__32471));
    Span4Mux_h I__5794 (
            .O(N__32471),
            .I(N__32468));
    Odrv4 I__5793 (
            .O(N__32468),
            .I(sDAC_mem_38Z0Z_6));
    CascadeMux I__5792 (
            .O(N__32465),
            .I(sDAC_data_2_13_bm_1_9_cascade_));
    InMux I__5791 (
            .O(N__32462),
            .I(N__32459));
    LocalMux I__5790 (
            .O(N__32459),
            .I(N__32456));
    Odrv12 I__5789 (
            .O(N__32456),
            .I(sDAC_mem_39Z0Z_6));
    InMux I__5788 (
            .O(N__32453),
            .I(N__32450));
    LocalMux I__5787 (
            .O(N__32450),
            .I(N__32447));
    Odrv4 I__5786 (
            .O(N__32447),
            .I(sDAC_data_RNO_5Z0Z_9));
    InMux I__5785 (
            .O(N__32444),
            .I(N__32441));
    LocalMux I__5784 (
            .O(N__32441),
            .I(sDAC_mem_6Z0Z_6));
    InMux I__5783 (
            .O(N__32438),
            .I(N__32435));
    LocalMux I__5782 (
            .O(N__32435),
            .I(N__32432));
    Span4Mux_h I__5781 (
            .O(N__32432),
            .I(N__32429));
    Span4Mux_v I__5780 (
            .O(N__32429),
            .I(N__32426));
    Odrv4 I__5779 (
            .O(N__32426),
            .I(sDAC_mem_40Z0Z_7));
    InMux I__5778 (
            .O(N__32423),
            .I(N__32420));
    LocalMux I__5777 (
            .O(N__32420),
            .I(N__32417));
    Span4Mux_v I__5776 (
            .O(N__32417),
            .I(N__32414));
    Span4Mux_h I__5775 (
            .O(N__32414),
            .I(N__32411));
    Odrv4 I__5774 (
            .O(N__32411),
            .I(sDAC_mem_8Z0Z_7));
    InMux I__5773 (
            .O(N__32408),
            .I(N__32405));
    LocalMux I__5772 (
            .O(N__32405),
            .I(N__32402));
    Sp12to4 I__5771 (
            .O(N__32402),
            .I(N__32399));
    Odrv12 I__5770 (
            .O(N__32399),
            .I(sDAC_mem_22Z0Z_0));
    InMux I__5769 (
            .O(N__32396),
            .I(N__32393));
    LocalMux I__5768 (
            .O(N__32393),
            .I(N__32390));
    Sp12to4 I__5767 (
            .O(N__32390),
            .I(N__32387));
    Odrv12 I__5766 (
            .O(N__32387),
            .I(sDAC_mem_22Z0Z_1));
    InMux I__5765 (
            .O(N__32384),
            .I(N__32381));
    LocalMux I__5764 (
            .O(N__32381),
            .I(sDAC_data_RNO_21Z0Z_4));
    InMux I__5763 (
            .O(N__32378),
            .I(N__32375));
    LocalMux I__5762 (
            .O(N__32375),
            .I(N__32372));
    Span12Mux_h I__5761 (
            .O(N__32372),
            .I(N__32369));
    Odrv12 I__5760 (
            .O(N__32369),
            .I(sDAC_mem_22Z0Z_2));
    InMux I__5759 (
            .O(N__32366),
            .I(N__32363));
    LocalMux I__5758 (
            .O(N__32363),
            .I(N__32360));
    Span12Mux_h I__5757 (
            .O(N__32360),
            .I(N__32357));
    Odrv12 I__5756 (
            .O(N__32357),
            .I(sDAC_mem_22Z0Z_3));
    InMux I__5755 (
            .O(N__32354),
            .I(N__32351));
    LocalMux I__5754 (
            .O(N__32351),
            .I(N__32348));
    Span4Mux_h I__5753 (
            .O(N__32348),
            .I(N__32345));
    Odrv4 I__5752 (
            .O(N__32345),
            .I(sDAC_data_RNO_21Z0Z_6));
    InMux I__5751 (
            .O(N__32342),
            .I(N__32339));
    LocalMux I__5750 (
            .O(N__32339),
            .I(N__32336));
    Span4Mux_v I__5749 (
            .O(N__32336),
            .I(N__32333));
    Odrv4 I__5748 (
            .O(N__32333),
            .I(sDAC_mem_36Z0Z_4));
    CascadeMux I__5747 (
            .O(N__32330),
            .I(sDAC_data_2_13_am_1_7_cascade_));
    InMux I__5746 (
            .O(N__32327),
            .I(N__32324));
    LocalMux I__5745 (
            .O(N__32324),
            .I(N__32321));
    Odrv4 I__5744 (
            .O(N__32321),
            .I(sDAC_data_RNO_4Z0Z_7));
    InMux I__5743 (
            .O(N__32318),
            .I(N__32315));
    LocalMux I__5742 (
            .O(N__32315),
            .I(sDAC_mem_4Z0Z_4));
    InMux I__5741 (
            .O(N__32312),
            .I(N__32309));
    LocalMux I__5740 (
            .O(N__32309),
            .I(N__32306));
    Span4Mux_v I__5739 (
            .O(N__32306),
            .I(N__32303));
    Odrv4 I__5738 (
            .O(N__32303),
            .I(sDAC_mem_36Z0Z_5));
    InMux I__5737 (
            .O(N__32300),
            .I(N__32297));
    LocalMux I__5736 (
            .O(N__32297),
            .I(N__32294));
    Odrv4 I__5735 (
            .O(N__32294),
            .I(sEEDACZ0Z_6));
    CascadeMux I__5734 (
            .O(N__32291),
            .I(sDAC_data_2_9_cascade_));
    InMux I__5733 (
            .O(N__32288),
            .I(N__32285));
    LocalMux I__5732 (
            .O(N__32285),
            .I(N__32282));
    Odrv4 I__5731 (
            .O(N__32282),
            .I(sDAC_dataZ0Z_9));
    InMux I__5730 (
            .O(N__32279),
            .I(N__32276));
    LocalMux I__5729 (
            .O(N__32276),
            .I(sDAC_data_2_14_ns_1_9));
    InMux I__5728 (
            .O(N__32273),
            .I(N__32270));
    LocalMux I__5727 (
            .O(N__32270),
            .I(N__32267));
    Odrv4 I__5726 (
            .O(N__32267),
            .I(sDAC_data_RNO_29Z0Z_9));
    InMux I__5725 (
            .O(N__32264),
            .I(N__32261));
    LocalMux I__5724 (
            .O(N__32261),
            .I(sDAC_data_RNO_28Z0Z_9));
    CascadeMux I__5723 (
            .O(N__32258),
            .I(sDAC_data_2_32_ns_1_9_cascade_));
    CascadeMux I__5722 (
            .O(N__32255),
            .I(sDAC_data_RNO_10Z0Z_9_cascade_));
    InMux I__5721 (
            .O(N__32252),
            .I(N__32249));
    LocalMux I__5720 (
            .O(N__32249),
            .I(N__32246));
    Span4Mux_h I__5719 (
            .O(N__32246),
            .I(N__32243));
    Span4Mux_v I__5718 (
            .O(N__32243),
            .I(N__32240));
    Odrv4 I__5717 (
            .O(N__32240),
            .I(sDAC_data_RNO_11Z0Z_9));
    InMux I__5716 (
            .O(N__32237),
            .I(N__32234));
    LocalMux I__5715 (
            .O(N__32234),
            .I(sDAC_data_2_41_ns_1_9));
    InMux I__5714 (
            .O(N__32231),
            .I(N__32228));
    LocalMux I__5713 (
            .O(N__32228),
            .I(N__32225));
    Odrv4 I__5712 (
            .O(N__32225),
            .I(sDAC_data_RNO_20Z0Z_8));
    InMux I__5711 (
            .O(N__32222),
            .I(N__32219));
    LocalMux I__5710 (
            .O(N__32219),
            .I(sDAC_mem_20Z0Z_5));
    InMux I__5709 (
            .O(N__32216),
            .I(N__32213));
    LocalMux I__5708 (
            .O(N__32213),
            .I(sDAC_data_RNO_20Z0Z_9));
    InMux I__5707 (
            .O(N__32210),
            .I(N__32207));
    LocalMux I__5706 (
            .O(N__32207),
            .I(sDAC_mem_20Z0Z_6));
    InMux I__5705 (
            .O(N__32204),
            .I(N__32201));
    LocalMux I__5704 (
            .O(N__32201),
            .I(sDAC_data_RNO_29Z0Z_7));
    InMux I__5703 (
            .O(N__32198),
            .I(N__32195));
    LocalMux I__5702 (
            .O(N__32195),
            .I(N__32192));
    Odrv4 I__5701 (
            .O(N__32192),
            .I(sDAC_data_RNO_28Z0Z_7));
    InMux I__5700 (
            .O(N__32189),
            .I(N__32186));
    LocalMux I__5699 (
            .O(N__32186),
            .I(sDAC_data_2_32_ns_1_7));
    CascadeMux I__5698 (
            .O(N__32183),
            .I(sDAC_data_2_14_ns_1_7_cascade_));
    InMux I__5697 (
            .O(N__32180),
            .I(N__32177));
    LocalMux I__5696 (
            .O(N__32177),
            .I(sDAC_data_RNO_5Z0Z_7));
    InMux I__5695 (
            .O(N__32174),
            .I(N__32171));
    LocalMux I__5694 (
            .O(N__32171),
            .I(N__32168));
    Span4Mux_v I__5693 (
            .O(N__32168),
            .I(N__32165));
    Span4Mux_v I__5692 (
            .O(N__32165),
            .I(N__32162));
    Odrv4 I__5691 (
            .O(N__32162),
            .I(sDAC_data_RNO_11Z0Z_7));
    InMux I__5690 (
            .O(N__32159),
            .I(N__32156));
    LocalMux I__5689 (
            .O(N__32156),
            .I(sDAC_data_RNO_10Z0Z_7));
    CascadeMux I__5688 (
            .O(N__32153),
            .I(sDAC_data_2_41_ns_1_7_cascade_));
    InMux I__5687 (
            .O(N__32150),
            .I(N__32147));
    LocalMux I__5686 (
            .O(N__32147),
            .I(sDAC_data_RNO_1Z0Z_7));
    InMux I__5685 (
            .O(N__32144),
            .I(N__32141));
    LocalMux I__5684 (
            .O(N__32141),
            .I(N__32138));
    Odrv4 I__5683 (
            .O(N__32138),
            .I(sEEDACZ0Z_4));
    CascadeMux I__5682 (
            .O(N__32135),
            .I(sDAC_data_2_7_cascade_));
    InMux I__5681 (
            .O(N__32132),
            .I(N__32129));
    LocalMux I__5680 (
            .O(N__32129),
            .I(N__32126));
    Odrv4 I__5679 (
            .O(N__32126),
            .I(sDAC_dataZ0Z_7));
    CascadeMux I__5678 (
            .O(N__32123),
            .I(sDAC_data_RNO_1Z0Z_9_cascade_));
    InMux I__5677 (
            .O(N__32120),
            .I(N__32117));
    LocalMux I__5676 (
            .O(N__32117),
            .I(N__32114));
    Odrv4 I__5675 (
            .O(N__32114),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_9 ));
    InMux I__5674 (
            .O(N__32111),
            .I(N__32108));
    LocalMux I__5673 (
            .O(N__32108),
            .I(N__32105));
    Span4Mux_v I__5672 (
            .O(N__32105),
            .I(N__32102));
    Odrv4 I__5671 (
            .O(N__32102),
            .I(sEEDACZ0Z_1));
    InMux I__5670 (
            .O(N__32099),
            .I(N__32096));
    LocalMux I__5669 (
            .O(N__32096),
            .I(N__32093));
    Span4Mux_h I__5668 (
            .O(N__32093),
            .I(N__32090));
    Odrv4 I__5667 (
            .O(N__32090),
            .I(sEEDACZ0Z_3));
    InMux I__5666 (
            .O(N__32087),
            .I(N__32084));
    LocalMux I__5665 (
            .O(N__32084),
            .I(N__32081));
    Span4Mux_v I__5664 (
            .O(N__32081),
            .I(N__32078));
    Span4Mux_h I__5663 (
            .O(N__32078),
            .I(N__32075));
    Odrv4 I__5662 (
            .O(N__32075),
            .I(sEEDACZ0Z_5));
    InMux I__5661 (
            .O(N__32072),
            .I(N__32069));
    LocalMux I__5660 (
            .O(N__32069),
            .I(N__32066));
    Span4Mux_v I__5659 (
            .O(N__32066),
            .I(N__32063));
    Span4Mux_v I__5658 (
            .O(N__32063),
            .I(N__32060));
    Odrv4 I__5657 (
            .O(N__32060),
            .I(sEEDACZ0Z_7));
    CEMux I__5656 (
            .O(N__32057),
            .I(N__32054));
    LocalMux I__5655 (
            .O(N__32054),
            .I(N__32051));
    Odrv4 I__5654 (
            .O(N__32051),
            .I(sEEDAC_1_sqmuxa));
    CascadeMux I__5653 (
            .O(N__32048),
            .I(N__32042));
    CascadeMux I__5652 (
            .O(N__32047),
            .I(N__32038));
    InMux I__5651 (
            .O(N__32046),
            .I(N__32034));
    InMux I__5650 (
            .O(N__32045),
            .I(N__32031));
    InMux I__5649 (
            .O(N__32042),
            .I(N__32028));
    CascadeMux I__5648 (
            .O(N__32041),
            .I(N__32024));
    InMux I__5647 (
            .O(N__32038),
            .I(N__32021));
    InMux I__5646 (
            .O(N__32037),
            .I(N__32015));
    LocalMux I__5645 (
            .O(N__32034),
            .I(N__32010));
    LocalMux I__5644 (
            .O(N__32031),
            .I(N__32010));
    LocalMux I__5643 (
            .O(N__32028),
            .I(N__32007));
    InMux I__5642 (
            .O(N__32027),
            .I(N__32004));
    InMux I__5641 (
            .O(N__32024),
            .I(N__32001));
    LocalMux I__5640 (
            .O(N__32021),
            .I(N__31998));
    InMux I__5639 (
            .O(N__32020),
            .I(N__31995));
    InMux I__5638 (
            .O(N__32019),
            .I(N__31992));
    InMux I__5637 (
            .O(N__32018),
            .I(N__31987));
    LocalMux I__5636 (
            .O(N__32015),
            .I(N__31984));
    Span4Mux_v I__5635 (
            .O(N__32010),
            .I(N__31981));
    Span4Mux_v I__5634 (
            .O(N__32007),
            .I(N__31976));
    LocalMux I__5633 (
            .O(N__32004),
            .I(N__31976));
    LocalMux I__5632 (
            .O(N__32001),
            .I(N__31973));
    Span4Mux_h I__5631 (
            .O(N__31998),
            .I(N__31966));
    LocalMux I__5630 (
            .O(N__31995),
            .I(N__31966));
    LocalMux I__5629 (
            .O(N__31992),
            .I(N__31966));
    InMux I__5628 (
            .O(N__31991),
            .I(N__31963));
    InMux I__5627 (
            .O(N__31990),
            .I(N__31960));
    LocalMux I__5626 (
            .O(N__31987),
            .I(N__31951));
    Span4Mux_h I__5625 (
            .O(N__31984),
            .I(N__31951));
    Span4Mux_h I__5624 (
            .O(N__31981),
            .I(N__31951));
    Span4Mux_v I__5623 (
            .O(N__31976),
            .I(N__31951));
    Span4Mux_v I__5622 (
            .O(N__31973),
            .I(N__31946));
    Span4Mux_v I__5621 (
            .O(N__31966),
            .I(N__31946));
    LocalMux I__5620 (
            .O(N__31963),
            .I(un7_spon_22));
    LocalMux I__5619 (
            .O(N__31960),
            .I(un7_spon_22));
    Odrv4 I__5618 (
            .O(N__31951),
            .I(un7_spon_22));
    Odrv4 I__5617 (
            .O(N__31946),
            .I(un7_spon_22));
    CascadeMux I__5616 (
            .O(N__31937),
            .I(N__31931));
    CascadeMux I__5615 (
            .O(N__31936),
            .I(N__31926));
    CascadeMux I__5614 (
            .O(N__31935),
            .I(N__31923));
    InMux I__5613 (
            .O(N__31934),
            .I(N__31920));
    InMux I__5612 (
            .O(N__31931),
            .I(N__31917));
    CascadeMux I__5611 (
            .O(N__31930),
            .I(N__31914));
    InMux I__5610 (
            .O(N__31929),
            .I(N__31910));
    InMux I__5609 (
            .O(N__31926),
            .I(N__31906));
    InMux I__5608 (
            .O(N__31923),
            .I(N__31902));
    LocalMux I__5607 (
            .O(N__31920),
            .I(N__31899));
    LocalMux I__5606 (
            .O(N__31917),
            .I(N__31896));
    InMux I__5605 (
            .O(N__31914),
            .I(N__31893));
    InMux I__5604 (
            .O(N__31913),
            .I(N__31890));
    LocalMux I__5603 (
            .O(N__31910),
            .I(N__31887));
    InMux I__5602 (
            .O(N__31909),
            .I(N__31884));
    LocalMux I__5601 (
            .O(N__31906),
            .I(N__31879));
    CascadeMux I__5600 (
            .O(N__31905),
            .I(N__31876));
    LocalMux I__5599 (
            .O(N__31902),
            .I(N__31873));
    Span4Mux_v I__5598 (
            .O(N__31899),
            .I(N__31866));
    Span4Mux_h I__5597 (
            .O(N__31896),
            .I(N__31866));
    LocalMux I__5596 (
            .O(N__31893),
            .I(N__31866));
    LocalMux I__5595 (
            .O(N__31890),
            .I(N__31863));
    Span4Mux_h I__5594 (
            .O(N__31887),
            .I(N__31858));
    LocalMux I__5593 (
            .O(N__31884),
            .I(N__31858));
    InMux I__5592 (
            .O(N__31883),
            .I(N__31855));
    InMux I__5591 (
            .O(N__31882),
            .I(N__31852));
    Span4Mux_h I__5590 (
            .O(N__31879),
            .I(N__31849));
    InMux I__5589 (
            .O(N__31876),
            .I(N__31846));
    Span4Mux_v I__5588 (
            .O(N__31873),
            .I(N__31843));
    Span4Mux_v I__5587 (
            .O(N__31866),
            .I(N__31838));
    Span4Mux_v I__5586 (
            .O(N__31863),
            .I(N__31838));
    Span4Mux_v I__5585 (
            .O(N__31858),
            .I(N__31835));
    LocalMux I__5584 (
            .O(N__31855),
            .I(un7_spon_23));
    LocalMux I__5583 (
            .O(N__31852),
            .I(un7_spon_23));
    Odrv4 I__5582 (
            .O(N__31849),
            .I(un7_spon_23));
    LocalMux I__5581 (
            .O(N__31846),
            .I(un7_spon_23));
    Odrv4 I__5580 (
            .O(N__31843),
            .I(un7_spon_23));
    Odrv4 I__5579 (
            .O(N__31838),
            .I(un7_spon_23));
    Odrv4 I__5578 (
            .O(N__31835),
            .I(un7_spon_23));
    InMux I__5577 (
            .O(N__31820),
            .I(bfn_14_20_0_));
    InMux I__5576 (
            .O(N__31817),
            .I(N__31814));
    LocalMux I__5575 (
            .O(N__31814),
            .I(N__31811));
    Span4Mux_v I__5574 (
            .O(N__31811),
            .I(N__31808));
    Span4Mux_v I__5573 (
            .O(N__31808),
            .I(N__31805));
    Odrv4 I__5572 (
            .O(N__31805),
            .I(un4_spoff_cry_23_THRU_CO));
    InMux I__5571 (
            .O(N__31802),
            .I(N__31799));
    LocalMux I__5570 (
            .O(N__31799),
            .I(N__31796));
    Odrv12 I__5569 (
            .O(N__31796),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_3 ));
    InMux I__5568 (
            .O(N__31793),
            .I(N__31790));
    LocalMux I__5567 (
            .O(N__31790),
            .I(N__31787));
    Span4Mux_h I__5566 (
            .O(N__31787),
            .I(N__31784));
    Span4Mux_v I__5565 (
            .O(N__31784),
            .I(N__31781));
    Odrv4 I__5564 (
            .O(N__31781),
            .I(sDAC_dataZ0Z_4));
    InMux I__5563 (
            .O(N__31778),
            .I(N__31775));
    LocalMux I__5562 (
            .O(N__31775),
            .I(N__31772));
    Odrv12 I__5561 (
            .O(N__31772),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_4 ));
    InMux I__5560 (
            .O(N__31769),
            .I(N__31766));
    LocalMux I__5559 (
            .O(N__31766),
            .I(N__31763));
    Odrv4 I__5558 (
            .O(N__31763),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_7 ));
    InMux I__5557 (
            .O(N__31760),
            .I(N__31757));
    LocalMux I__5556 (
            .O(N__31757),
            .I(N__31754));
    Span4Mux_h I__5555 (
            .O(N__31754),
            .I(N__31751));
    Odrv4 I__5554 (
            .O(N__31751),
            .I(sDAC_dataZ0Z_8));
    CascadeMux I__5553 (
            .O(N__31748),
            .I(N__31744));
    InMux I__5552 (
            .O(N__31747),
            .I(N__31740));
    InMux I__5551 (
            .O(N__31744),
            .I(N__31737));
    CascadeMux I__5550 (
            .O(N__31743),
            .I(N__31734));
    LocalMux I__5549 (
            .O(N__31740),
            .I(N__31729));
    LocalMux I__5548 (
            .O(N__31737),
            .I(N__31726));
    InMux I__5547 (
            .O(N__31734),
            .I(N__31723));
    CascadeMux I__5546 (
            .O(N__31733),
            .I(N__31719));
    InMux I__5545 (
            .O(N__31732),
            .I(N__31714));
    Span4Mux_h I__5544 (
            .O(N__31729),
            .I(N__31707));
    Span4Mux_h I__5543 (
            .O(N__31726),
            .I(N__31707));
    LocalMux I__5542 (
            .O(N__31723),
            .I(N__31707));
    InMux I__5541 (
            .O(N__31722),
            .I(N__31704));
    InMux I__5540 (
            .O(N__31719),
            .I(N__31701));
    InMux I__5539 (
            .O(N__31718),
            .I(N__31697));
    InMux I__5538 (
            .O(N__31717),
            .I(N__31694));
    LocalMux I__5537 (
            .O(N__31714),
            .I(N__31691));
    Span4Mux_v I__5536 (
            .O(N__31707),
            .I(N__31688));
    LocalMux I__5535 (
            .O(N__31704),
            .I(N__31685));
    LocalMux I__5534 (
            .O(N__31701),
            .I(N__31682));
    InMux I__5533 (
            .O(N__31700),
            .I(N__31679));
    LocalMux I__5532 (
            .O(N__31697),
            .I(un7_spon_12));
    LocalMux I__5531 (
            .O(N__31694),
            .I(un7_spon_12));
    Odrv12 I__5530 (
            .O(N__31691),
            .I(un7_spon_12));
    Odrv4 I__5529 (
            .O(N__31688),
            .I(un7_spon_12));
    Odrv4 I__5528 (
            .O(N__31685),
            .I(un7_spon_12));
    Odrv12 I__5527 (
            .O(N__31682),
            .I(un7_spon_12));
    LocalMux I__5526 (
            .O(N__31679),
            .I(un7_spon_12));
    CascadeMux I__5525 (
            .O(N__31664),
            .I(N__31661));
    InMux I__5524 (
            .O(N__31661),
            .I(N__31655));
    InMux I__5523 (
            .O(N__31660),
            .I(N__31652));
    CascadeMux I__5522 (
            .O(N__31659),
            .I(N__31649));
    CascadeMux I__5521 (
            .O(N__31658),
            .I(N__31646));
    LocalMux I__5520 (
            .O(N__31655),
            .I(N__31640));
    LocalMux I__5519 (
            .O(N__31652),
            .I(N__31637));
    InMux I__5518 (
            .O(N__31649),
            .I(N__31634));
    InMux I__5517 (
            .O(N__31646),
            .I(N__31631));
    InMux I__5516 (
            .O(N__31645),
            .I(N__31627));
    InMux I__5515 (
            .O(N__31644),
            .I(N__31624));
    InMux I__5514 (
            .O(N__31643),
            .I(N__31621));
    Span4Mux_h I__5513 (
            .O(N__31640),
            .I(N__31614));
    Span4Mux_h I__5512 (
            .O(N__31637),
            .I(N__31614));
    LocalMux I__5511 (
            .O(N__31634),
            .I(N__31614));
    LocalMux I__5510 (
            .O(N__31631),
            .I(N__31611));
    InMux I__5509 (
            .O(N__31630),
            .I(N__31607));
    LocalMux I__5508 (
            .O(N__31627),
            .I(N__31602));
    LocalMux I__5507 (
            .O(N__31624),
            .I(N__31602));
    LocalMux I__5506 (
            .O(N__31621),
            .I(N__31599));
    Span4Mux_v I__5505 (
            .O(N__31614),
            .I(N__31594));
    Span4Mux_v I__5504 (
            .O(N__31611),
            .I(N__31594));
    InMux I__5503 (
            .O(N__31610),
            .I(N__31591));
    LocalMux I__5502 (
            .O(N__31607),
            .I(un7_spon_13));
    Odrv12 I__5501 (
            .O(N__31602),
            .I(un7_spon_13));
    Odrv4 I__5500 (
            .O(N__31599),
            .I(un7_spon_13));
    Odrv4 I__5499 (
            .O(N__31594),
            .I(un7_spon_13));
    LocalMux I__5498 (
            .O(N__31591),
            .I(un7_spon_13));
    CascadeMux I__5497 (
            .O(N__31580),
            .I(N__31575));
    CascadeMux I__5496 (
            .O(N__31579),
            .I(N__31570));
    InMux I__5495 (
            .O(N__31578),
            .I(N__31566));
    InMux I__5494 (
            .O(N__31575),
            .I(N__31563));
    CascadeMux I__5493 (
            .O(N__31574),
            .I(N__31560));
    CascadeMux I__5492 (
            .O(N__31573),
            .I(N__31557));
    InMux I__5491 (
            .O(N__31570),
            .I(N__31554));
    InMux I__5490 (
            .O(N__31569),
            .I(N__31551));
    LocalMux I__5489 (
            .O(N__31566),
            .I(N__31547));
    LocalMux I__5488 (
            .O(N__31563),
            .I(N__31544));
    InMux I__5487 (
            .O(N__31560),
            .I(N__31541));
    InMux I__5486 (
            .O(N__31557),
            .I(N__31538));
    LocalMux I__5485 (
            .O(N__31554),
            .I(N__31534));
    LocalMux I__5484 (
            .O(N__31551),
            .I(N__31531));
    InMux I__5483 (
            .O(N__31550),
            .I(N__31528));
    Span4Mux_h I__5482 (
            .O(N__31547),
            .I(N__31521));
    Span4Mux_h I__5481 (
            .O(N__31544),
            .I(N__31521));
    LocalMux I__5480 (
            .O(N__31541),
            .I(N__31521));
    LocalMux I__5479 (
            .O(N__31538),
            .I(N__31518));
    InMux I__5478 (
            .O(N__31537),
            .I(N__31514));
    Span4Mux_h I__5477 (
            .O(N__31534),
            .I(N__31511));
    Span4Mux_h I__5476 (
            .O(N__31531),
            .I(N__31508));
    LocalMux I__5475 (
            .O(N__31528),
            .I(N__31505));
    Span4Mux_v I__5474 (
            .O(N__31521),
            .I(N__31500));
    Span4Mux_v I__5473 (
            .O(N__31518),
            .I(N__31500));
    InMux I__5472 (
            .O(N__31517),
            .I(N__31497));
    LocalMux I__5471 (
            .O(N__31514),
            .I(un7_spon_14));
    Odrv4 I__5470 (
            .O(N__31511),
            .I(un7_spon_14));
    Odrv4 I__5469 (
            .O(N__31508),
            .I(un7_spon_14));
    Odrv4 I__5468 (
            .O(N__31505),
            .I(un7_spon_14));
    Odrv4 I__5467 (
            .O(N__31500),
            .I(un7_spon_14));
    LocalMux I__5466 (
            .O(N__31497),
            .I(un7_spon_14));
    CascadeMux I__5465 (
            .O(N__31484),
            .I(N__31481));
    InMux I__5464 (
            .O(N__31481),
            .I(N__31476));
    InMux I__5463 (
            .O(N__31480),
            .I(N__31473));
    CascadeMux I__5462 (
            .O(N__31479),
            .I(N__31469));
    LocalMux I__5461 (
            .O(N__31476),
            .I(N__31464));
    LocalMux I__5460 (
            .O(N__31473),
            .I(N__31461));
    InMux I__5459 (
            .O(N__31472),
            .I(N__31458));
    InMux I__5458 (
            .O(N__31469),
            .I(N__31455));
    CascadeMux I__5457 (
            .O(N__31468),
            .I(N__31451));
    CascadeMux I__5456 (
            .O(N__31467),
            .I(N__31447));
    Span4Mux_h I__5455 (
            .O(N__31464),
            .I(N__31440));
    Span4Mux_h I__5454 (
            .O(N__31461),
            .I(N__31440));
    LocalMux I__5453 (
            .O(N__31458),
            .I(N__31440));
    LocalMux I__5452 (
            .O(N__31455),
            .I(N__31437));
    InMux I__5451 (
            .O(N__31454),
            .I(N__31434));
    InMux I__5450 (
            .O(N__31451),
            .I(N__31431));
    InMux I__5449 (
            .O(N__31450),
            .I(N__31427));
    InMux I__5448 (
            .O(N__31447),
            .I(N__31424));
    Span4Mux_v I__5447 (
            .O(N__31440),
            .I(N__31421));
    Span4Mux_v I__5446 (
            .O(N__31437),
            .I(N__31418));
    LocalMux I__5445 (
            .O(N__31434),
            .I(N__31413));
    LocalMux I__5444 (
            .O(N__31431),
            .I(N__31413));
    InMux I__5443 (
            .O(N__31430),
            .I(N__31410));
    LocalMux I__5442 (
            .O(N__31427),
            .I(un7_spon_15));
    LocalMux I__5441 (
            .O(N__31424),
            .I(un7_spon_15));
    Odrv4 I__5440 (
            .O(N__31421),
            .I(un7_spon_15));
    Odrv4 I__5439 (
            .O(N__31418),
            .I(un7_spon_15));
    Odrv12 I__5438 (
            .O(N__31413),
            .I(un7_spon_15));
    LocalMux I__5437 (
            .O(N__31410),
            .I(un7_spon_15));
    CascadeMux I__5436 (
            .O(N__31397),
            .I(N__31394));
    InMux I__5435 (
            .O(N__31394),
            .I(N__31390));
    CascadeMux I__5434 (
            .O(N__31393),
            .I(N__31384));
    LocalMux I__5433 (
            .O(N__31390),
            .I(N__31381));
    InMux I__5432 (
            .O(N__31389),
            .I(N__31378));
    InMux I__5431 (
            .O(N__31388),
            .I(N__31373));
    CascadeMux I__5430 (
            .O(N__31387),
            .I(N__31370));
    InMux I__5429 (
            .O(N__31384),
            .I(N__31367));
    Span4Mux_v I__5428 (
            .O(N__31381),
            .I(N__31362));
    LocalMux I__5427 (
            .O(N__31378),
            .I(N__31359));
    InMux I__5426 (
            .O(N__31377),
            .I(N__31354));
    InMux I__5425 (
            .O(N__31376),
            .I(N__31354));
    LocalMux I__5424 (
            .O(N__31373),
            .I(N__31351));
    InMux I__5423 (
            .O(N__31370),
            .I(N__31348));
    LocalMux I__5422 (
            .O(N__31367),
            .I(N__31345));
    InMux I__5421 (
            .O(N__31366),
            .I(N__31342));
    InMux I__5420 (
            .O(N__31365),
            .I(N__31339));
    Span4Mux_h I__5419 (
            .O(N__31362),
            .I(N__31327));
    Span4Mux_h I__5418 (
            .O(N__31359),
            .I(N__31327));
    LocalMux I__5417 (
            .O(N__31354),
            .I(N__31327));
    Span4Mux_v I__5416 (
            .O(N__31351),
            .I(N__31327));
    LocalMux I__5415 (
            .O(N__31348),
            .I(N__31324));
    Span4Mux_v I__5414 (
            .O(N__31345),
            .I(N__31319));
    LocalMux I__5413 (
            .O(N__31342),
            .I(N__31319));
    LocalMux I__5412 (
            .O(N__31339),
            .I(N__31316));
    InMux I__5411 (
            .O(N__31338),
            .I(N__31313));
    InMux I__5410 (
            .O(N__31337),
            .I(N__31310));
    InMux I__5409 (
            .O(N__31336),
            .I(N__31307));
    Span4Mux_v I__5408 (
            .O(N__31327),
            .I(N__31302));
    Span4Mux_h I__5407 (
            .O(N__31324),
            .I(N__31302));
    Span4Mux_v I__5406 (
            .O(N__31319),
            .I(N__31297));
    Span4Mux_v I__5405 (
            .O(N__31316),
            .I(N__31297));
    LocalMux I__5404 (
            .O(N__31313),
            .I(un7_spon_16));
    LocalMux I__5403 (
            .O(N__31310),
            .I(un7_spon_16));
    LocalMux I__5402 (
            .O(N__31307),
            .I(un7_spon_16));
    Odrv4 I__5401 (
            .O(N__31302),
            .I(un7_spon_16));
    Odrv4 I__5400 (
            .O(N__31297),
            .I(un7_spon_16));
    CascadeMux I__5399 (
            .O(N__31286),
            .I(N__31280));
    InMux I__5398 (
            .O(N__31285),
            .I(N__31277));
    CascadeMux I__5397 (
            .O(N__31284),
            .I(N__31273));
    InMux I__5396 (
            .O(N__31283),
            .I(N__31270));
    InMux I__5395 (
            .O(N__31280),
            .I(N__31263));
    LocalMux I__5394 (
            .O(N__31277),
            .I(N__31258));
    InMux I__5393 (
            .O(N__31276),
            .I(N__31255));
    InMux I__5392 (
            .O(N__31273),
            .I(N__31252));
    LocalMux I__5391 (
            .O(N__31270),
            .I(N__31249));
    InMux I__5390 (
            .O(N__31269),
            .I(N__31246));
    CascadeMux I__5389 (
            .O(N__31268),
            .I(N__31243));
    CascadeMux I__5388 (
            .O(N__31267),
            .I(N__31240));
    InMux I__5387 (
            .O(N__31266),
            .I(N__31236));
    LocalMux I__5386 (
            .O(N__31263),
            .I(N__31233));
    InMux I__5385 (
            .O(N__31262),
            .I(N__31230));
    InMux I__5384 (
            .O(N__31261),
            .I(N__31227));
    Span4Mux_v I__5383 (
            .O(N__31258),
            .I(N__31222));
    LocalMux I__5382 (
            .O(N__31255),
            .I(N__31222));
    LocalMux I__5381 (
            .O(N__31252),
            .I(N__31219));
    Span4Mux_v I__5380 (
            .O(N__31249),
            .I(N__31214));
    LocalMux I__5379 (
            .O(N__31246),
            .I(N__31214));
    InMux I__5378 (
            .O(N__31243),
            .I(N__31211));
    InMux I__5377 (
            .O(N__31240),
            .I(N__31206));
    InMux I__5376 (
            .O(N__31239),
            .I(N__31206));
    LocalMux I__5375 (
            .O(N__31236),
            .I(N__31203));
    Span4Mux_v I__5374 (
            .O(N__31233),
            .I(N__31200));
    LocalMux I__5373 (
            .O(N__31230),
            .I(N__31189));
    LocalMux I__5372 (
            .O(N__31227),
            .I(N__31189));
    Span4Mux_v I__5371 (
            .O(N__31222),
            .I(N__31189));
    Span4Mux_h I__5370 (
            .O(N__31219),
            .I(N__31189));
    Span4Mux_v I__5369 (
            .O(N__31214),
            .I(N__31189));
    LocalMux I__5368 (
            .O(N__31211),
            .I(un7_spon_17));
    LocalMux I__5367 (
            .O(N__31206),
            .I(un7_spon_17));
    Odrv12 I__5366 (
            .O(N__31203),
            .I(un7_spon_17));
    Odrv4 I__5365 (
            .O(N__31200),
            .I(un7_spon_17));
    Odrv4 I__5364 (
            .O(N__31189),
            .I(un7_spon_17));
    CascadeMux I__5363 (
            .O(N__31178),
            .I(N__31173));
    CascadeMux I__5362 (
            .O(N__31177),
            .I(N__31170));
    CascadeMux I__5361 (
            .O(N__31176),
            .I(N__31167));
    InMux I__5360 (
            .O(N__31173),
            .I(N__31164));
    InMux I__5359 (
            .O(N__31170),
            .I(N__31157));
    InMux I__5358 (
            .O(N__31167),
            .I(N__31154));
    LocalMux I__5357 (
            .O(N__31164),
            .I(N__31151));
    InMux I__5356 (
            .O(N__31163),
            .I(N__31145));
    InMux I__5355 (
            .O(N__31162),
            .I(N__31142));
    InMux I__5354 (
            .O(N__31161),
            .I(N__31137));
    InMux I__5353 (
            .O(N__31160),
            .I(N__31137));
    LocalMux I__5352 (
            .O(N__31157),
            .I(N__31134));
    LocalMux I__5351 (
            .O(N__31154),
            .I(N__31131));
    Span4Mux_v I__5350 (
            .O(N__31151),
            .I(N__31128));
    InMux I__5349 (
            .O(N__31150),
            .I(N__31125));
    InMux I__5348 (
            .O(N__31149),
            .I(N__31120));
    InMux I__5347 (
            .O(N__31148),
            .I(N__31117));
    LocalMux I__5346 (
            .O(N__31145),
            .I(N__31114));
    LocalMux I__5345 (
            .O(N__31142),
            .I(N__31111));
    LocalMux I__5344 (
            .O(N__31137),
            .I(N__31108));
    Span4Mux_h I__5343 (
            .O(N__31134),
            .I(N__31105));
    Span4Mux_v I__5342 (
            .O(N__31131),
            .I(N__31098));
    Span4Mux_h I__5341 (
            .O(N__31128),
            .I(N__31098));
    LocalMux I__5340 (
            .O(N__31125),
            .I(N__31098));
    InMux I__5339 (
            .O(N__31124),
            .I(N__31095));
    InMux I__5338 (
            .O(N__31123),
            .I(N__31092));
    LocalMux I__5337 (
            .O(N__31120),
            .I(N__31089));
    LocalMux I__5336 (
            .O(N__31117),
            .I(N__31076));
    Span4Mux_h I__5335 (
            .O(N__31114),
            .I(N__31076));
    Span4Mux_h I__5334 (
            .O(N__31111),
            .I(N__31076));
    Span4Mux_v I__5333 (
            .O(N__31108),
            .I(N__31076));
    Span4Mux_v I__5332 (
            .O(N__31105),
            .I(N__31076));
    Span4Mux_v I__5331 (
            .O(N__31098),
            .I(N__31076));
    LocalMux I__5330 (
            .O(N__31095),
            .I(un7_spon_18));
    LocalMux I__5329 (
            .O(N__31092),
            .I(un7_spon_18));
    Odrv12 I__5328 (
            .O(N__31089),
            .I(un7_spon_18));
    Odrv4 I__5327 (
            .O(N__31076),
            .I(un7_spon_18));
    InMux I__5326 (
            .O(N__31067),
            .I(N__31064));
    LocalMux I__5325 (
            .O(N__31064),
            .I(sEEPonPoffZ0Z_4));
    CascadeMux I__5324 (
            .O(N__31061),
            .I(N__31056));
    CascadeMux I__5323 (
            .O(N__31060),
            .I(N__31053));
    InMux I__5322 (
            .O(N__31059),
            .I(N__31049));
    InMux I__5321 (
            .O(N__31056),
            .I(N__31045));
    InMux I__5320 (
            .O(N__31053),
            .I(N__31042));
    CascadeMux I__5319 (
            .O(N__31052),
            .I(N__31039));
    LocalMux I__5318 (
            .O(N__31049),
            .I(N__31035));
    CascadeMux I__5317 (
            .O(N__31048),
            .I(N__31030));
    LocalMux I__5316 (
            .O(N__31045),
            .I(N__31026));
    LocalMux I__5315 (
            .O(N__31042),
            .I(N__31023));
    InMux I__5314 (
            .O(N__31039),
            .I(N__31020));
    CascadeMux I__5313 (
            .O(N__31038),
            .I(N__31017));
    Span4Mux_v I__5312 (
            .O(N__31035),
            .I(N__31013));
    InMux I__5311 (
            .O(N__31034),
            .I(N__31008));
    InMux I__5310 (
            .O(N__31033),
            .I(N__31008));
    InMux I__5309 (
            .O(N__31030),
            .I(N__31005));
    InMux I__5308 (
            .O(N__31029),
            .I(N__31002));
    Span4Mux_h I__5307 (
            .O(N__31026),
            .I(N__30996));
    Span4Mux_v I__5306 (
            .O(N__31023),
            .I(N__30991));
    LocalMux I__5305 (
            .O(N__31020),
            .I(N__30991));
    InMux I__5304 (
            .O(N__31017),
            .I(N__30988));
    CascadeMux I__5303 (
            .O(N__31016),
            .I(N__30985));
    Span4Mux_v I__5302 (
            .O(N__31013),
            .I(N__30975));
    LocalMux I__5301 (
            .O(N__31008),
            .I(N__30975));
    LocalMux I__5300 (
            .O(N__31005),
            .I(N__30975));
    LocalMux I__5299 (
            .O(N__31002),
            .I(N__30975));
    InMux I__5298 (
            .O(N__31001),
            .I(N__30972));
    InMux I__5297 (
            .O(N__31000),
            .I(N__30969));
    InMux I__5296 (
            .O(N__30999),
            .I(N__30966));
    Span4Mux_v I__5295 (
            .O(N__30996),
            .I(N__30959));
    Span4Mux_h I__5294 (
            .O(N__30991),
            .I(N__30959));
    LocalMux I__5293 (
            .O(N__30988),
            .I(N__30959));
    InMux I__5292 (
            .O(N__30985),
            .I(N__30956));
    InMux I__5291 (
            .O(N__30984),
            .I(N__30952));
    Span4Mux_v I__5290 (
            .O(N__30975),
            .I(N__30949));
    LocalMux I__5289 (
            .O(N__30972),
            .I(N__30946));
    LocalMux I__5288 (
            .O(N__30969),
            .I(N__30939));
    LocalMux I__5287 (
            .O(N__30966),
            .I(N__30939));
    Span4Mux_v I__5286 (
            .O(N__30959),
            .I(N__30939));
    LocalMux I__5285 (
            .O(N__30956),
            .I(N__30936));
    InMux I__5284 (
            .O(N__30955),
            .I(N__30933));
    LocalMux I__5283 (
            .O(N__30952),
            .I(un7_spon_4));
    Odrv4 I__5282 (
            .O(N__30949),
            .I(un7_spon_4));
    Odrv12 I__5281 (
            .O(N__30946),
            .I(un7_spon_4));
    Odrv4 I__5280 (
            .O(N__30939),
            .I(un7_spon_4));
    Odrv12 I__5279 (
            .O(N__30936),
            .I(un7_spon_4));
    LocalMux I__5278 (
            .O(N__30933),
            .I(un7_spon_4));
    InMux I__5277 (
            .O(N__30920),
            .I(N__30917));
    LocalMux I__5276 (
            .O(N__30917),
            .I(sEEPonPoff_i_4));
    InMux I__5275 (
            .O(N__30914),
            .I(N__30911));
    LocalMux I__5274 (
            .O(N__30911),
            .I(sEEPonPoffZ0Z_5));
    CascadeMux I__5273 (
            .O(N__30908),
            .I(N__30904));
    CascadeMux I__5272 (
            .O(N__30907),
            .I(N__30901));
    InMux I__5271 (
            .O(N__30904),
            .I(N__30895));
    InMux I__5270 (
            .O(N__30901),
            .I(N__30892));
    CascadeMux I__5269 (
            .O(N__30900),
            .I(N__30889));
    CascadeMux I__5268 (
            .O(N__30899),
            .I(N__30885));
    InMux I__5267 (
            .O(N__30898),
            .I(N__30882));
    LocalMux I__5266 (
            .O(N__30895),
            .I(N__30876));
    LocalMux I__5265 (
            .O(N__30892),
            .I(N__30873));
    InMux I__5264 (
            .O(N__30889),
            .I(N__30870));
    InMux I__5263 (
            .O(N__30888),
            .I(N__30867));
    InMux I__5262 (
            .O(N__30885),
            .I(N__30864));
    LocalMux I__5261 (
            .O(N__30882),
            .I(N__30860));
    InMux I__5260 (
            .O(N__30881),
            .I(N__30857));
    InMux I__5259 (
            .O(N__30880),
            .I(N__30852));
    InMux I__5258 (
            .O(N__30879),
            .I(N__30852));
    Span4Mux_h I__5257 (
            .O(N__30876),
            .I(N__30845));
    Span4Mux_h I__5256 (
            .O(N__30873),
            .I(N__30845));
    LocalMux I__5255 (
            .O(N__30870),
            .I(N__30845));
    LocalMux I__5254 (
            .O(N__30867),
            .I(N__30842));
    LocalMux I__5253 (
            .O(N__30864),
            .I(N__30839));
    InMux I__5252 (
            .O(N__30863),
            .I(N__30835));
    Span4Mux_h I__5251 (
            .O(N__30860),
            .I(N__30832));
    LocalMux I__5250 (
            .O(N__30857),
            .I(N__30829));
    LocalMux I__5249 (
            .O(N__30852),
            .I(N__30824));
    Span4Mux_v I__5248 (
            .O(N__30845),
            .I(N__30824));
    Span4Mux_h I__5247 (
            .O(N__30842),
            .I(N__30819));
    Span4Mux_v I__5246 (
            .O(N__30839),
            .I(N__30819));
    InMux I__5245 (
            .O(N__30838),
            .I(N__30816));
    LocalMux I__5244 (
            .O(N__30835),
            .I(un7_spon_5));
    Odrv4 I__5243 (
            .O(N__30832),
            .I(un7_spon_5));
    Odrv4 I__5242 (
            .O(N__30829),
            .I(un7_spon_5));
    Odrv4 I__5241 (
            .O(N__30824),
            .I(un7_spon_5));
    Odrv4 I__5240 (
            .O(N__30819),
            .I(un7_spon_5));
    LocalMux I__5239 (
            .O(N__30816),
            .I(un7_spon_5));
    InMux I__5238 (
            .O(N__30803),
            .I(N__30800));
    LocalMux I__5237 (
            .O(N__30800),
            .I(sEEPonPoff_i_5));
    InMux I__5236 (
            .O(N__30797),
            .I(N__30794));
    LocalMux I__5235 (
            .O(N__30794),
            .I(sEEPonPoffZ0Z_6));
    CascadeMux I__5234 (
            .O(N__30791),
            .I(N__30787));
    CascadeMux I__5233 (
            .O(N__30790),
            .I(N__30782));
    InMux I__5232 (
            .O(N__30787),
            .I(N__30778));
    CascadeMux I__5231 (
            .O(N__30786),
            .I(N__30775));
    CascadeMux I__5230 (
            .O(N__30785),
            .I(N__30770));
    InMux I__5229 (
            .O(N__30782),
            .I(N__30766));
    InMux I__5228 (
            .O(N__30781),
            .I(N__30763));
    LocalMux I__5227 (
            .O(N__30778),
            .I(N__30759));
    InMux I__5226 (
            .O(N__30775),
            .I(N__30756));
    CascadeMux I__5225 (
            .O(N__30774),
            .I(N__30753));
    InMux I__5224 (
            .O(N__30773),
            .I(N__30747));
    InMux I__5223 (
            .O(N__30770),
            .I(N__30747));
    InMux I__5222 (
            .O(N__30769),
            .I(N__30744));
    LocalMux I__5221 (
            .O(N__30766),
            .I(N__30739));
    LocalMux I__5220 (
            .O(N__30763),
            .I(N__30739));
    InMux I__5219 (
            .O(N__30762),
            .I(N__30736));
    Span4Mux_h I__5218 (
            .O(N__30759),
            .I(N__30731));
    LocalMux I__5217 (
            .O(N__30756),
            .I(N__30731));
    InMux I__5216 (
            .O(N__30753),
            .I(N__30728));
    InMux I__5215 (
            .O(N__30752),
            .I(N__30724));
    LocalMux I__5214 (
            .O(N__30747),
            .I(N__30719));
    LocalMux I__5213 (
            .O(N__30744),
            .I(N__30719));
    Span12Mux_v I__5212 (
            .O(N__30739),
            .I(N__30714));
    LocalMux I__5211 (
            .O(N__30736),
            .I(N__30714));
    Span4Mux_v I__5210 (
            .O(N__30731),
            .I(N__30711));
    LocalMux I__5209 (
            .O(N__30728),
            .I(N__30708));
    InMux I__5208 (
            .O(N__30727),
            .I(N__30705));
    LocalMux I__5207 (
            .O(N__30724),
            .I(un7_spon_6));
    Odrv4 I__5206 (
            .O(N__30719),
            .I(un7_spon_6));
    Odrv12 I__5205 (
            .O(N__30714),
            .I(un7_spon_6));
    Odrv4 I__5204 (
            .O(N__30711),
            .I(un7_spon_6));
    Odrv12 I__5203 (
            .O(N__30708),
            .I(un7_spon_6));
    LocalMux I__5202 (
            .O(N__30705),
            .I(un7_spon_6));
    InMux I__5201 (
            .O(N__30692),
            .I(N__30689));
    LocalMux I__5200 (
            .O(N__30689),
            .I(sEEPonPoff_i_6));
    CascadeMux I__5199 (
            .O(N__30686),
            .I(N__30683));
    InMux I__5198 (
            .O(N__30683),
            .I(N__30679));
    CascadeMux I__5197 (
            .O(N__30682),
            .I(N__30676));
    LocalMux I__5196 (
            .O(N__30679),
            .I(N__30671));
    InMux I__5195 (
            .O(N__30676),
            .I(N__30668));
    InMux I__5194 (
            .O(N__30675),
            .I(N__30664));
    InMux I__5193 (
            .O(N__30674),
            .I(N__30661));
    Span4Mux_h I__5192 (
            .O(N__30671),
            .I(N__30656));
    LocalMux I__5191 (
            .O(N__30668),
            .I(N__30656));
    InMux I__5190 (
            .O(N__30667),
            .I(N__30653));
    LocalMux I__5189 (
            .O(N__30664),
            .I(N__30644));
    LocalMux I__5188 (
            .O(N__30661),
            .I(N__30644));
    Span4Mux_h I__5187 (
            .O(N__30656),
            .I(N__30641));
    LocalMux I__5186 (
            .O(N__30653),
            .I(N__30638));
    InMux I__5185 (
            .O(N__30652),
            .I(N__30635));
    InMux I__5184 (
            .O(N__30651),
            .I(N__30631));
    InMux I__5183 (
            .O(N__30650),
            .I(N__30628));
    InMux I__5182 (
            .O(N__30649),
            .I(N__30624));
    Span4Mux_h I__5181 (
            .O(N__30644),
            .I(N__30621));
    Span4Mux_v I__5180 (
            .O(N__30641),
            .I(N__30616));
    Span4Mux_h I__5179 (
            .O(N__30638),
            .I(N__30616));
    LocalMux I__5178 (
            .O(N__30635),
            .I(N__30613));
    InMux I__5177 (
            .O(N__30634),
            .I(N__30610));
    LocalMux I__5176 (
            .O(N__30631),
            .I(N__30605));
    LocalMux I__5175 (
            .O(N__30628),
            .I(N__30605));
    InMux I__5174 (
            .O(N__30627),
            .I(N__30602));
    LocalMux I__5173 (
            .O(N__30624),
            .I(un7_spon_7));
    Odrv4 I__5172 (
            .O(N__30621),
            .I(un7_spon_7));
    Odrv4 I__5171 (
            .O(N__30616),
            .I(un7_spon_7));
    Odrv12 I__5170 (
            .O(N__30613),
            .I(un7_spon_7));
    LocalMux I__5169 (
            .O(N__30610),
            .I(un7_spon_7));
    Odrv12 I__5168 (
            .O(N__30605),
            .I(un7_spon_7));
    LocalMux I__5167 (
            .O(N__30602),
            .I(un7_spon_7));
    InMux I__5166 (
            .O(N__30587),
            .I(N__30584));
    LocalMux I__5165 (
            .O(N__30584),
            .I(sEEPonPoffZ0Z_7));
    InMux I__5164 (
            .O(N__30581),
            .I(N__30578));
    LocalMux I__5163 (
            .O(N__30578),
            .I(sEEPonPoff_i_7));
    CascadeMux I__5162 (
            .O(N__30575),
            .I(N__30572));
    InMux I__5161 (
            .O(N__30572),
            .I(N__30567));
    InMux I__5160 (
            .O(N__30571),
            .I(N__30564));
    CascadeMux I__5159 (
            .O(N__30570),
            .I(N__30559));
    LocalMux I__5158 (
            .O(N__30567),
            .I(N__30556));
    LocalMux I__5157 (
            .O(N__30564),
            .I(N__30552));
    InMux I__5156 (
            .O(N__30563),
            .I(N__30548));
    CascadeMux I__5155 (
            .O(N__30562),
            .I(N__30545));
    InMux I__5154 (
            .O(N__30559),
            .I(N__30542));
    Span4Mux_v I__5153 (
            .O(N__30556),
            .I(N__30538));
    InMux I__5152 (
            .O(N__30555),
            .I(N__30535));
    Span4Mux_v I__5151 (
            .O(N__30552),
            .I(N__30530));
    InMux I__5150 (
            .O(N__30551),
            .I(N__30527));
    LocalMux I__5149 (
            .O(N__30548),
            .I(N__30524));
    InMux I__5148 (
            .O(N__30545),
            .I(N__30521));
    LocalMux I__5147 (
            .O(N__30542),
            .I(N__30518));
    InMux I__5146 (
            .O(N__30541),
            .I(N__30514));
    Span4Mux_v I__5145 (
            .O(N__30538),
            .I(N__30509));
    LocalMux I__5144 (
            .O(N__30535),
            .I(N__30509));
    InMux I__5143 (
            .O(N__30534),
            .I(N__30504));
    InMux I__5142 (
            .O(N__30533),
            .I(N__30504));
    Span4Mux_v I__5141 (
            .O(N__30530),
            .I(N__30499));
    LocalMux I__5140 (
            .O(N__30527),
            .I(N__30499));
    Span4Mux_h I__5139 (
            .O(N__30524),
            .I(N__30496));
    LocalMux I__5138 (
            .O(N__30521),
            .I(N__30493));
    Span4Mux_h I__5137 (
            .O(N__30518),
            .I(N__30490));
    InMux I__5136 (
            .O(N__30517),
            .I(N__30487));
    LocalMux I__5135 (
            .O(N__30514),
            .I(un7_spon_8));
    Odrv4 I__5134 (
            .O(N__30509),
            .I(un7_spon_8));
    LocalMux I__5133 (
            .O(N__30504),
            .I(un7_spon_8));
    Odrv4 I__5132 (
            .O(N__30499),
            .I(un7_spon_8));
    Odrv4 I__5131 (
            .O(N__30496),
            .I(un7_spon_8));
    Odrv12 I__5130 (
            .O(N__30493),
            .I(un7_spon_8));
    Odrv4 I__5129 (
            .O(N__30490),
            .I(un7_spon_8));
    LocalMux I__5128 (
            .O(N__30487),
            .I(un7_spon_8));
    CascadeMux I__5127 (
            .O(N__30470),
            .I(N__30467));
    InMux I__5126 (
            .O(N__30467),
            .I(N__30462));
    InMux I__5125 (
            .O(N__30466),
            .I(N__30459));
    CascadeMux I__5124 (
            .O(N__30465),
            .I(N__30453));
    LocalMux I__5123 (
            .O(N__30462),
            .I(N__30450));
    LocalMux I__5122 (
            .O(N__30459),
            .I(N__30447));
    InMux I__5121 (
            .O(N__30458),
            .I(N__30442));
    InMux I__5120 (
            .O(N__30457),
            .I(N__30439));
    CascadeMux I__5119 (
            .O(N__30456),
            .I(N__30436));
    InMux I__5118 (
            .O(N__30453),
            .I(N__30433));
    Span4Mux_v I__5117 (
            .O(N__30450),
            .I(N__30430));
    Span4Mux_v I__5116 (
            .O(N__30447),
            .I(N__30427));
    CascadeMux I__5115 (
            .O(N__30446),
            .I(N__30423));
    InMux I__5114 (
            .O(N__30445),
            .I(N__30419));
    LocalMux I__5113 (
            .O(N__30442),
            .I(N__30414));
    LocalMux I__5112 (
            .O(N__30439),
            .I(N__30414));
    InMux I__5111 (
            .O(N__30436),
            .I(N__30411));
    LocalMux I__5110 (
            .O(N__30433),
            .I(N__30408));
    Span4Mux_v I__5109 (
            .O(N__30430),
            .I(N__30402));
    Span4Mux_v I__5108 (
            .O(N__30427),
            .I(N__30402));
    InMux I__5107 (
            .O(N__30426),
            .I(N__30399));
    InMux I__5106 (
            .O(N__30423),
            .I(N__30394));
    InMux I__5105 (
            .O(N__30422),
            .I(N__30394));
    LocalMux I__5104 (
            .O(N__30419),
            .I(N__30391));
    Span4Mux_h I__5103 (
            .O(N__30414),
            .I(N__30388));
    LocalMux I__5102 (
            .O(N__30411),
            .I(N__30385));
    Span4Mux_h I__5101 (
            .O(N__30408),
            .I(N__30382));
    InMux I__5100 (
            .O(N__30407),
            .I(N__30379));
    Odrv4 I__5099 (
            .O(N__30402),
            .I(un7_spon_9));
    LocalMux I__5098 (
            .O(N__30399),
            .I(un7_spon_9));
    LocalMux I__5097 (
            .O(N__30394),
            .I(un7_spon_9));
    Odrv4 I__5096 (
            .O(N__30391),
            .I(un7_spon_9));
    Odrv4 I__5095 (
            .O(N__30388),
            .I(un7_spon_9));
    Odrv12 I__5094 (
            .O(N__30385),
            .I(un7_spon_9));
    Odrv4 I__5093 (
            .O(N__30382),
            .I(un7_spon_9));
    LocalMux I__5092 (
            .O(N__30379),
            .I(un7_spon_9));
    CascadeMux I__5091 (
            .O(N__30362),
            .I(N__30357));
    CascadeMux I__5090 (
            .O(N__30361),
            .I(N__30354));
    InMux I__5089 (
            .O(N__30360),
            .I(N__30350));
    InMux I__5088 (
            .O(N__30357),
            .I(N__30347));
    InMux I__5087 (
            .O(N__30354),
            .I(N__30342));
    CascadeMux I__5086 (
            .O(N__30353),
            .I(N__30338));
    LocalMux I__5085 (
            .O(N__30350),
            .I(N__30334));
    LocalMux I__5084 (
            .O(N__30347),
            .I(N__30331));
    InMux I__5083 (
            .O(N__30346),
            .I(N__30328));
    InMux I__5082 (
            .O(N__30345),
            .I(N__30325));
    LocalMux I__5081 (
            .O(N__30342),
            .I(N__30322));
    CascadeMux I__5080 (
            .O(N__30341),
            .I(N__30319));
    InMux I__5079 (
            .O(N__30338),
            .I(N__30316));
    InMux I__5078 (
            .O(N__30337),
            .I(N__30311));
    Span4Mux_v I__5077 (
            .O(N__30334),
            .I(N__30308));
    Span4Mux_v I__5076 (
            .O(N__30331),
            .I(N__30303));
    LocalMux I__5075 (
            .O(N__30328),
            .I(N__30303));
    LocalMux I__5074 (
            .O(N__30325),
            .I(N__30300));
    Span4Mux_v I__5073 (
            .O(N__30322),
            .I(N__30297));
    InMux I__5072 (
            .O(N__30319),
            .I(N__30294));
    LocalMux I__5071 (
            .O(N__30316),
            .I(N__30291));
    InMux I__5070 (
            .O(N__30315),
            .I(N__30287));
    InMux I__5069 (
            .O(N__30314),
            .I(N__30284));
    LocalMux I__5068 (
            .O(N__30311),
            .I(N__30281));
    Span4Mux_v I__5067 (
            .O(N__30308),
            .I(N__30272));
    Span4Mux_v I__5066 (
            .O(N__30303),
            .I(N__30272));
    Span4Mux_h I__5065 (
            .O(N__30300),
            .I(N__30272));
    Span4Mux_h I__5064 (
            .O(N__30297),
            .I(N__30272));
    LocalMux I__5063 (
            .O(N__30294),
            .I(N__30269));
    Span4Mux_h I__5062 (
            .O(N__30291),
            .I(N__30266));
    InMux I__5061 (
            .O(N__30290),
            .I(N__30263));
    LocalMux I__5060 (
            .O(N__30287),
            .I(un7_spon_10));
    LocalMux I__5059 (
            .O(N__30284),
            .I(un7_spon_10));
    Odrv4 I__5058 (
            .O(N__30281),
            .I(un7_spon_10));
    Odrv4 I__5057 (
            .O(N__30272),
            .I(un7_spon_10));
    Odrv12 I__5056 (
            .O(N__30269),
            .I(un7_spon_10));
    Odrv4 I__5055 (
            .O(N__30266),
            .I(un7_spon_10));
    LocalMux I__5054 (
            .O(N__30263),
            .I(un7_spon_10));
    InMux I__5053 (
            .O(N__30248),
            .I(N__30245));
    LocalMux I__5052 (
            .O(N__30245),
            .I(sEEPonPoffZ0Z_0));
    CascadeMux I__5051 (
            .O(N__30242),
            .I(N__30238));
    InMux I__5050 (
            .O(N__30241),
            .I(N__30234));
    InMux I__5049 (
            .O(N__30238),
            .I(N__30230));
    CascadeMux I__5048 (
            .O(N__30237),
            .I(N__30226));
    LocalMux I__5047 (
            .O(N__30234),
            .I(N__30223));
    InMux I__5046 (
            .O(N__30233),
            .I(N__30220));
    LocalMux I__5045 (
            .O(N__30230),
            .I(N__30217));
    CascadeMux I__5044 (
            .O(N__30229),
            .I(N__30213));
    InMux I__5043 (
            .O(N__30226),
            .I(N__30210));
    Span4Mux_v I__5042 (
            .O(N__30223),
            .I(N__30207));
    LocalMux I__5041 (
            .O(N__30220),
            .I(N__30201));
    Span4Mux_v I__5040 (
            .O(N__30217),
            .I(N__30198));
    InMux I__5039 (
            .O(N__30216),
            .I(N__30195));
    InMux I__5038 (
            .O(N__30213),
            .I(N__30192));
    LocalMux I__5037 (
            .O(N__30210),
            .I(N__30189));
    Span4Mux_v I__5036 (
            .O(N__30207),
            .I(N__30185));
    InMux I__5035 (
            .O(N__30206),
            .I(N__30182));
    InMux I__5034 (
            .O(N__30205),
            .I(N__30177));
    InMux I__5033 (
            .O(N__30204),
            .I(N__30177));
    Span4Mux_h I__5032 (
            .O(N__30201),
            .I(N__30174));
    Span4Mux_v I__5031 (
            .O(N__30198),
            .I(N__30169));
    LocalMux I__5030 (
            .O(N__30195),
            .I(N__30169));
    LocalMux I__5029 (
            .O(N__30192),
            .I(N__30166));
    Span4Mux_h I__5028 (
            .O(N__30189),
            .I(N__30163));
    InMux I__5027 (
            .O(N__30188),
            .I(N__30160));
    Odrv4 I__5026 (
            .O(N__30185),
            .I(un7_spon_0));
    LocalMux I__5025 (
            .O(N__30182),
            .I(un7_spon_0));
    LocalMux I__5024 (
            .O(N__30177),
            .I(un7_spon_0));
    Odrv4 I__5023 (
            .O(N__30174),
            .I(un7_spon_0));
    Odrv4 I__5022 (
            .O(N__30169),
            .I(un7_spon_0));
    Odrv12 I__5021 (
            .O(N__30166),
            .I(un7_spon_0));
    Odrv4 I__5020 (
            .O(N__30163),
            .I(un7_spon_0));
    LocalMux I__5019 (
            .O(N__30160),
            .I(un7_spon_0));
    InMux I__5018 (
            .O(N__30143),
            .I(N__30140));
    LocalMux I__5017 (
            .O(N__30140),
            .I(sEEPonPoff_i_0));
    CascadeMux I__5016 (
            .O(N__30137),
            .I(N__30134));
    InMux I__5015 (
            .O(N__30134),
            .I(N__30131));
    LocalMux I__5014 (
            .O(N__30131),
            .I(N__30127));
    CascadeMux I__5013 (
            .O(N__30130),
            .I(N__30124));
    Span4Mux_v I__5012 (
            .O(N__30127),
            .I(N__30121));
    InMux I__5011 (
            .O(N__30124),
            .I(N__30118));
    Span4Mux_h I__5010 (
            .O(N__30121),
            .I(N__30112));
    LocalMux I__5009 (
            .O(N__30118),
            .I(N__30112));
    CascadeMux I__5008 (
            .O(N__30117),
            .I(N__30106));
    Span4Mux_v I__5007 (
            .O(N__30112),
            .I(N__30103));
    InMux I__5006 (
            .O(N__30111),
            .I(N__30100));
    InMux I__5005 (
            .O(N__30110),
            .I(N__30097));
    CascadeMux I__5004 (
            .O(N__30109),
            .I(N__30093));
    InMux I__5003 (
            .O(N__30106),
            .I(N__30090));
    Span4Mux_h I__5002 (
            .O(N__30103),
            .I(N__30082));
    LocalMux I__5001 (
            .O(N__30100),
            .I(N__30082));
    LocalMux I__5000 (
            .O(N__30097),
            .I(N__30082));
    InMux I__4999 (
            .O(N__30096),
            .I(N__30077));
    InMux I__4998 (
            .O(N__30093),
            .I(N__30074));
    LocalMux I__4997 (
            .O(N__30090),
            .I(N__30071));
    InMux I__4996 (
            .O(N__30089),
            .I(N__30067));
    Span4Mux_v I__4995 (
            .O(N__30082),
            .I(N__30064));
    InMux I__4994 (
            .O(N__30081),
            .I(N__30059));
    InMux I__4993 (
            .O(N__30080),
            .I(N__30059));
    LocalMux I__4992 (
            .O(N__30077),
            .I(N__30056));
    LocalMux I__4991 (
            .O(N__30074),
            .I(N__30053));
    Span4Mux_h I__4990 (
            .O(N__30071),
            .I(N__30050));
    InMux I__4989 (
            .O(N__30070),
            .I(N__30047));
    LocalMux I__4988 (
            .O(N__30067),
            .I(un7_spon_1));
    Odrv4 I__4987 (
            .O(N__30064),
            .I(un7_spon_1));
    LocalMux I__4986 (
            .O(N__30059),
            .I(un7_spon_1));
    Odrv12 I__4985 (
            .O(N__30056),
            .I(un7_spon_1));
    Odrv12 I__4984 (
            .O(N__30053),
            .I(un7_spon_1));
    Odrv4 I__4983 (
            .O(N__30050),
            .I(un7_spon_1));
    LocalMux I__4982 (
            .O(N__30047),
            .I(un7_spon_1));
    InMux I__4981 (
            .O(N__30032),
            .I(N__30029));
    LocalMux I__4980 (
            .O(N__30029),
            .I(sEEPonPoffZ0Z_1));
    InMux I__4979 (
            .O(N__30026),
            .I(N__30023));
    LocalMux I__4978 (
            .O(N__30023),
            .I(sEEPonPoff_i_1));
    InMux I__4977 (
            .O(N__30020),
            .I(N__30017));
    LocalMux I__4976 (
            .O(N__30017),
            .I(sEEPonPoffZ0Z_2));
    CascadeMux I__4975 (
            .O(N__30014),
            .I(N__30010));
    CascadeMux I__4974 (
            .O(N__30013),
            .I(N__30007));
    InMux I__4973 (
            .O(N__30010),
            .I(N__30002));
    InMux I__4972 (
            .O(N__30007),
            .I(N__29999));
    CascadeMux I__4971 (
            .O(N__30006),
            .I(N__29993));
    InMux I__4970 (
            .O(N__30005),
            .I(N__29990));
    LocalMux I__4969 (
            .O(N__30002),
            .I(N__29987));
    LocalMux I__4968 (
            .O(N__29999),
            .I(N__29984));
    InMux I__4967 (
            .O(N__29998),
            .I(N__29980));
    CascadeMux I__4966 (
            .O(N__29997),
            .I(N__29977));
    CascadeMux I__4965 (
            .O(N__29996),
            .I(N__29974));
    InMux I__4964 (
            .O(N__29993),
            .I(N__29971));
    LocalMux I__4963 (
            .O(N__29990),
            .I(N__29966));
    Span4Mux_h I__4962 (
            .O(N__29987),
            .I(N__29961));
    Span4Mux_h I__4961 (
            .O(N__29984),
            .I(N__29961));
    InMux I__4960 (
            .O(N__29983),
            .I(N__29958));
    LocalMux I__4959 (
            .O(N__29980),
            .I(N__29955));
    InMux I__4958 (
            .O(N__29977),
            .I(N__29952));
    InMux I__4957 (
            .O(N__29974),
            .I(N__29949));
    LocalMux I__4956 (
            .O(N__29971),
            .I(N__29946));
    InMux I__4955 (
            .O(N__29970),
            .I(N__29942));
    InMux I__4954 (
            .O(N__29969),
            .I(N__29939));
    Span4Mux_v I__4953 (
            .O(N__29966),
            .I(N__29936));
    Span4Mux_v I__4952 (
            .O(N__29961),
            .I(N__29931));
    LocalMux I__4951 (
            .O(N__29958),
            .I(N__29931));
    Span4Mux_h I__4950 (
            .O(N__29955),
            .I(N__29928));
    LocalMux I__4949 (
            .O(N__29952),
            .I(N__29925));
    LocalMux I__4948 (
            .O(N__29949),
            .I(N__29922));
    Span4Mux_h I__4947 (
            .O(N__29946),
            .I(N__29919));
    InMux I__4946 (
            .O(N__29945),
            .I(N__29916));
    LocalMux I__4945 (
            .O(N__29942),
            .I(un7_spon_2));
    LocalMux I__4944 (
            .O(N__29939),
            .I(un7_spon_2));
    Odrv4 I__4943 (
            .O(N__29936),
            .I(un7_spon_2));
    Odrv4 I__4942 (
            .O(N__29931),
            .I(un7_spon_2));
    Odrv4 I__4941 (
            .O(N__29928),
            .I(un7_spon_2));
    Odrv12 I__4940 (
            .O(N__29925),
            .I(un7_spon_2));
    Odrv12 I__4939 (
            .O(N__29922),
            .I(un7_spon_2));
    Odrv4 I__4938 (
            .O(N__29919),
            .I(un7_spon_2));
    LocalMux I__4937 (
            .O(N__29916),
            .I(un7_spon_2));
    InMux I__4936 (
            .O(N__29897),
            .I(N__29894));
    LocalMux I__4935 (
            .O(N__29894),
            .I(sEEPonPoff_i_2));
    InMux I__4934 (
            .O(N__29891),
            .I(N__29888));
    LocalMux I__4933 (
            .O(N__29888),
            .I(sEEPonPoffZ0Z_3));
    CascadeMux I__4932 (
            .O(N__29885),
            .I(N__29881));
    CascadeMux I__4931 (
            .O(N__29884),
            .I(N__29878));
    InMux I__4930 (
            .O(N__29881),
            .I(N__29874));
    InMux I__4929 (
            .O(N__29878),
            .I(N__29868));
    CascadeMux I__4928 (
            .O(N__29877),
            .I(N__29864));
    LocalMux I__4927 (
            .O(N__29874),
            .I(N__29861));
    InMux I__4926 (
            .O(N__29873),
            .I(N__29858));
    InMux I__4925 (
            .O(N__29872),
            .I(N__29855));
    InMux I__4924 (
            .O(N__29871),
            .I(N__29852));
    LocalMux I__4923 (
            .O(N__29868),
            .I(N__29848));
    InMux I__4922 (
            .O(N__29867),
            .I(N__29845));
    InMux I__4921 (
            .O(N__29864),
            .I(N__29842));
    Span4Mux_v I__4920 (
            .O(N__29861),
            .I(N__29833));
    LocalMux I__4919 (
            .O(N__29858),
            .I(N__29833));
    LocalMux I__4918 (
            .O(N__29855),
            .I(N__29833));
    LocalMux I__4917 (
            .O(N__29852),
            .I(N__29830));
    InMux I__4916 (
            .O(N__29851),
            .I(N__29827));
    Span4Mux_h I__4915 (
            .O(N__29848),
            .I(N__29822));
    LocalMux I__4914 (
            .O(N__29845),
            .I(N__29822));
    LocalMux I__4913 (
            .O(N__29842),
            .I(N__29819));
    InMux I__4912 (
            .O(N__29841),
            .I(N__29815));
    InMux I__4911 (
            .O(N__29840),
            .I(N__29812));
    Span4Mux_v I__4910 (
            .O(N__29833),
            .I(N__29807));
    Span4Mux_h I__4909 (
            .O(N__29830),
            .I(N__29807));
    LocalMux I__4908 (
            .O(N__29827),
            .I(N__29802));
    Span4Mux_v I__4907 (
            .O(N__29822),
            .I(N__29802));
    Span4Mux_h I__4906 (
            .O(N__29819),
            .I(N__29799));
    InMux I__4905 (
            .O(N__29818),
            .I(N__29796));
    LocalMux I__4904 (
            .O(N__29815),
            .I(un7_spon_3));
    LocalMux I__4903 (
            .O(N__29812),
            .I(un7_spon_3));
    Odrv4 I__4902 (
            .O(N__29807),
            .I(un7_spon_3));
    Odrv4 I__4901 (
            .O(N__29802),
            .I(un7_spon_3));
    Odrv4 I__4900 (
            .O(N__29799),
            .I(un7_spon_3));
    LocalMux I__4899 (
            .O(N__29796),
            .I(un7_spon_3));
    InMux I__4898 (
            .O(N__29783),
            .I(N__29780));
    LocalMux I__4897 (
            .O(N__29780),
            .I(sEEPonPoff_i_3));
    InMux I__4896 (
            .O(N__29777),
            .I(N__29774));
    LocalMux I__4895 (
            .O(N__29774),
            .I(N__29771));
    Odrv4 I__4894 (
            .O(N__29771),
            .I(sDAC_mem_27Z0Z_2));
    InMux I__4893 (
            .O(N__29768),
            .I(N__29765));
    LocalMux I__4892 (
            .O(N__29765),
            .I(N__29762));
    Span4Mux_h I__4891 (
            .O(N__29762),
            .I(N__29759));
    Odrv4 I__4890 (
            .O(N__29759),
            .I(sDAC_mem_27Z0Z_4));
    InMux I__4889 (
            .O(N__29756),
            .I(N__29753));
    LocalMux I__4888 (
            .O(N__29753),
            .I(N__29750));
    Odrv4 I__4887 (
            .O(N__29750),
            .I(sDAC_mem_27Z0Z_5));
    InMux I__4886 (
            .O(N__29747),
            .I(N__29744));
    LocalMux I__4885 (
            .O(N__29744),
            .I(N__29741));
    Span4Mux_v I__4884 (
            .O(N__29741),
            .I(N__29738));
    Odrv4 I__4883 (
            .O(N__29738),
            .I(sDAC_mem_27Z0Z_6));
    InMux I__4882 (
            .O(N__29735),
            .I(N__29732));
    LocalMux I__4881 (
            .O(N__29732),
            .I(N__29729));
    Odrv4 I__4880 (
            .O(N__29729),
            .I(sDAC_mem_27Z0Z_7));
    CEMux I__4879 (
            .O(N__29726),
            .I(N__29723));
    LocalMux I__4878 (
            .O(N__29723),
            .I(N__29720));
    Span12Mux_h I__4877 (
            .O(N__29720),
            .I(N__29717));
    Odrv12 I__4876 (
            .O(N__29717),
            .I(sDAC_mem_27_1_sqmuxa));
    InMux I__4875 (
            .O(N__29714),
            .I(N__29711));
    LocalMux I__4874 (
            .O(N__29711),
            .I(sDAC_mem_28Z0Z_6));
    InMux I__4873 (
            .O(N__29708),
            .I(N__29705));
    LocalMux I__4872 (
            .O(N__29705),
            .I(N__29702));
    Odrv12 I__4871 (
            .O(N__29702),
            .I(sDAC_mem_31Z0Z_0));
    InMux I__4870 (
            .O(N__29699),
            .I(N__29696));
    LocalMux I__4869 (
            .O(N__29696),
            .I(N__29693));
    Span4Mux_v I__4868 (
            .O(N__29693),
            .I(N__29690));
    Span4Mux_h I__4867 (
            .O(N__29690),
            .I(N__29687));
    Odrv4 I__4866 (
            .O(N__29687),
            .I(sDAC_mem_30Z0Z_0));
    InMux I__4865 (
            .O(N__29684),
            .I(N__29681));
    LocalMux I__4864 (
            .O(N__29681),
            .I(N__29678));
    Odrv12 I__4863 (
            .O(N__29678),
            .I(sDAC_mem_31Z0Z_3));
    InMux I__4862 (
            .O(N__29675),
            .I(N__29672));
    LocalMux I__4861 (
            .O(N__29672),
            .I(N__29669));
    Span12Mux_h I__4860 (
            .O(N__29669),
            .I(N__29666));
    Odrv12 I__4859 (
            .O(N__29666),
            .I(sDAC_mem_30Z0Z_3));
    InMux I__4858 (
            .O(N__29663),
            .I(N__29660));
    LocalMux I__4857 (
            .O(N__29660),
            .I(N__29657));
    Span4Mux_h I__4856 (
            .O(N__29657),
            .I(N__29654));
    Odrv4 I__4855 (
            .O(N__29654),
            .I(sDAC_mem_31Z0Z_6));
    InMux I__4854 (
            .O(N__29651),
            .I(N__29648));
    LocalMux I__4853 (
            .O(N__29648),
            .I(N__29645));
    Span4Mux_h I__4852 (
            .O(N__29645),
            .I(N__29642));
    Span4Mux_h I__4851 (
            .O(N__29642),
            .I(N__29639));
    Odrv4 I__4850 (
            .O(N__29639),
            .I(sDAC_mem_30Z0Z_6));
    InMux I__4849 (
            .O(N__29636),
            .I(N__29633));
    LocalMux I__4848 (
            .O(N__29633),
            .I(N__29630));
    Span4Mux_v I__4847 (
            .O(N__29630),
            .I(N__29627));
    Odrv4 I__4846 (
            .O(N__29627),
            .I(sDAC_data_RNO_24Z0Z_9));
    InMux I__4845 (
            .O(N__29624),
            .I(N__29621));
    LocalMux I__4844 (
            .O(N__29621),
            .I(N__29618));
    Span4Mux_h I__4843 (
            .O(N__29618),
            .I(N__29615));
    Span4Mux_h I__4842 (
            .O(N__29615),
            .I(N__29612));
    Odrv4 I__4841 (
            .O(N__29612),
            .I(sDAC_mem_16Z0Z_0));
    InMux I__4840 (
            .O(N__29609),
            .I(N__29606));
    LocalMux I__4839 (
            .O(N__29606),
            .I(N__29603));
    Span4Mux_h I__4838 (
            .O(N__29603),
            .I(N__29600));
    Span4Mux_h I__4837 (
            .O(N__29600),
            .I(N__29597));
    Odrv4 I__4836 (
            .O(N__29597),
            .I(sDAC_mem_16Z0Z_1));
    InMux I__4835 (
            .O(N__29594),
            .I(N__29591));
    LocalMux I__4834 (
            .O(N__29591),
            .I(N__29588));
    Span4Mux_v I__4833 (
            .O(N__29588),
            .I(N__29585));
    Odrv4 I__4832 (
            .O(N__29585),
            .I(sDAC_data_RNO_28Z0Z_4));
    InMux I__4831 (
            .O(N__29582),
            .I(N__29579));
    LocalMux I__4830 (
            .O(N__29579),
            .I(N__29576));
    Span12Mux_h I__4829 (
            .O(N__29576),
            .I(N__29573));
    Odrv12 I__4828 (
            .O(N__29573),
            .I(sDAC_mem_16Z0Z_2));
    InMux I__4827 (
            .O(N__29570),
            .I(N__29567));
    LocalMux I__4826 (
            .O(N__29567),
            .I(N__29564));
    Odrv4 I__4825 (
            .O(N__29564),
            .I(sDAC_mem_27Z0Z_1));
    InMux I__4824 (
            .O(N__29561),
            .I(N__29558));
    LocalMux I__4823 (
            .O(N__29558),
            .I(N__29551));
    InMux I__4822 (
            .O(N__29557),
            .I(N__29548));
    InMux I__4821 (
            .O(N__29556),
            .I(N__29545));
    InMux I__4820 (
            .O(N__29555),
            .I(N__29540));
    InMux I__4819 (
            .O(N__29554),
            .I(N__29540));
    Span12Mux_v I__4818 (
            .O(N__29551),
            .I(N__29535));
    LocalMux I__4817 (
            .O(N__29548),
            .I(N__29535));
    LocalMux I__4816 (
            .O(N__29545),
            .I(N_106));
    LocalMux I__4815 (
            .O(N__29540),
            .I(N_106));
    Odrv12 I__4814 (
            .O(N__29535),
            .I(N_106));
    InMux I__4813 (
            .O(N__29528),
            .I(bfn_14_13_0_));
    InMux I__4812 (
            .O(N__29525),
            .I(N__29522));
    LocalMux I__4811 (
            .O(N__29522),
            .I(N__29519));
    Span4Mux_h I__4810 (
            .O(N__29519),
            .I(N__29516));
    Odrv4 I__4809 (
            .O(N__29516),
            .I(sDAC_mem_24Z0Z_7));
    InMux I__4808 (
            .O(N__29513),
            .I(N__29510));
    LocalMux I__4807 (
            .O(N__29510),
            .I(N__29507));
    Span4Mux_h I__4806 (
            .O(N__29507),
            .I(N__29504));
    Span4Mux_h I__4805 (
            .O(N__29504),
            .I(N__29501));
    Odrv4 I__4804 (
            .O(N__29501),
            .I(sDAC_mem_26Z0Z_7));
    InMux I__4803 (
            .O(N__29498),
            .I(N__29495));
    LocalMux I__4802 (
            .O(N__29495),
            .I(N__29492));
    Span4Mux_v I__4801 (
            .O(N__29492),
            .I(N__29489));
    Span4Mux_h I__4800 (
            .O(N__29489),
            .I(N__29486));
    Span4Mux_v I__4799 (
            .O(N__29486),
            .I(N__29483));
    Odrv4 I__4798 (
            .O(N__29483),
            .I(sDAC_dataZ0Z_10));
    InMux I__4797 (
            .O(N__29480),
            .I(N__29477));
    LocalMux I__4796 (
            .O(N__29477),
            .I(N__29474));
    Span4Mux_h I__4795 (
            .O(N__29474),
            .I(N__29471));
    Odrv4 I__4794 (
            .O(N__29471),
            .I(sDAC_mem_24Z0Z_2));
    InMux I__4793 (
            .O(N__29468),
            .I(N__29465));
    LocalMux I__4792 (
            .O(N__29465),
            .I(sDAC_data_RNO_30Z0Z_5));
    InMux I__4791 (
            .O(N__29462),
            .I(N__29459));
    LocalMux I__4790 (
            .O(N__29459),
            .I(N__29456));
    Span4Mux_v I__4789 (
            .O(N__29456),
            .I(N__29453));
    Odrv4 I__4788 (
            .O(N__29453),
            .I(sDAC_mem_24Z0Z_5));
    InMux I__4787 (
            .O(N__29450),
            .I(N__29447));
    LocalMux I__4786 (
            .O(N__29447),
            .I(N__29444));
    Span4Mux_h I__4785 (
            .O(N__29444),
            .I(N__29441));
    Odrv4 I__4784 (
            .O(N__29441),
            .I(sDAC_data_RNO_30Z0Z_8));
    InMux I__4783 (
            .O(N__29438),
            .I(N__29435));
    LocalMux I__4782 (
            .O(N__29435),
            .I(N__29432));
    Span4Mux_h I__4781 (
            .O(N__29432),
            .I(N__29429));
    Span4Mux_h I__4780 (
            .O(N__29429),
            .I(N__29426));
    Odrv4 I__4779 (
            .O(N__29426),
            .I(sDAC_mem_29Z0Z_6));
    InMux I__4778 (
            .O(N__29423),
            .I(N__29420));
    LocalMux I__4777 (
            .O(N__29420),
            .I(N__29417));
    Span4Mux_v I__4776 (
            .O(N__29417),
            .I(N__29414));
    Odrv4 I__4775 (
            .O(N__29414),
            .I(sDAC_data_RNO_23Z0Z_9));
    InMux I__4774 (
            .O(N__29411),
            .I(N__29408));
    LocalMux I__4773 (
            .O(N__29408),
            .I(N__29404));
    CascadeMux I__4772 (
            .O(N__29407),
            .I(N__29401));
    Span4Mux_h I__4771 (
            .O(N__29404),
            .I(N__29398));
    InMux I__4770 (
            .O(N__29401),
            .I(N__29395));
    Odrv4 I__4769 (
            .O(N__29398),
            .I(sEEACQZ0Z_15));
    LocalMux I__4768 (
            .O(N__29395),
            .I(sEEACQZ0Z_15));
    CascadeMux I__4767 (
            .O(N__29390),
            .I(N__29387));
    InMux I__4766 (
            .O(N__29387),
            .I(N__29384));
    LocalMux I__4765 (
            .O(N__29384),
            .I(N__29381));
    Odrv4 I__4764 (
            .O(N__29381),
            .I(sEEACQ_i_15));
    InMux I__4763 (
            .O(N__29378),
            .I(N__29374));
    CascadeMux I__4762 (
            .O(N__29377),
            .I(N__29371));
    LocalMux I__4761 (
            .O(N__29374),
            .I(N__29368));
    InMux I__4760 (
            .O(N__29371),
            .I(N__29365));
    Span4Mux_h I__4759 (
            .O(N__29368),
            .I(N__29362));
    LocalMux I__4758 (
            .O(N__29365),
            .I(N__29357));
    Span4Mux_v I__4757 (
            .O(N__29362),
            .I(N__29357));
    Odrv4 I__4756 (
            .O(N__29357),
            .I(sEEACQZ0Z_7));
    CascadeMux I__4755 (
            .O(N__29354),
            .I(N__29351));
    InMux I__4754 (
            .O(N__29351),
            .I(N__29348));
    LocalMux I__4753 (
            .O(N__29348),
            .I(sEEACQ_i_7));
    InMux I__4752 (
            .O(N__29345),
            .I(N__29342));
    LocalMux I__4751 (
            .O(N__29342),
            .I(N__29338));
    CascadeMux I__4750 (
            .O(N__29341),
            .I(N__29335));
    Span12Mux_v I__4749 (
            .O(N__29338),
            .I(N__29332));
    InMux I__4748 (
            .O(N__29335),
            .I(N__29329));
    Odrv12 I__4747 (
            .O(N__29332),
            .I(sEEACQZ0Z_8));
    LocalMux I__4746 (
            .O(N__29329),
            .I(sEEACQZ0Z_8));
    CascadeMux I__4745 (
            .O(N__29324),
            .I(N__29321));
    InMux I__4744 (
            .O(N__29321),
            .I(N__29318));
    LocalMux I__4743 (
            .O(N__29318),
            .I(sEEACQ_i_8));
    InMux I__4742 (
            .O(N__29315),
            .I(N__29312));
    LocalMux I__4741 (
            .O(N__29312),
            .I(N__29309));
    Span4Mux_h I__4740 (
            .O(N__29309),
            .I(N__29305));
    CascadeMux I__4739 (
            .O(N__29308),
            .I(N__29302));
    Span4Mux_v I__4738 (
            .O(N__29305),
            .I(N__29299));
    InMux I__4737 (
            .O(N__29302),
            .I(N__29296));
    Odrv4 I__4736 (
            .O(N__29299),
            .I(sEEACQZ0Z_9));
    LocalMux I__4735 (
            .O(N__29296),
            .I(sEEACQZ0Z_9));
    CascadeMux I__4734 (
            .O(N__29291),
            .I(N__29288));
    InMux I__4733 (
            .O(N__29288),
            .I(N__29285));
    LocalMux I__4732 (
            .O(N__29285),
            .I(sEEACQ_i_9));
    InMux I__4731 (
            .O(N__29282),
            .I(N__29279));
    LocalMux I__4730 (
            .O(N__29279),
            .I(N__29275));
    CascadeMux I__4729 (
            .O(N__29278),
            .I(N__29272));
    Span4Mux_h I__4728 (
            .O(N__29275),
            .I(N__29269));
    InMux I__4727 (
            .O(N__29272),
            .I(N__29266));
    Span4Mux_v I__4726 (
            .O(N__29269),
            .I(N__29261));
    LocalMux I__4725 (
            .O(N__29266),
            .I(N__29261));
    Odrv4 I__4724 (
            .O(N__29261),
            .I(sEEACQZ0Z_10));
    CascadeMux I__4723 (
            .O(N__29258),
            .I(N__29255));
    InMux I__4722 (
            .O(N__29255),
            .I(N__29252));
    LocalMux I__4721 (
            .O(N__29252),
            .I(sEEACQ_i_10));
    InMux I__4720 (
            .O(N__29249),
            .I(N__29245));
    CascadeMux I__4719 (
            .O(N__29248),
            .I(N__29242));
    LocalMux I__4718 (
            .O(N__29245),
            .I(N__29239));
    InMux I__4717 (
            .O(N__29242),
            .I(N__29236));
    Span4Mux_h I__4716 (
            .O(N__29239),
            .I(N__29233));
    LocalMux I__4715 (
            .O(N__29236),
            .I(N__29230));
    Odrv4 I__4714 (
            .O(N__29233),
            .I(sEEACQZ0Z_11));
    Odrv4 I__4713 (
            .O(N__29230),
            .I(sEEACQZ0Z_11));
    CascadeMux I__4712 (
            .O(N__29225),
            .I(N__29222));
    InMux I__4711 (
            .O(N__29222),
            .I(N__29219));
    LocalMux I__4710 (
            .O(N__29219),
            .I(sEEACQ_i_11));
    InMux I__4709 (
            .O(N__29216),
            .I(N__29213));
    LocalMux I__4708 (
            .O(N__29213),
            .I(N__29209));
    CascadeMux I__4707 (
            .O(N__29212),
            .I(N__29206));
    Span4Mux_h I__4706 (
            .O(N__29209),
            .I(N__29203));
    InMux I__4705 (
            .O(N__29206),
            .I(N__29200));
    Odrv4 I__4704 (
            .O(N__29203),
            .I(sEEACQZ0Z_12));
    LocalMux I__4703 (
            .O(N__29200),
            .I(sEEACQZ0Z_12));
    CascadeMux I__4702 (
            .O(N__29195),
            .I(N__29192));
    InMux I__4701 (
            .O(N__29192),
            .I(N__29189));
    LocalMux I__4700 (
            .O(N__29189),
            .I(sEEACQ_i_12));
    InMux I__4699 (
            .O(N__29186),
            .I(N__29183));
    LocalMux I__4698 (
            .O(N__29183),
            .I(N__29179));
    CascadeMux I__4697 (
            .O(N__29182),
            .I(N__29176));
    Span4Mux_h I__4696 (
            .O(N__29179),
            .I(N__29173));
    InMux I__4695 (
            .O(N__29176),
            .I(N__29170));
    Odrv4 I__4694 (
            .O(N__29173),
            .I(sEEACQZ0Z_13));
    LocalMux I__4693 (
            .O(N__29170),
            .I(sEEACQZ0Z_13));
    CascadeMux I__4692 (
            .O(N__29165),
            .I(N__29162));
    InMux I__4691 (
            .O(N__29162),
            .I(N__29159));
    LocalMux I__4690 (
            .O(N__29159),
            .I(sEEACQ_i_13));
    InMux I__4689 (
            .O(N__29156),
            .I(N__29152));
    CascadeMux I__4688 (
            .O(N__29155),
            .I(N__29149));
    LocalMux I__4687 (
            .O(N__29152),
            .I(N__29146));
    InMux I__4686 (
            .O(N__29149),
            .I(N__29143));
    Span4Mux_h I__4685 (
            .O(N__29146),
            .I(N__29140));
    LocalMux I__4684 (
            .O(N__29143),
            .I(N__29137));
    Odrv4 I__4683 (
            .O(N__29140),
            .I(sEEACQZ0Z_14));
    Odrv4 I__4682 (
            .O(N__29137),
            .I(sEEACQZ0Z_14));
    InMux I__4681 (
            .O(N__29132),
            .I(N__29129));
    LocalMux I__4680 (
            .O(N__29129),
            .I(sEEACQ_i_14));
    InMux I__4679 (
            .O(N__29126),
            .I(N__29123));
    LocalMux I__4678 (
            .O(N__29123),
            .I(sDAC_mem_12Z0Z_3));
    InMux I__4677 (
            .O(N__29120),
            .I(N__29116));
    CascadeMux I__4676 (
            .O(N__29119),
            .I(N__29113));
    LocalMux I__4675 (
            .O(N__29116),
            .I(N__29110));
    InMux I__4674 (
            .O(N__29113),
            .I(N__29107));
    Span4Mux_h I__4673 (
            .O(N__29110),
            .I(N__29104));
    LocalMux I__4672 (
            .O(N__29107),
            .I(N__29101));
    Odrv4 I__4671 (
            .O(N__29104),
            .I(sEEACQZ0Z_0));
    Odrv4 I__4670 (
            .O(N__29101),
            .I(sEEACQZ0Z_0));
    CascadeMux I__4669 (
            .O(N__29096),
            .I(N__29093));
    InMux I__4668 (
            .O(N__29093),
            .I(N__29090));
    LocalMux I__4667 (
            .O(N__29090),
            .I(sEEACQ_i_0));
    InMux I__4666 (
            .O(N__29087),
            .I(N__29083));
    CascadeMux I__4665 (
            .O(N__29086),
            .I(N__29080));
    LocalMux I__4664 (
            .O(N__29083),
            .I(N__29077));
    InMux I__4663 (
            .O(N__29080),
            .I(N__29074));
    Span4Mux_h I__4662 (
            .O(N__29077),
            .I(N__29071));
    LocalMux I__4661 (
            .O(N__29074),
            .I(N__29068));
    Odrv4 I__4660 (
            .O(N__29071),
            .I(sEEACQZ0Z_1));
    Odrv4 I__4659 (
            .O(N__29068),
            .I(sEEACQZ0Z_1));
    CascadeMux I__4658 (
            .O(N__29063),
            .I(N__29060));
    InMux I__4657 (
            .O(N__29060),
            .I(N__29057));
    LocalMux I__4656 (
            .O(N__29057),
            .I(sEEACQ_i_1));
    InMux I__4655 (
            .O(N__29054),
            .I(N__29051));
    LocalMux I__4654 (
            .O(N__29051),
            .I(N__29047));
    CascadeMux I__4653 (
            .O(N__29050),
            .I(N__29044));
    Span4Mux_h I__4652 (
            .O(N__29047),
            .I(N__29041));
    InMux I__4651 (
            .O(N__29044),
            .I(N__29038));
    Odrv4 I__4650 (
            .O(N__29041),
            .I(sEEACQZ0Z_2));
    LocalMux I__4649 (
            .O(N__29038),
            .I(sEEACQZ0Z_2));
    InMux I__4648 (
            .O(N__29033),
            .I(N__29030));
    LocalMux I__4647 (
            .O(N__29030),
            .I(sEEACQ_i_2));
    InMux I__4646 (
            .O(N__29027),
            .I(N__29024));
    LocalMux I__4645 (
            .O(N__29024),
            .I(N__29020));
    CascadeMux I__4644 (
            .O(N__29023),
            .I(N__29017));
    Span4Mux_h I__4643 (
            .O(N__29020),
            .I(N__29014));
    InMux I__4642 (
            .O(N__29017),
            .I(N__29011));
    Odrv4 I__4641 (
            .O(N__29014),
            .I(sEEACQZ0Z_3));
    LocalMux I__4640 (
            .O(N__29011),
            .I(sEEACQZ0Z_3));
    CascadeMux I__4639 (
            .O(N__29006),
            .I(N__29003));
    InMux I__4638 (
            .O(N__29003),
            .I(N__29000));
    LocalMux I__4637 (
            .O(N__29000),
            .I(sEEACQ_i_3));
    InMux I__4636 (
            .O(N__28997),
            .I(N__28993));
    CascadeMux I__4635 (
            .O(N__28996),
            .I(N__28990));
    LocalMux I__4634 (
            .O(N__28993),
            .I(N__28987));
    InMux I__4633 (
            .O(N__28990),
            .I(N__28984));
    Span4Mux_h I__4632 (
            .O(N__28987),
            .I(N__28981));
    LocalMux I__4631 (
            .O(N__28984),
            .I(N__28978));
    Odrv4 I__4630 (
            .O(N__28981),
            .I(sEEACQZ0Z_4));
    Odrv4 I__4629 (
            .O(N__28978),
            .I(sEEACQZ0Z_4));
    CascadeMux I__4628 (
            .O(N__28973),
            .I(N__28970));
    InMux I__4627 (
            .O(N__28970),
            .I(N__28967));
    LocalMux I__4626 (
            .O(N__28967),
            .I(sEEACQ_i_4));
    InMux I__4625 (
            .O(N__28964),
            .I(N__28961));
    LocalMux I__4624 (
            .O(N__28961),
            .I(N__28957));
    CascadeMux I__4623 (
            .O(N__28960),
            .I(N__28954));
    Span4Mux_h I__4622 (
            .O(N__28957),
            .I(N__28951));
    InMux I__4621 (
            .O(N__28954),
            .I(N__28948));
    Odrv4 I__4620 (
            .O(N__28951),
            .I(sEEACQZ0Z_5));
    LocalMux I__4619 (
            .O(N__28948),
            .I(sEEACQZ0Z_5));
    CascadeMux I__4618 (
            .O(N__28943),
            .I(N__28940));
    InMux I__4617 (
            .O(N__28940),
            .I(N__28937));
    LocalMux I__4616 (
            .O(N__28937),
            .I(sEEACQ_i_5));
    InMux I__4615 (
            .O(N__28934),
            .I(N__28931));
    LocalMux I__4614 (
            .O(N__28931),
            .I(N__28927));
    CascadeMux I__4613 (
            .O(N__28930),
            .I(N__28924));
    Span12Mux_v I__4612 (
            .O(N__28927),
            .I(N__28921));
    InMux I__4611 (
            .O(N__28924),
            .I(N__28918));
    Odrv12 I__4610 (
            .O(N__28921),
            .I(sEEACQZ0Z_6));
    LocalMux I__4609 (
            .O(N__28918),
            .I(sEEACQZ0Z_6));
    CascadeMux I__4608 (
            .O(N__28913),
            .I(N__28910));
    InMux I__4607 (
            .O(N__28910),
            .I(N__28907));
    LocalMux I__4606 (
            .O(N__28907),
            .I(sEEACQ_i_6));
    InMux I__4605 (
            .O(N__28904),
            .I(N__28901));
    LocalMux I__4604 (
            .O(N__28901),
            .I(sDAC_data_2_14_ns_1_4));
    InMux I__4603 (
            .O(N__28898),
            .I(N__28895));
    LocalMux I__4602 (
            .O(N__28895),
            .I(sDAC_data_2_32_ns_1_4));
    InMux I__4601 (
            .O(N__28892),
            .I(N__28889));
    LocalMux I__4600 (
            .O(N__28889),
            .I(N__28886));
    Odrv12 I__4599 (
            .O(N__28886),
            .I(sDAC_mem_15Z0Z_2));
    InMux I__4598 (
            .O(N__28883),
            .I(N__28880));
    LocalMux I__4597 (
            .O(N__28880),
            .I(N__28877));
    Span4Mux_h I__4596 (
            .O(N__28877),
            .I(N__28874));
    Odrv4 I__4595 (
            .O(N__28874),
            .I(sDAC_mem_14Z0Z_2));
    CascadeMux I__4594 (
            .O(N__28871),
            .I(sDAC_data_RNO_18Z0Z_5_cascade_));
    InMux I__4593 (
            .O(N__28868),
            .I(N__28865));
    LocalMux I__4592 (
            .O(N__28865),
            .I(sDAC_data_RNO_19Z0Z_5));
    CascadeMux I__4591 (
            .O(N__28862),
            .I(sDAC_data_RNO_18Z0Z_6_cascade_));
    InMux I__4590 (
            .O(N__28859),
            .I(N__28856));
    LocalMux I__4589 (
            .O(N__28856),
            .I(N__28853));
    Span4Mux_h I__4588 (
            .O(N__28853),
            .I(N__28850));
    Odrv4 I__4587 (
            .O(N__28850),
            .I(sDAC_data_2_24_ns_1_6));
    InMux I__4586 (
            .O(N__28847),
            .I(N__28844));
    LocalMux I__4585 (
            .O(N__28844),
            .I(N__28841));
    Odrv12 I__4584 (
            .O(N__28841),
            .I(sDAC_mem_15Z0Z_3));
    InMux I__4583 (
            .O(N__28838),
            .I(N__28835));
    LocalMux I__4582 (
            .O(N__28835),
            .I(N__28832));
    Span4Mux_h I__4581 (
            .O(N__28832),
            .I(N__28829));
    Odrv4 I__4580 (
            .O(N__28829),
            .I(sDAC_mem_14Z0Z_3));
    InMux I__4579 (
            .O(N__28826),
            .I(N__28823));
    LocalMux I__4578 (
            .O(N__28823),
            .I(sDAC_data_RNO_19Z0Z_6));
    InMux I__4577 (
            .O(N__28820),
            .I(N__28817));
    LocalMux I__4576 (
            .O(N__28817),
            .I(sDAC_mem_12Z0Z_2));
    InMux I__4575 (
            .O(N__28814),
            .I(N__28811));
    LocalMux I__4574 (
            .O(N__28811),
            .I(sDAC_data_RNO_28Z0Z_8));
    InMux I__4573 (
            .O(N__28808),
            .I(N__28805));
    LocalMux I__4572 (
            .O(N__28805),
            .I(sDAC_mem_16Z0Z_5));
    InMux I__4571 (
            .O(N__28802),
            .I(N__28799));
    LocalMux I__4570 (
            .O(N__28799),
            .I(sDAC_mem_16Z0Z_6));
    CascadeMux I__4569 (
            .O(N__28796),
            .I(sDAC_data_RNO_10Z0Z_4_cascade_));
    InMux I__4568 (
            .O(N__28793),
            .I(N__28790));
    LocalMux I__4567 (
            .O(N__28790),
            .I(N__28787));
    Span4Mux_h I__4566 (
            .O(N__28787),
            .I(N__28784));
    Odrv4 I__4565 (
            .O(N__28784),
            .I(sDAC_data_RNO_11Z0Z_4));
    InMux I__4564 (
            .O(N__28781),
            .I(N__28778));
    LocalMux I__4563 (
            .O(N__28778),
            .I(N__28775));
    Span4Mux_h I__4562 (
            .O(N__28775),
            .I(N__28772));
    Odrv4 I__4561 (
            .O(N__28772),
            .I(sDAC_data_RNO_5Z0Z_4));
    InMux I__4560 (
            .O(N__28769),
            .I(N__28766));
    LocalMux I__4559 (
            .O(N__28766),
            .I(sDAC_data_RNO_2Z0Z_4));
    CascadeMux I__4558 (
            .O(N__28763),
            .I(sDAC_data_RNO_1Z0Z_4_cascade_));
    InMux I__4557 (
            .O(N__28760),
            .I(N__28757));
    LocalMux I__4556 (
            .O(N__28757),
            .I(sDAC_data_2_41_ns_1_4));
    CascadeMux I__4555 (
            .O(N__28754),
            .I(sDAC_data_2_4_cascade_));
    InMux I__4554 (
            .O(N__28751),
            .I(N__28748));
    LocalMux I__4553 (
            .O(N__28748),
            .I(sDAC_data_RNO_15Z0Z_4));
    InMux I__4552 (
            .O(N__28745),
            .I(N__28742));
    LocalMux I__4551 (
            .O(N__28742),
            .I(N__28739));
    Span4Mux_h I__4550 (
            .O(N__28739),
            .I(N__28736));
    Odrv4 I__4549 (
            .O(N__28736),
            .I(sDAC_mem_38Z0Z_3));
    InMux I__4548 (
            .O(N__28733),
            .I(N__28730));
    LocalMux I__4547 (
            .O(N__28730),
            .I(N__28727));
    Span4Mux_h I__4546 (
            .O(N__28727),
            .I(N__28724));
    Odrv4 I__4545 (
            .O(N__28724),
            .I(sDAC_mem_39Z0Z_3));
    CascadeMux I__4544 (
            .O(N__28721),
            .I(sDAC_data_2_13_bm_1_6_cascade_));
    InMux I__4543 (
            .O(N__28718),
            .I(N__28715));
    LocalMux I__4542 (
            .O(N__28715),
            .I(sDAC_data_RNO_5Z0Z_6));
    InMux I__4541 (
            .O(N__28712),
            .I(N__28709));
    LocalMux I__4540 (
            .O(N__28709),
            .I(sDAC_mem_6Z0Z_3));
    InMux I__4539 (
            .O(N__28706),
            .I(N__28703));
    LocalMux I__4538 (
            .O(N__28703),
            .I(N__28700));
    Odrv12 I__4537 (
            .O(N__28700),
            .I(sDAC_mem_38Z0Z_4));
    InMux I__4536 (
            .O(N__28697),
            .I(N__28694));
    LocalMux I__4535 (
            .O(N__28694),
            .I(N__28691));
    Span4Mux_v I__4534 (
            .O(N__28691),
            .I(N__28688));
    Sp12to4 I__4533 (
            .O(N__28688),
            .I(N__28685));
    Odrv12 I__4532 (
            .O(N__28685),
            .I(sDAC_mem_39Z0Z_4));
    CascadeMux I__4531 (
            .O(N__28682),
            .I(sDAC_data_2_13_bm_1_7_cascade_));
    InMux I__4530 (
            .O(N__28679),
            .I(N__28676));
    LocalMux I__4529 (
            .O(N__28676),
            .I(N__28673));
    Odrv4 I__4528 (
            .O(N__28673),
            .I(sDAC_data_RNO_28Z0Z_6));
    InMux I__4527 (
            .O(N__28670),
            .I(N__28667));
    LocalMux I__4526 (
            .O(N__28667),
            .I(sDAC_mem_16Z0Z_3));
    InMux I__4525 (
            .O(N__28664),
            .I(N__28661));
    LocalMux I__4524 (
            .O(N__28661),
            .I(sDAC_mem_16Z0Z_4));
    CascadeMux I__4523 (
            .O(N__28658),
            .I(sDAC_data_RNO_18Z0Z_8_cascade_));
    InMux I__4522 (
            .O(N__28655),
            .I(N__28652));
    LocalMux I__4521 (
            .O(N__28652),
            .I(sDAC_data_2_24_ns_1_8));
    InMux I__4520 (
            .O(N__28649),
            .I(N__28646));
    LocalMux I__4519 (
            .O(N__28646),
            .I(N__28643));
    Span4Mux_h I__4518 (
            .O(N__28643),
            .I(N__28640));
    Odrv4 I__4517 (
            .O(N__28640),
            .I(sDAC_mem_15Z0Z_5));
    InMux I__4516 (
            .O(N__28637),
            .I(N__28634));
    LocalMux I__4515 (
            .O(N__28634),
            .I(N__28631));
    Span4Mux_h I__4514 (
            .O(N__28631),
            .I(N__28628));
    Odrv4 I__4513 (
            .O(N__28628),
            .I(sDAC_mem_14Z0Z_5));
    InMux I__4512 (
            .O(N__28625),
            .I(N__28622));
    LocalMux I__4511 (
            .O(N__28622),
            .I(sDAC_data_RNO_19Z0Z_8));
    InMux I__4510 (
            .O(N__28619),
            .I(N__28616));
    LocalMux I__4509 (
            .O(N__28616),
            .I(sDAC_mem_12Z0Z_4));
    InMux I__4508 (
            .O(N__28613),
            .I(N__28610));
    LocalMux I__4507 (
            .O(N__28610),
            .I(sDAC_mem_12Z0Z_5));
    InMux I__4506 (
            .O(N__28607),
            .I(N__28604));
    LocalMux I__4505 (
            .O(N__28604),
            .I(N__28601));
    Odrv12 I__4504 (
            .O(N__28601),
            .I(sDAC_mem_38Z0Z_2));
    InMux I__4503 (
            .O(N__28598),
            .I(N__28595));
    LocalMux I__4502 (
            .O(N__28595),
            .I(N__28592));
    Span4Mux_h I__4501 (
            .O(N__28592),
            .I(N__28589));
    Odrv4 I__4500 (
            .O(N__28589),
            .I(sDAC_mem_39Z0Z_2));
    CascadeMux I__4499 (
            .O(N__28586),
            .I(sDAC_data_2_13_bm_1_5_cascade_));
    InMux I__4498 (
            .O(N__28583),
            .I(N__28580));
    LocalMux I__4497 (
            .O(N__28580),
            .I(sDAC_mem_6Z0Z_2));
    InMux I__4496 (
            .O(N__28577),
            .I(N__28574));
    LocalMux I__4495 (
            .O(N__28574),
            .I(sDAC_mem_18Z0Z_3));
    InMux I__4494 (
            .O(N__28571),
            .I(N__28568));
    LocalMux I__4493 (
            .O(N__28568),
            .I(sDAC_mem_18Z0Z_4));
    InMux I__4492 (
            .O(N__28565),
            .I(N__28562));
    LocalMux I__4491 (
            .O(N__28562),
            .I(N__28559));
    Odrv4 I__4490 (
            .O(N__28559),
            .I(sDAC_data_RNO_29Z0Z_8));
    InMux I__4489 (
            .O(N__28556),
            .I(N__28553));
    LocalMux I__4488 (
            .O(N__28553),
            .I(sDAC_mem_18Z0Z_5));
    InMux I__4487 (
            .O(N__28550),
            .I(N__28547));
    LocalMux I__4486 (
            .O(N__28547),
            .I(sDAC_mem_18Z0Z_6));
    CEMux I__4485 (
            .O(N__28544),
            .I(N__28541));
    LocalMux I__4484 (
            .O(N__28541),
            .I(N__28537));
    CEMux I__4483 (
            .O(N__28540),
            .I(N__28534));
    Span4Mux_h I__4482 (
            .O(N__28537),
            .I(N__28531));
    LocalMux I__4481 (
            .O(N__28534),
            .I(N__28528));
    Span4Mux_v I__4480 (
            .O(N__28531),
            .I(N__28523));
    Span4Mux_v I__4479 (
            .O(N__28528),
            .I(N__28523));
    Span4Mux_h I__4478 (
            .O(N__28523),
            .I(N__28520));
    Odrv4 I__4477 (
            .O(N__28520),
            .I(sDAC_mem_18_1_sqmuxa));
    InMux I__4476 (
            .O(N__28517),
            .I(N__28514));
    LocalMux I__4475 (
            .O(N__28514),
            .I(N__28511));
    Span12Mux_v I__4474 (
            .O(N__28511),
            .I(N__28508));
    Odrv12 I__4473 (
            .O(N__28508),
            .I(sDAC_mem_15Z0Z_4));
    InMux I__4472 (
            .O(N__28505),
            .I(N__28502));
    LocalMux I__4471 (
            .O(N__28502),
            .I(N__28499));
    Span4Mux_h I__4470 (
            .O(N__28499),
            .I(N__28496));
    Odrv4 I__4469 (
            .O(N__28496),
            .I(sDAC_mem_14Z0Z_4));
    CascadeMux I__4468 (
            .O(N__28493),
            .I(sDAC_data_RNO_18Z0Z_7_cascade_));
    InMux I__4467 (
            .O(N__28490),
            .I(N__28487));
    LocalMux I__4466 (
            .O(N__28487),
            .I(sDAC_data_RNO_19Z0Z_7));
    CEMux I__4465 (
            .O(N__28484),
            .I(N__28481));
    LocalMux I__4464 (
            .O(N__28481),
            .I(sDAC_mem_36_1_sqmuxa));
    InMux I__4463 (
            .O(N__28478),
            .I(N__28475));
    LocalMux I__4462 (
            .O(N__28475),
            .I(sDAC_data_RNO_29Z0Z_6));
    InMux I__4461 (
            .O(N__28472),
            .I(sRAM_pointer_read_cry_9));
    InMux I__4460 (
            .O(N__28469),
            .I(sRAM_pointer_read_cry_10));
    InMux I__4459 (
            .O(N__28466),
            .I(sRAM_pointer_read_cry_11));
    InMux I__4458 (
            .O(N__28463),
            .I(sRAM_pointer_read_cry_12));
    InMux I__4457 (
            .O(N__28460),
            .I(sRAM_pointer_read_cry_13));
    InMux I__4456 (
            .O(N__28457),
            .I(sRAM_pointer_read_cry_14));
    InMux I__4455 (
            .O(N__28454),
            .I(bfn_13_20_0_));
    InMux I__4454 (
            .O(N__28451),
            .I(sRAM_pointer_read_cry_16));
    InMux I__4453 (
            .O(N__28448),
            .I(sRAM_pointer_read_cry_17));
    CEMux I__4452 (
            .O(N__28445),
            .I(N__28436));
    CEMux I__4451 (
            .O(N__28444),
            .I(N__28436));
    CEMux I__4450 (
            .O(N__28443),
            .I(N__28436));
    GlobalMux I__4449 (
            .O(N__28436),
            .I(N__28433));
    gio2CtrlBuf I__4448 (
            .O(N__28433),
            .I(N_28_g));
    InMux I__4447 (
            .O(N__28430),
            .I(sRAM_pointer_read_cry_0));
    InMux I__4446 (
            .O(N__28427),
            .I(sRAM_pointer_read_cry_1));
    InMux I__4445 (
            .O(N__28424),
            .I(sRAM_pointer_read_cry_2));
    InMux I__4444 (
            .O(N__28421),
            .I(sRAM_pointer_read_cry_3));
    InMux I__4443 (
            .O(N__28418),
            .I(sRAM_pointer_read_cry_4));
    InMux I__4442 (
            .O(N__28415),
            .I(sRAM_pointer_read_cry_5));
    InMux I__4441 (
            .O(N__28412),
            .I(sRAM_pointer_read_cry_6));
    InMux I__4440 (
            .O(N__28409),
            .I(bfn_13_19_0_));
    InMux I__4439 (
            .O(N__28406),
            .I(sRAM_pointer_read_cry_8));
    InMux I__4438 (
            .O(N__28403),
            .I(N__28400));
    LocalMux I__4437 (
            .O(N__28400),
            .I(un1_sacqtime_cry_20_sf));
    InMux I__4436 (
            .O(N__28397),
            .I(N__28394));
    LocalMux I__4435 (
            .O(N__28394),
            .I(un1_sacqtime_cry_21_sf));
    InMux I__4434 (
            .O(N__28391),
            .I(N__28388));
    LocalMux I__4433 (
            .O(N__28388),
            .I(un1_sacqtime_cry_22_sf));
    InMux I__4432 (
            .O(N__28385),
            .I(N__28382));
    LocalMux I__4431 (
            .O(N__28382),
            .I(un1_sacqtime_cry_23_sf));
    InMux I__4430 (
            .O(N__28379),
            .I(bfn_13_17_0_));
    CascadeMux I__4429 (
            .O(N__28376),
            .I(N__28373));
    InMux I__4428 (
            .O(N__28373),
            .I(N__28367));
    InMux I__4427 (
            .O(N__28372),
            .I(N__28367));
    LocalMux I__4426 (
            .O(N__28367),
            .I(sADC_clk_prevZ0));
    CascadeMux I__4425 (
            .O(N__28364),
            .I(N_71_cascade_));
    InMux I__4424 (
            .O(N__28361),
            .I(bfn_13_18_0_));
    InMux I__4423 (
            .O(N__28358),
            .I(N__28354));
    CascadeMux I__4422 (
            .O(N__28357),
            .I(N__28351));
    LocalMux I__4421 (
            .O(N__28354),
            .I(N__28348));
    InMux I__4420 (
            .O(N__28351),
            .I(N__28345));
    Span4Mux_v I__4419 (
            .O(N__28348),
            .I(N__28342));
    LocalMux I__4418 (
            .O(N__28345),
            .I(sCounter_i_11));
    Odrv4 I__4417 (
            .O(N__28342),
            .I(sCounter_i_11));
    InMux I__4416 (
            .O(N__28337),
            .I(N__28333));
    InMux I__4415 (
            .O(N__28336),
            .I(N__28330));
    LocalMux I__4414 (
            .O(N__28333),
            .I(N__28327));
    LocalMux I__4413 (
            .O(N__28330),
            .I(N__28322));
    Span4Mux_v I__4412 (
            .O(N__28327),
            .I(N__28322));
    Odrv4 I__4411 (
            .O(N__28322),
            .I(sCounter_i_12));
    InMux I__4410 (
            .O(N__28319),
            .I(N__28315));
    CascadeMux I__4409 (
            .O(N__28318),
            .I(N__28312));
    LocalMux I__4408 (
            .O(N__28315),
            .I(N__28309));
    InMux I__4407 (
            .O(N__28312),
            .I(N__28306));
    Span4Mux_v I__4406 (
            .O(N__28309),
            .I(N__28303));
    LocalMux I__4405 (
            .O(N__28306),
            .I(sCounter_i_13));
    Odrv4 I__4404 (
            .O(N__28303),
            .I(sCounter_i_13));
    InMux I__4403 (
            .O(N__28298),
            .I(N__28294));
    CascadeMux I__4402 (
            .O(N__28297),
            .I(N__28291));
    LocalMux I__4401 (
            .O(N__28294),
            .I(N__28288));
    InMux I__4400 (
            .O(N__28291),
            .I(N__28285));
    Span4Mux_v I__4399 (
            .O(N__28288),
            .I(N__28282));
    LocalMux I__4398 (
            .O(N__28285),
            .I(sCounter_i_14));
    Odrv4 I__4397 (
            .O(N__28282),
            .I(sCounter_i_14));
    InMux I__4396 (
            .O(N__28277),
            .I(N__28274));
    LocalMux I__4395 (
            .O(N__28274),
            .I(N__28270));
    InMux I__4394 (
            .O(N__28273),
            .I(N__28267));
    Span4Mux_v I__4393 (
            .O(N__28270),
            .I(N__28264));
    LocalMux I__4392 (
            .O(N__28267),
            .I(sCounter_i_15));
    Odrv4 I__4391 (
            .O(N__28264),
            .I(sCounter_i_15));
    InMux I__4390 (
            .O(N__28259),
            .I(N__28256));
    LocalMux I__4389 (
            .O(N__28256),
            .I(un1_sacqtime_cry_16_sf));
    InMux I__4388 (
            .O(N__28253),
            .I(N__28250));
    LocalMux I__4387 (
            .O(N__28250),
            .I(un1_sacqtime_cry_17_sf));
    InMux I__4386 (
            .O(N__28247),
            .I(N__28244));
    LocalMux I__4385 (
            .O(N__28244),
            .I(un1_sacqtime_cry_18_sf));
    InMux I__4384 (
            .O(N__28241),
            .I(N__28238));
    LocalMux I__4383 (
            .O(N__28238),
            .I(un1_sacqtime_cry_19_sf));
    InMux I__4382 (
            .O(N__28235),
            .I(N__28231));
    CascadeMux I__4381 (
            .O(N__28234),
            .I(N__28228));
    LocalMux I__4380 (
            .O(N__28231),
            .I(N__28225));
    InMux I__4379 (
            .O(N__28228),
            .I(N__28222));
    Span4Mux_v I__4378 (
            .O(N__28225),
            .I(N__28219));
    LocalMux I__4377 (
            .O(N__28222),
            .I(sCounter_i_3));
    Odrv4 I__4376 (
            .O(N__28219),
            .I(sCounter_i_3));
    InMux I__4375 (
            .O(N__28214),
            .I(N__28210));
    CascadeMux I__4374 (
            .O(N__28213),
            .I(N__28207));
    LocalMux I__4373 (
            .O(N__28210),
            .I(N__28204));
    InMux I__4372 (
            .O(N__28207),
            .I(N__28201));
    Span4Mux_v I__4371 (
            .O(N__28204),
            .I(N__28198));
    LocalMux I__4370 (
            .O(N__28201),
            .I(sCounter_i_4));
    Odrv4 I__4369 (
            .O(N__28198),
            .I(sCounter_i_4));
    InMux I__4368 (
            .O(N__28193),
            .I(N__28190));
    LocalMux I__4367 (
            .O(N__28190),
            .I(N__28186));
    InMux I__4366 (
            .O(N__28189),
            .I(N__28183));
    Span4Mux_v I__4365 (
            .O(N__28186),
            .I(N__28180));
    LocalMux I__4364 (
            .O(N__28183),
            .I(sCounter_i_5));
    Odrv4 I__4363 (
            .O(N__28180),
            .I(sCounter_i_5));
    InMux I__4362 (
            .O(N__28175),
            .I(N__28171));
    CascadeMux I__4361 (
            .O(N__28174),
            .I(N__28168));
    LocalMux I__4360 (
            .O(N__28171),
            .I(N__28165));
    InMux I__4359 (
            .O(N__28168),
            .I(N__28162));
    Span4Mux_v I__4358 (
            .O(N__28165),
            .I(N__28159));
    LocalMux I__4357 (
            .O(N__28162),
            .I(sCounter_i_6));
    Odrv4 I__4356 (
            .O(N__28159),
            .I(sCounter_i_6));
    InMux I__4355 (
            .O(N__28154),
            .I(N__28151));
    LocalMux I__4354 (
            .O(N__28151),
            .I(N__28147));
    InMux I__4353 (
            .O(N__28150),
            .I(N__28144));
    Span4Mux_v I__4352 (
            .O(N__28147),
            .I(N__28141));
    LocalMux I__4351 (
            .O(N__28144),
            .I(sCounter_i_7));
    Odrv4 I__4350 (
            .O(N__28141),
            .I(sCounter_i_7));
    InMux I__4349 (
            .O(N__28136),
            .I(N__28132));
    CascadeMux I__4348 (
            .O(N__28135),
            .I(N__28129));
    LocalMux I__4347 (
            .O(N__28132),
            .I(N__28126));
    InMux I__4346 (
            .O(N__28129),
            .I(N__28123));
    Span4Mux_v I__4345 (
            .O(N__28126),
            .I(N__28120));
    LocalMux I__4344 (
            .O(N__28123),
            .I(sCounter_i_8));
    Odrv4 I__4343 (
            .O(N__28120),
            .I(sCounter_i_8));
    InMux I__4342 (
            .O(N__28115),
            .I(N__28112));
    LocalMux I__4341 (
            .O(N__28112),
            .I(N__28108));
    InMux I__4340 (
            .O(N__28111),
            .I(N__28105));
    Span4Mux_v I__4339 (
            .O(N__28108),
            .I(N__28102));
    LocalMux I__4338 (
            .O(N__28105),
            .I(sCounter_i_9));
    Odrv4 I__4337 (
            .O(N__28102),
            .I(sCounter_i_9));
    InMux I__4336 (
            .O(N__28097),
            .I(N__28093));
    CascadeMux I__4335 (
            .O(N__28096),
            .I(N__28090));
    LocalMux I__4334 (
            .O(N__28093),
            .I(N__28087));
    InMux I__4333 (
            .O(N__28090),
            .I(N__28084));
    Span4Mux_v I__4332 (
            .O(N__28087),
            .I(N__28081));
    LocalMux I__4331 (
            .O(N__28084),
            .I(sCounter_i_10));
    Odrv4 I__4330 (
            .O(N__28081),
            .I(sCounter_i_10));
    InMux I__4329 (
            .O(N__28076),
            .I(N__28073));
    LocalMux I__4328 (
            .O(N__28073),
            .I(sDAC_data_RNO_31Z0Z_5));
    InMux I__4327 (
            .O(N__28070),
            .I(N__28067));
    LocalMux I__4326 (
            .O(N__28067),
            .I(sDAC_mem_26Z0Z_2));
    InMux I__4325 (
            .O(N__28064),
            .I(N__28061));
    LocalMux I__4324 (
            .O(N__28061),
            .I(N__28058));
    Odrv4 I__4323 (
            .O(N__28058),
            .I(sDAC_data_RNO_31Z0Z_8));
    InMux I__4322 (
            .O(N__28055),
            .I(N__28052));
    LocalMux I__4321 (
            .O(N__28052),
            .I(sDAC_mem_26Z0Z_5));
    CEMux I__4320 (
            .O(N__28049),
            .I(N__28046));
    LocalMux I__4319 (
            .O(N__28046),
            .I(N__28042));
    CEMux I__4318 (
            .O(N__28045),
            .I(N__28039));
    Span4Mux_h I__4317 (
            .O(N__28042),
            .I(N__28034));
    LocalMux I__4316 (
            .O(N__28039),
            .I(N__28034));
    Span4Mux_v I__4315 (
            .O(N__28034),
            .I(N__28031));
    Span4Mux_h I__4314 (
            .O(N__28031),
            .I(N__28028));
    Odrv4 I__4313 (
            .O(N__28028),
            .I(sDAC_mem_26_1_sqmuxa));
    InMux I__4312 (
            .O(N__28025),
            .I(N__28022));
    LocalMux I__4311 (
            .O(N__28022),
            .I(N__28019));
    Span4Mux_h I__4310 (
            .O(N__28019),
            .I(N__28016));
    Span4Mux_v I__4309 (
            .O(N__28016),
            .I(N__28013));
    Span4Mux_v I__4308 (
            .O(N__28013),
            .I(N__28010));
    Odrv4 I__4307 (
            .O(N__28010),
            .I(\spi_master_inst.sclk_gen_u0.delay_clk_iZ0 ));
    InMux I__4306 (
            .O(N__28007),
            .I(N__28004));
    LocalMux I__4305 (
            .O(N__28004),
            .I(N__28001));
    Span4Mux_h I__4304 (
            .O(N__28001),
            .I(N__27997));
    InMux I__4303 (
            .O(N__28000),
            .I(N__27994));
    Span4Mux_h I__4302 (
            .O(N__27997),
            .I(N__27990));
    LocalMux I__4301 (
            .O(N__27994),
            .I(N__27986));
    InMux I__4300 (
            .O(N__27993),
            .I(N__27983));
    Span4Mux_v I__4299 (
            .O(N__27990),
            .I(N__27980));
    InMux I__4298 (
            .O(N__27989),
            .I(N__27977));
    Odrv4 I__4297 (
            .O(N__27986),
            .I(\spi_master_inst.sclk_gen_u0.div_clk_iZ0 ));
    LocalMux I__4296 (
            .O(N__27983),
            .I(\spi_master_inst.sclk_gen_u0.div_clk_iZ0 ));
    Odrv4 I__4295 (
            .O(N__27980),
            .I(\spi_master_inst.sclk_gen_u0.div_clk_iZ0 ));
    LocalMux I__4294 (
            .O(N__27977),
            .I(\spi_master_inst.sclk_gen_u0.div_clk_iZ0 ));
    CEMux I__4293 (
            .O(N__27968),
            .I(N__27965));
    LocalMux I__4292 (
            .O(N__27965),
            .I(N__27962));
    Odrv4 I__4291 (
            .O(N__27962),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i ));
    InMux I__4290 (
            .O(N__27959),
            .I(N__27953));
    InMux I__4289 (
            .O(N__27958),
            .I(N__27953));
    LocalMux I__4288 (
            .O(N__27953),
            .I(N__27950));
    Span4Mux_h I__4287 (
            .O(N__27950),
            .I(N__27947));
    Span4Mux_h I__4286 (
            .O(N__27947),
            .I(N__27944));
    Span4Mux_h I__4285 (
            .O(N__27944),
            .I(N__27940));
    InMux I__4284 (
            .O(N__27943),
            .I(N__27937));
    Span4Mux_v I__4283 (
            .O(N__27940),
            .I(N__27934));
    LocalMux I__4282 (
            .O(N__27937),
            .I(\spi_master_inst.sclk_gen_u0.falling_count_start_iZ0 ));
    Odrv4 I__4281 (
            .O(N__27934),
            .I(\spi_master_inst.sclk_gen_u0.falling_count_start_iZ0 ));
    InMux I__4280 (
            .O(N__27929),
            .I(N__27911));
    InMux I__4279 (
            .O(N__27928),
            .I(N__27911));
    InMux I__4278 (
            .O(N__27927),
            .I(N__27911));
    InMux I__4277 (
            .O(N__27926),
            .I(N__27911));
    InMux I__4276 (
            .O(N__27925),
            .I(N__27911));
    InMux I__4275 (
            .O(N__27924),
            .I(N__27904));
    InMux I__4274 (
            .O(N__27923),
            .I(N__27904));
    InMux I__4273 (
            .O(N__27922),
            .I(N__27904));
    LocalMux I__4272 (
            .O(N__27911),
            .I(N__27899));
    LocalMux I__4271 (
            .O(N__27904),
            .I(N__27899));
    Odrv4 I__4270 (
            .O(N__27899),
            .I(\spi_master_inst.sclk_gen_u0.falling_count_start_i_i ));
    InMux I__4269 (
            .O(N__27896),
            .I(N__27893));
    LocalMux I__4268 (
            .O(N__27893),
            .I(N__27889));
    InMux I__4267 (
            .O(N__27892),
            .I(N__27886));
    Span4Mux_v I__4266 (
            .O(N__27889),
            .I(N__27883));
    LocalMux I__4265 (
            .O(N__27886),
            .I(sCounter_i_0));
    Odrv4 I__4264 (
            .O(N__27883),
            .I(sCounter_i_0));
    InMux I__4263 (
            .O(N__27878),
            .I(N__27874));
    CascadeMux I__4262 (
            .O(N__27877),
            .I(N__27871));
    LocalMux I__4261 (
            .O(N__27874),
            .I(N__27868));
    InMux I__4260 (
            .O(N__27871),
            .I(N__27865));
    Span4Mux_v I__4259 (
            .O(N__27868),
            .I(N__27862));
    LocalMux I__4258 (
            .O(N__27865),
            .I(sCounter_i_1));
    Odrv4 I__4257 (
            .O(N__27862),
            .I(sCounter_i_1));
    InMux I__4256 (
            .O(N__27857),
            .I(N__27853));
    CascadeMux I__4255 (
            .O(N__27856),
            .I(N__27850));
    LocalMux I__4254 (
            .O(N__27853),
            .I(N__27847));
    InMux I__4253 (
            .O(N__27850),
            .I(N__27844));
    Span4Mux_v I__4252 (
            .O(N__27847),
            .I(N__27841));
    LocalMux I__4251 (
            .O(N__27844),
            .I(sCounter_i_2));
    Odrv4 I__4250 (
            .O(N__27841),
            .I(sCounter_i_2));
    InMux I__4249 (
            .O(N__27836),
            .I(N__27833));
    LocalMux I__4248 (
            .O(N__27833),
            .I(N__27830));
    Span4Mux_h I__4247 (
            .O(N__27830),
            .I(N__27827));
    Odrv4 I__4246 (
            .O(N__27827),
            .I(sDAC_mem_26Z0Z_1));
    CascadeMux I__4245 (
            .O(N__27824),
            .I(sDAC_data_RNO_30Z0Z_4_cascade_));
    InMux I__4244 (
            .O(N__27821),
            .I(N__27818));
    LocalMux I__4243 (
            .O(N__27818),
            .I(sDAC_data_RNO_31Z0Z_4));
    CascadeMux I__4242 (
            .O(N__27815),
            .I(sDAC_data_2_39_ns_1_4_cascade_));
    InMux I__4241 (
            .O(N__27812),
            .I(N__27809));
    LocalMux I__4240 (
            .O(N__27809),
            .I(N__27806));
    Span4Mux_h I__4239 (
            .O(N__27806),
            .I(N__27803));
    Odrv4 I__4238 (
            .O(N__27803),
            .I(sDAC_mem_28Z0Z_1));
    InMux I__4237 (
            .O(N__27800),
            .I(N__27797));
    LocalMux I__4236 (
            .O(N__27797),
            .I(N__27794));
    Span12Mux_h I__4235 (
            .O(N__27794),
            .I(N__27791));
    Odrv12 I__4234 (
            .O(N__27791),
            .I(sDAC_mem_29Z0Z_1));
    InMux I__4233 (
            .O(N__27788),
            .I(N__27785));
    LocalMux I__4232 (
            .O(N__27785),
            .I(sDAC_data_RNO_23Z0Z_4));
    InMux I__4231 (
            .O(N__27782),
            .I(N__27779));
    LocalMux I__4230 (
            .O(N__27779),
            .I(N__27776));
    Span4Mux_h I__4229 (
            .O(N__27776),
            .I(N__27773));
    Odrv4 I__4228 (
            .O(N__27773),
            .I(sDAC_mem_31Z0Z_1));
    InMux I__4227 (
            .O(N__27770),
            .I(N__27767));
    LocalMux I__4226 (
            .O(N__27767),
            .I(N__27764));
    Span12Mux_h I__4225 (
            .O(N__27764),
            .I(N__27761));
    Odrv12 I__4224 (
            .O(N__27761),
            .I(sDAC_mem_30Z0Z_1));
    InMux I__4223 (
            .O(N__27758),
            .I(N__27755));
    LocalMux I__4222 (
            .O(N__27755),
            .I(sDAC_data_RNO_24Z0Z_4));
    InMux I__4221 (
            .O(N__27752),
            .I(N__27749));
    LocalMux I__4220 (
            .O(N__27749),
            .I(sDAC_mem_24Z0Z_1));
    CEMux I__4219 (
            .O(N__27746),
            .I(N__27742));
    CEMux I__4218 (
            .O(N__27745),
            .I(N__27738));
    LocalMux I__4217 (
            .O(N__27742),
            .I(N__27735));
    CEMux I__4216 (
            .O(N__27741),
            .I(N__27732));
    LocalMux I__4215 (
            .O(N__27738),
            .I(N__27729));
    Span4Mux_v I__4214 (
            .O(N__27735),
            .I(N__27726));
    LocalMux I__4213 (
            .O(N__27732),
            .I(N__27723));
    Span4Mux_v I__4212 (
            .O(N__27729),
            .I(N__27720));
    Span4Mux_h I__4211 (
            .O(N__27726),
            .I(N__27715));
    Span4Mux_v I__4210 (
            .O(N__27723),
            .I(N__27715));
    Odrv4 I__4209 (
            .O(N__27720),
            .I(sDAC_mem_24_1_sqmuxa));
    Odrv4 I__4208 (
            .O(N__27715),
            .I(sDAC_mem_24_1_sqmuxa));
    InMux I__4207 (
            .O(N__27710),
            .I(N__27707));
    LocalMux I__4206 (
            .O(N__27707),
            .I(N__27704));
    Span4Mux_h I__4205 (
            .O(N__27704),
            .I(N__27701));
    Span4Mux_h I__4204 (
            .O(N__27701),
            .I(N__27698));
    Odrv4 I__4203 (
            .O(N__27698),
            .I(sDAC_mem_26Z0Z_6));
    InMux I__4202 (
            .O(N__27695),
            .I(N__27692));
    LocalMux I__4201 (
            .O(N__27692),
            .I(sDAC_data_RNO_31Z0Z_9));
    CascadeMux I__4200 (
            .O(N__27689),
            .I(sDAC_data_RNO_30Z0Z_7_cascade_));
    CascadeMux I__4199 (
            .O(N__27686),
            .I(sDAC_data_2_39_ns_1_7_cascade_));
    InMux I__4198 (
            .O(N__27683),
            .I(N__27680));
    LocalMux I__4197 (
            .O(N__27680),
            .I(N__27677));
    Span4Mux_h I__4196 (
            .O(N__27677),
            .I(N__27674));
    Odrv4 I__4195 (
            .O(N__27674),
            .I(sDAC_mem_26Z0Z_4));
    InMux I__4194 (
            .O(N__27671),
            .I(N__27668));
    LocalMux I__4193 (
            .O(N__27668),
            .I(sDAC_data_RNO_31Z0Z_7));
    InMux I__4192 (
            .O(N__27665),
            .I(N__27662));
    LocalMux I__4191 (
            .O(N__27662),
            .I(N__27659));
    Span4Mux_v I__4190 (
            .O(N__27659),
            .I(N__27656));
    Span4Mux_h I__4189 (
            .O(N__27656),
            .I(N__27653));
    Odrv4 I__4188 (
            .O(N__27653),
            .I(sDAC_mem_29Z0Z_4));
    InMux I__4187 (
            .O(N__27650),
            .I(N__27647));
    LocalMux I__4186 (
            .O(N__27647),
            .I(N__27644));
    Span4Mux_h I__4185 (
            .O(N__27644),
            .I(N__27641));
    Span4Mux_v I__4184 (
            .O(N__27641),
            .I(N__27638));
    Odrv4 I__4183 (
            .O(N__27638),
            .I(sDAC_mem_28Z0Z_4));
    InMux I__4182 (
            .O(N__27635),
            .I(N__27632));
    LocalMux I__4181 (
            .O(N__27632),
            .I(sDAC_data_RNO_23Z0Z_7));
    InMux I__4180 (
            .O(N__27629),
            .I(N__27626));
    LocalMux I__4179 (
            .O(N__27626),
            .I(N__27623));
    Span4Mux_h I__4178 (
            .O(N__27623),
            .I(N__27620));
    Odrv4 I__4177 (
            .O(N__27620),
            .I(sDAC_mem_30Z0Z_4));
    InMux I__4176 (
            .O(N__27617),
            .I(N__27614));
    LocalMux I__4175 (
            .O(N__27614),
            .I(N__27611));
    Span4Mux_v I__4174 (
            .O(N__27611),
            .I(N__27608));
    Span4Mux_h I__4173 (
            .O(N__27608),
            .I(N__27605));
    Odrv4 I__4172 (
            .O(N__27605),
            .I(sDAC_mem_31Z0Z_4));
    InMux I__4171 (
            .O(N__27602),
            .I(N__27599));
    LocalMux I__4170 (
            .O(N__27599),
            .I(sDAC_data_RNO_24Z0Z_7));
    InMux I__4169 (
            .O(N__27596),
            .I(N__27593));
    LocalMux I__4168 (
            .O(N__27593),
            .I(sDAC_mem_24Z0Z_4));
    InMux I__4167 (
            .O(N__27590),
            .I(N__27587));
    LocalMux I__4166 (
            .O(N__27587),
            .I(sDAC_data_2_39_ns_1_8));
    InMux I__4165 (
            .O(N__27584),
            .I(N__27581));
    LocalMux I__4164 (
            .O(N__27581),
            .I(sDAC_mem_12Z0Z_0));
    InMux I__4163 (
            .O(N__27578),
            .I(N__27575));
    LocalMux I__4162 (
            .O(N__27575),
            .I(sDAC_mem_12Z0Z_1));
    InMux I__4161 (
            .O(N__27572),
            .I(N__27569));
    LocalMux I__4160 (
            .O(N__27569),
            .I(N__27566));
    Span4Mux_h I__4159 (
            .O(N__27566),
            .I(N__27563));
    Odrv4 I__4158 (
            .O(N__27563),
            .I(sDAC_mem_31Z0Z_5));
    InMux I__4157 (
            .O(N__27560),
            .I(N__27557));
    LocalMux I__4156 (
            .O(N__27557),
            .I(N__27554));
    Span4Mux_h I__4155 (
            .O(N__27554),
            .I(N__27551));
    Span4Mux_v I__4154 (
            .O(N__27551),
            .I(N__27548));
    Odrv4 I__4153 (
            .O(N__27548),
            .I(sDAC_mem_30Z0Z_5));
    InMux I__4152 (
            .O(N__27545),
            .I(N__27542));
    LocalMux I__4151 (
            .O(N__27542),
            .I(N__27539));
    Span4Mux_v I__4150 (
            .O(N__27539),
            .I(N__27536));
    Span4Mux_h I__4149 (
            .O(N__27536),
            .I(N__27533));
    Odrv4 I__4148 (
            .O(N__27533),
            .I(sDAC_mem_29Z0Z_5));
    InMux I__4147 (
            .O(N__27530),
            .I(N__27527));
    LocalMux I__4146 (
            .O(N__27527),
            .I(sDAC_data_RNO_24Z0Z_8));
    CascadeMux I__4145 (
            .O(N__27524),
            .I(sDAC_data_RNO_23Z0Z_8_cascade_));
    InMux I__4144 (
            .O(N__27521),
            .I(N__27518));
    LocalMux I__4143 (
            .O(N__27518),
            .I(N__27515));
    Odrv4 I__4142 (
            .O(N__27515),
            .I(sDAC_data_RNO_11Z0Z_8));
    InMux I__4141 (
            .O(N__27512),
            .I(N__27509));
    LocalMux I__4140 (
            .O(N__27509),
            .I(sDAC_mem_28Z0Z_5));
    InMux I__4139 (
            .O(N__27506),
            .I(N__27503));
    LocalMux I__4138 (
            .O(N__27503),
            .I(N__27500));
    Span4Mux_v I__4137 (
            .O(N__27500),
            .I(N__27497));
    Span4Mux_h I__4136 (
            .O(N__27497),
            .I(N__27494));
    Odrv4 I__4135 (
            .O(N__27494),
            .I(sDAC_mem_24Z0Z_6));
    CascadeMux I__4134 (
            .O(N__27491),
            .I(sDAC_data_RNO_30Z0Z_9_cascade_));
    CascadeMux I__4133 (
            .O(N__27488),
            .I(sDAC_data_2_39_ns_1_9_cascade_));
    InMux I__4132 (
            .O(N__27485),
            .I(N__27482));
    LocalMux I__4131 (
            .O(N__27482),
            .I(N__27479));
    Odrv12 I__4130 (
            .O(N__27479),
            .I(sDAC_mem_40Z0Z_1));
    InMux I__4129 (
            .O(N__27476),
            .I(N__27473));
    LocalMux I__4128 (
            .O(N__27473),
            .I(N__27470));
    Span4Mux_v I__4127 (
            .O(N__27470),
            .I(N__27467));
    Odrv4 I__4126 (
            .O(N__27467),
            .I(sDAC_mem_8Z0Z_1));
    CascadeMux I__4125 (
            .O(N__27464),
            .I(sDAC_data_2_20_am_1_4_cascade_));
    CascadeMux I__4124 (
            .O(N__27461),
            .I(sDAC_data_RNO_7Z0Z_4_cascade_));
    InMux I__4123 (
            .O(N__27458),
            .I(N__27455));
    LocalMux I__4122 (
            .O(N__27455),
            .I(sDAC_data_RNO_8Z0Z_4));
    InMux I__4121 (
            .O(N__27452),
            .I(N__27449));
    LocalMux I__4120 (
            .O(N__27449),
            .I(N__27446));
    Odrv4 I__4119 (
            .O(N__27446),
            .I(sDAC_mem_15Z0Z_0));
    InMux I__4118 (
            .O(N__27443),
            .I(N__27440));
    LocalMux I__4117 (
            .O(N__27440),
            .I(N__27437));
    Span4Mux_v I__4116 (
            .O(N__27437),
            .I(N__27434));
    Odrv4 I__4115 (
            .O(N__27434),
            .I(sDAC_mem_14Z0Z_0));
    CascadeMux I__4114 (
            .O(N__27431),
            .I(sDAC_data_RNO_18Z0Z_3_cascade_));
    InMux I__4113 (
            .O(N__27428),
            .I(N__27425));
    LocalMux I__4112 (
            .O(N__27425),
            .I(sDAC_data_RNO_19Z0Z_3));
    CascadeMux I__4111 (
            .O(N__27422),
            .I(sDAC_data_RNO_18Z0Z_4_cascade_));
    InMux I__4110 (
            .O(N__27419),
            .I(N__27416));
    LocalMux I__4109 (
            .O(N__27416),
            .I(sDAC_data_2_24_ns_1_4));
    InMux I__4108 (
            .O(N__27413),
            .I(N__27410));
    LocalMux I__4107 (
            .O(N__27410),
            .I(N__27407));
    Odrv4 I__4106 (
            .O(N__27407),
            .I(sDAC_mem_15Z0Z_1));
    InMux I__4105 (
            .O(N__27404),
            .I(N__27401));
    LocalMux I__4104 (
            .O(N__27401),
            .I(N__27398));
    Span4Mux_v I__4103 (
            .O(N__27398),
            .I(N__27395));
    Odrv4 I__4102 (
            .O(N__27395),
            .I(sDAC_mem_14Z0Z_1));
    InMux I__4101 (
            .O(N__27392),
            .I(N__27389));
    LocalMux I__4100 (
            .O(N__27389),
            .I(sDAC_data_RNO_19Z0Z_4));
    CascadeMux I__4099 (
            .O(N__27386),
            .I(sDAC_data_2_8_cascade_));
    CascadeMux I__4098 (
            .O(N__27383),
            .I(sDAC_data_2_32_ns_1_8_cascade_));
    CascadeMux I__4097 (
            .O(N__27380),
            .I(sDAC_data_RNO_10Z0Z_8_cascade_));
    InMux I__4096 (
            .O(N__27377),
            .I(N__27374));
    LocalMux I__4095 (
            .O(N__27374),
            .I(sDAC_data_2_41_ns_1_8));
    InMux I__4094 (
            .O(N__27371),
            .I(N__27368));
    LocalMux I__4093 (
            .O(N__27368),
            .I(sDAC_mem_34Z0Z_1));
    InMux I__4092 (
            .O(N__27365),
            .I(N__27362));
    LocalMux I__4091 (
            .O(N__27362),
            .I(N__27359));
    Odrv4 I__4090 (
            .O(N__27359),
            .I(sDAC_mem_2Z0Z_1));
    InMux I__4089 (
            .O(N__27356),
            .I(N__27353));
    LocalMux I__4088 (
            .O(N__27353),
            .I(sDAC_mem_3Z0Z_1));
    InMux I__4087 (
            .O(N__27350),
            .I(N__27347));
    LocalMux I__4086 (
            .O(N__27347),
            .I(N__27344));
    Span4Mux_h I__4085 (
            .O(N__27344),
            .I(N__27341));
    Span4Mux_h I__4084 (
            .O(N__27341),
            .I(N__27338));
    Odrv4 I__4083 (
            .O(N__27338),
            .I(sDAC_mem_35Z0Z_1));
    CascadeMux I__4082 (
            .O(N__27335),
            .I(sDAC_data_2_6_bm_1_4_cascade_));
    InMux I__4081 (
            .O(N__27332),
            .I(N__27329));
    LocalMux I__4080 (
            .O(N__27329),
            .I(N__27326));
    Span4Mux_v I__4079 (
            .O(N__27326),
            .I(N__27323));
    Odrv4 I__4078 (
            .O(N__27323),
            .I(sDAC_mem_42Z0Z_1));
    InMux I__4077 (
            .O(N__27320),
            .I(N__27317));
    LocalMux I__4076 (
            .O(N__27317),
            .I(N__27314));
    Span4Mux_v I__4075 (
            .O(N__27314),
            .I(N__27311));
    Odrv4 I__4074 (
            .O(N__27311),
            .I(sDAC_mem_10Z0Z_1));
    CascadeMux I__4073 (
            .O(N__27308),
            .I(sDAC_data_RNO_17Z0Z_4_cascade_));
    InMux I__4072 (
            .O(N__27305),
            .I(N__27302));
    LocalMux I__4071 (
            .O(N__27302),
            .I(N__27299));
    Span4Mux_h I__4070 (
            .O(N__27299),
            .I(N__27296));
    Span4Mux_h I__4069 (
            .O(N__27296),
            .I(N__27293));
    Odrv4 I__4068 (
            .O(N__27293),
            .I(sDAC_mem_11Z0Z_1));
    InMux I__4067 (
            .O(N__27290),
            .I(N__27287));
    LocalMux I__4066 (
            .O(N__27287),
            .I(N__27284));
    Span4Mux_v I__4065 (
            .O(N__27284),
            .I(N__27281));
    Odrv4 I__4064 (
            .O(N__27281),
            .I(sDAC_mem_42Z0Z_5));
    InMux I__4063 (
            .O(N__27278),
            .I(N__27275));
    LocalMux I__4062 (
            .O(N__27275),
            .I(N__27272));
    Span4Mux_v I__4061 (
            .O(N__27272),
            .I(N__27269));
    Odrv4 I__4060 (
            .O(N__27269),
            .I(sDAC_mem_10Z0Z_5));
    CascadeMux I__4059 (
            .O(N__27266),
            .I(sDAC_data_RNO_17Z0Z_8_cascade_));
    InMux I__4058 (
            .O(N__27263),
            .I(N__27260));
    LocalMux I__4057 (
            .O(N__27260),
            .I(N__27257));
    Odrv12 I__4056 (
            .O(N__27257),
            .I(sDAC_mem_11Z0Z_5));
    InMux I__4055 (
            .O(N__27254),
            .I(N__27251));
    LocalMux I__4054 (
            .O(N__27251),
            .I(N__27248));
    Odrv4 I__4053 (
            .O(N__27248),
            .I(sDAC_mem_40Z0Z_5));
    InMux I__4052 (
            .O(N__27245),
            .I(N__27242));
    LocalMux I__4051 (
            .O(N__27242),
            .I(N__27239));
    Odrv4 I__4050 (
            .O(N__27239),
            .I(sDAC_mem_8Z0Z_5));
    CascadeMux I__4049 (
            .O(N__27236),
            .I(sDAC_data_2_20_am_1_8_cascade_));
    CascadeMux I__4048 (
            .O(N__27233),
            .I(sDAC_data_RNO_7Z0Z_8_cascade_));
    InMux I__4047 (
            .O(N__27230),
            .I(N__27227));
    LocalMux I__4046 (
            .O(N__27227),
            .I(sDAC_data_RNO_8Z0Z_8));
    InMux I__4045 (
            .O(N__27224),
            .I(N__27221));
    LocalMux I__4044 (
            .O(N__27221),
            .I(sDAC_data_RNO_15Z0Z_8));
    CascadeMux I__4043 (
            .O(N__27218),
            .I(sDAC_data_2_14_ns_1_8_cascade_));
    InMux I__4042 (
            .O(N__27215),
            .I(N__27212));
    LocalMux I__4041 (
            .O(N__27212),
            .I(sDAC_data_RNO_2Z0Z_8));
    CascadeMux I__4040 (
            .O(N__27209),
            .I(sDAC_data_RNO_1Z0Z_8_cascade_));
    CascadeMux I__4039 (
            .O(N__27206),
            .I(sDAC_data_2_32_ns_1_6_cascade_));
    InMux I__4038 (
            .O(N__27203),
            .I(N__27200));
    LocalMux I__4037 (
            .O(N__27200),
            .I(sDAC_data_RNO_15Z0Z_6));
    CascadeMux I__4036 (
            .O(N__27197),
            .I(sDAC_data_2_14_ns_1_6_cascade_));
    InMux I__4035 (
            .O(N__27194),
            .I(N__27191));
    LocalMux I__4034 (
            .O(N__27191),
            .I(sDAC_data_RNO_10Z0Z_6));
    InMux I__4033 (
            .O(N__27188),
            .I(N__27185));
    LocalMux I__4032 (
            .O(N__27185),
            .I(sDAC_data_RNO_2Z0Z_6));
    CascadeMux I__4031 (
            .O(N__27182),
            .I(sDAC_data_2_41_ns_1_6_cascade_));
    InMux I__4030 (
            .O(N__27179),
            .I(N__27176));
    LocalMux I__4029 (
            .O(N__27176),
            .I(sDAC_data_RNO_1Z0Z_6));
    CascadeMux I__4028 (
            .O(N__27173),
            .I(sDAC_data_2_6_cascade_));
    InMux I__4027 (
            .O(N__27170),
            .I(N__27167));
    LocalMux I__4026 (
            .O(N__27167),
            .I(N__27164));
    Odrv12 I__4025 (
            .O(N__27164),
            .I(sDAC_dataZ0Z_6));
    InMux I__4024 (
            .O(N__27161),
            .I(N__27158));
    LocalMux I__4023 (
            .O(N__27158),
            .I(N__27155));
    Span4Mux_h I__4022 (
            .O(N__27155),
            .I(N__27152));
    Odrv4 I__4021 (
            .O(N__27152),
            .I(sDAC_mem_34Z0Z_5));
    InMux I__4020 (
            .O(N__27149),
            .I(N__27146));
    LocalMux I__4019 (
            .O(N__27146),
            .I(sDAC_mem_2Z0Z_5));
    InMux I__4018 (
            .O(N__27143),
            .I(N__27140));
    LocalMux I__4017 (
            .O(N__27140),
            .I(N__27137));
    Odrv12 I__4016 (
            .O(N__27137),
            .I(sDAC_mem_35Z0Z_5));
    CascadeMux I__4015 (
            .O(N__27134),
            .I(sDAC_data_2_6_bm_1_8_cascade_));
    InMux I__4014 (
            .O(N__27131),
            .I(N__27128));
    LocalMux I__4013 (
            .O(N__27128),
            .I(sDAC_mem_3Z0Z_5));
    CEMux I__4012 (
            .O(N__27125),
            .I(N__27122));
    LocalMux I__4011 (
            .O(N__27122),
            .I(N__27119));
    Odrv12 I__4010 (
            .O(N__27119),
            .I(sDAC_mem_40_1_sqmuxa));
    CEMux I__4009 (
            .O(N__27116),
            .I(N__27113));
    LocalMux I__4008 (
            .O(N__27113),
            .I(sDAC_mem_8_1_sqmuxa));
    InMux I__4007 (
            .O(N__27110),
            .I(N__27107));
    LocalMux I__4006 (
            .O(N__27107),
            .I(N__27103));
    InMux I__4005 (
            .O(N__27106),
            .I(N__27100));
    Span4Mux_h I__4004 (
            .O(N__27103),
            .I(N__27095));
    LocalMux I__4003 (
            .O(N__27100),
            .I(N__27095));
    Span4Mux_h I__4002 (
            .O(N__27095),
            .I(N__27087));
    InMux I__4001 (
            .O(N__27094),
            .I(N__27084));
    InMux I__4000 (
            .O(N__27093),
            .I(N__27081));
    InMux I__3999 (
            .O(N__27092),
            .I(N__27078));
    InMux I__3998 (
            .O(N__27091),
            .I(N__27073));
    InMux I__3997 (
            .O(N__27090),
            .I(N__27073));
    Odrv4 I__3996 (
            .O(N__27087),
            .I(N_317));
    LocalMux I__3995 (
            .O(N__27084),
            .I(N_317));
    LocalMux I__3994 (
            .O(N__27081),
            .I(N_317));
    LocalMux I__3993 (
            .O(N__27078),
            .I(N_317));
    LocalMux I__3992 (
            .O(N__27073),
            .I(N_317));
    InMux I__3991 (
            .O(N__27062),
            .I(N__27058));
    CascadeMux I__3990 (
            .O(N__27061),
            .I(N__27054));
    LocalMux I__3989 (
            .O(N__27058),
            .I(N__27051));
    InMux I__3988 (
            .O(N__27057),
            .I(N__27046));
    InMux I__3987 (
            .O(N__27054),
            .I(N__27046));
    Span4Mux_v I__3986 (
            .O(N__27051),
            .I(N__27043));
    LocalMux I__3985 (
            .O(N__27046),
            .I(N__27040));
    Span4Mux_v I__3984 (
            .O(N__27043),
            .I(N__27037));
    Span4Mux_h I__3983 (
            .O(N__27040),
            .I(N__27034));
    Span4Mux_v I__3982 (
            .O(N__27037),
            .I(N__27031));
    Span4Mux_v I__3981 (
            .O(N__27034),
            .I(N__27028));
    Odrv4 I__3980 (
            .O(N__27031),
            .I(sAddress_RNI6VH7_4Z0Z_1));
    Odrv4 I__3979 (
            .O(N__27028),
            .I(sAddress_RNI6VH7_4Z0Z_1));
    CascadeMux I__3978 (
            .O(N__27023),
            .I(N__27016));
    InMux I__3977 (
            .O(N__27022),
            .I(N__27006));
    InMux I__3976 (
            .O(N__27021),
            .I(N__27006));
    InMux I__3975 (
            .O(N__27020),
            .I(N__27006));
    InMux I__3974 (
            .O(N__27019),
            .I(N__27006));
    InMux I__3973 (
            .O(N__27016),
            .I(N__27003));
    InMux I__3972 (
            .O(N__27015),
            .I(N__27000));
    LocalMux I__3971 (
            .O(N__27006),
            .I(N__26997));
    LocalMux I__3970 (
            .O(N__27003),
            .I(N__26992));
    LocalMux I__3969 (
            .O(N__27000),
            .I(N__26992));
    Span12Mux_v I__3968 (
            .O(N__26997),
            .I(N__26989));
    Odrv4 I__3967 (
            .O(N__26992),
            .I(sAddress_RNI70I7Z0Z_1));
    Odrv12 I__3966 (
            .O(N__26989),
            .I(sAddress_RNI70I7Z0Z_1));
    InMux I__3965 (
            .O(N__26984),
            .I(N__26981));
    LocalMux I__3964 (
            .O(N__26981),
            .I(N__26978));
    Span4Mux_h I__3963 (
            .O(N__26978),
            .I(N__26974));
    CascadeMux I__3962 (
            .O(N__26977),
            .I(N__26971));
    Span4Mux_v I__3961 (
            .O(N__26974),
            .I(N__26968));
    InMux I__3960 (
            .O(N__26971),
            .I(N__26965));
    Odrv4 I__3959 (
            .O(N__26968),
            .I(sAddress_RNIAM2A_0Z0Z_1));
    LocalMux I__3958 (
            .O(N__26965),
            .I(sAddress_RNIAM2A_0Z0Z_1));
    InMux I__3957 (
            .O(N__26960),
            .I(N__26957));
    LocalMux I__3956 (
            .O(N__26957),
            .I(N__26954));
    Span4Mux_v I__3955 (
            .O(N__26954),
            .I(N__26951));
    Span4Mux_h I__3954 (
            .O(N__26951),
            .I(N__26946));
    InMux I__3953 (
            .O(N__26950),
            .I(N__26943));
    InMux I__3952 (
            .O(N__26949),
            .I(N__26940));
    Odrv4 I__3951 (
            .O(N__26946),
            .I(sTrigCounterZ0Z_1));
    LocalMux I__3950 (
            .O(N__26943),
            .I(sTrigCounterZ0Z_1));
    LocalMux I__3949 (
            .O(N__26940),
            .I(sTrigCounterZ0Z_1));
    IoInMux I__3948 (
            .O(N__26933),
            .I(N__26930));
    LocalMux I__3947 (
            .O(N__26930),
            .I(N__26927));
    Span4Mux_s2_h I__3946 (
            .O(N__26927),
            .I(N__26924));
    Span4Mux_h I__3945 (
            .O(N__26924),
            .I(N__26921));
    Sp12to4 I__3944 (
            .O(N__26921),
            .I(N__26918));
    Span12Mux_v I__3943 (
            .O(N__26918),
            .I(N__26915));
    Odrv12 I__3942 (
            .O(N__26915),
            .I(RAM_DATA_1Z0Z_14));
    InMux I__3941 (
            .O(N__26912),
            .I(N__26909));
    LocalMux I__3940 (
            .O(N__26909),
            .I(N__26906));
    Span4Mux_v I__3939 (
            .O(N__26906),
            .I(N__26903));
    Sp12to4 I__3938 (
            .O(N__26903),
            .I(N__26900));
    Span12Mux_h I__3937 (
            .O(N__26900),
            .I(N__26897));
    Odrv12 I__3936 (
            .O(N__26897),
            .I(ADC2_c));
    IoInMux I__3935 (
            .O(N__26894),
            .I(N__26891));
    LocalMux I__3934 (
            .O(N__26891),
            .I(N__26888));
    Span12Mux_s8_v I__3933 (
            .O(N__26888),
            .I(N__26885));
    Span12Mux_h I__3932 (
            .O(N__26885),
            .I(N__26882));
    Odrv12 I__3931 (
            .O(N__26882),
            .I(RAM_DATA_1Z0Z_2));
    InMux I__3930 (
            .O(N__26879),
            .I(N__26876));
    LocalMux I__3929 (
            .O(N__26876),
            .I(N__26873));
    Span4Mux_v I__3928 (
            .O(N__26873),
            .I(N__26870));
    Sp12to4 I__3927 (
            .O(N__26870),
            .I(N__26867));
    Span12Mux_h I__3926 (
            .O(N__26867),
            .I(N__26864));
    Odrv12 I__3925 (
            .O(N__26864),
            .I(ADC6_c));
    IoInMux I__3924 (
            .O(N__26861),
            .I(N__26858));
    LocalMux I__3923 (
            .O(N__26858),
            .I(N__26855));
    Span4Mux_s2_v I__3922 (
            .O(N__26855),
            .I(N__26852));
    Span4Mux_h I__3921 (
            .O(N__26852),
            .I(N__26849));
    Span4Mux_v I__3920 (
            .O(N__26849),
            .I(N__26846));
    Sp12to4 I__3919 (
            .O(N__26846),
            .I(N__26843));
    Odrv12 I__3918 (
            .O(N__26843),
            .I(RAM_DATA_1Z0Z_6));
    InMux I__3917 (
            .O(N__26840),
            .I(N__26837));
    LocalMux I__3916 (
            .O(N__26837),
            .I(N__26834));
    Span4Mux_v I__3915 (
            .O(N__26834),
            .I(N__26831));
    Span4Mux_h I__3914 (
            .O(N__26831),
            .I(N__26828));
    Span4Mux_h I__3913 (
            .O(N__26828),
            .I(N__26825));
    Odrv4 I__3912 (
            .O(N__26825),
            .I(ADC0_c));
    IoInMux I__3911 (
            .O(N__26822),
            .I(N__26819));
    LocalMux I__3910 (
            .O(N__26819),
            .I(N__26816));
    Span4Mux_s2_v I__3909 (
            .O(N__26816),
            .I(N__26813));
    Span4Mux_v I__3908 (
            .O(N__26813),
            .I(N__26810));
    Sp12to4 I__3907 (
            .O(N__26810),
            .I(N__26807));
    Odrv12 I__3906 (
            .O(N__26807),
            .I(RAM_DATA_1Z0Z_0));
    InMux I__3905 (
            .O(N__26804),
            .I(N__26801));
    LocalMux I__3904 (
            .O(N__26801),
            .I(N__26798));
    Odrv4 I__3903 (
            .O(N__26798),
            .I(sDAC_mem_40Z0Z_3));
    CascadeMux I__3902 (
            .O(N__26795),
            .I(N__26792));
    InMux I__3901 (
            .O(N__26792),
            .I(N__26789));
    LocalMux I__3900 (
            .O(N__26789),
            .I(N__26786));
    Span12Mux_v I__3899 (
            .O(N__26786),
            .I(N__26783));
    Odrv12 I__3898 (
            .O(N__26783),
            .I(sEEPoffZ0Z_15));
    InMux I__3897 (
            .O(N__26780),
            .I(N__26777));
    LocalMux I__3896 (
            .O(N__26777),
            .I(N__26774));
    Span4Mux_v I__3895 (
            .O(N__26774),
            .I(N__26771));
    Odrv4 I__3894 (
            .O(N__26771),
            .I(sEEPoffZ0Z_8));
    CascadeMux I__3893 (
            .O(N__26768),
            .I(N__26765));
    InMux I__3892 (
            .O(N__26765),
            .I(N__26762));
    LocalMux I__3891 (
            .O(N__26762),
            .I(N__26759));
    Odrv12 I__3890 (
            .O(N__26759),
            .I(sEEPoffZ0Z_9));
    CEMux I__3889 (
            .O(N__26756),
            .I(N__26752));
    CEMux I__3888 (
            .O(N__26755),
            .I(N__26749));
    LocalMux I__3887 (
            .O(N__26752),
            .I(sAddress_RNIA6242_2Z0Z_0));
    LocalMux I__3886 (
            .O(N__26749),
            .I(sAddress_RNIA6242_2Z0Z_0));
    IoInMux I__3885 (
            .O(N__26744),
            .I(N__26741));
    LocalMux I__3884 (
            .O(N__26741),
            .I(N__26738));
    IoSpan4Mux I__3883 (
            .O(N__26738),
            .I(N__26735));
    Span4Mux_s3_h I__3882 (
            .O(N__26735),
            .I(N__26732));
    Span4Mux_h I__3881 (
            .O(N__26732),
            .I(N__26729));
    Span4Mux_h I__3880 (
            .O(N__26729),
            .I(N__26726));
    Span4Mux_h I__3879 (
            .O(N__26726),
            .I(N__26723));
    Odrv4 I__3878 (
            .O(N__26723),
            .I(un4_sacqtime_cry_23_c_RNI2CQMZ0));
    InMux I__3877 (
            .O(N__26720),
            .I(N__26717));
    LocalMux I__3876 (
            .O(N__26717),
            .I(N__26714));
    Span4Mux_v I__3875 (
            .O(N__26714),
            .I(N__26711));
    Sp12to4 I__3874 (
            .O(N__26711),
            .I(N__26708));
    Span12Mux_h I__3873 (
            .O(N__26708),
            .I(N__26705));
    Odrv12 I__3872 (
            .O(N__26705),
            .I(ADC5_c));
    IoInMux I__3871 (
            .O(N__26702),
            .I(N__26699));
    LocalMux I__3870 (
            .O(N__26699),
            .I(N__26696));
    IoSpan4Mux I__3869 (
            .O(N__26696),
            .I(N__26693));
    IoSpan4Mux I__3868 (
            .O(N__26693),
            .I(N__26690));
    Span4Mux_s2_v I__3867 (
            .O(N__26690),
            .I(N__26687));
    Sp12to4 I__3866 (
            .O(N__26687),
            .I(N__26684));
    Span12Mux_s8_v I__3865 (
            .O(N__26684),
            .I(N__26681));
    Odrv12 I__3864 (
            .O(N__26681),
            .I(RAM_DATA_1Z0Z_5));
    InMux I__3863 (
            .O(N__26678),
            .I(N__26675));
    LocalMux I__3862 (
            .O(N__26675),
            .I(N__26672));
    Span4Mux_v I__3861 (
            .O(N__26672),
            .I(N__26669));
    Sp12to4 I__3860 (
            .O(N__26669),
            .I(N__26666));
    Span12Mux_h I__3859 (
            .O(N__26666),
            .I(N__26663));
    Odrv12 I__3858 (
            .O(N__26663),
            .I(ADC1_c));
    IoInMux I__3857 (
            .O(N__26660),
            .I(N__26657));
    LocalMux I__3856 (
            .O(N__26657),
            .I(N__26654));
    Span12Mux_s11_v I__3855 (
            .O(N__26654),
            .I(N__26651));
    Span12Mux_h I__3854 (
            .O(N__26651),
            .I(N__26648));
    Odrv12 I__3853 (
            .O(N__26648),
            .I(RAM_DATA_1Z0Z_1));
    InMux I__3852 (
            .O(N__26645),
            .I(N__26642));
    LocalMux I__3851 (
            .O(N__26642),
            .I(N__26639));
    Span4Mux_v I__3850 (
            .O(N__26639),
            .I(N__26636));
    Sp12to4 I__3849 (
            .O(N__26636),
            .I(N__26633));
    Span12Mux_h I__3848 (
            .O(N__26633),
            .I(N__26630));
    Odrv12 I__3847 (
            .O(N__26630),
            .I(ADC9_c));
    IoInMux I__3846 (
            .O(N__26627),
            .I(N__26624));
    LocalMux I__3845 (
            .O(N__26624),
            .I(N__26621));
    Span12Mux_s4_h I__3844 (
            .O(N__26621),
            .I(N__26618));
    Span12Mux_v I__3843 (
            .O(N__26618),
            .I(N__26615));
    Span12Mux_h I__3842 (
            .O(N__26615),
            .I(N__26612));
    Odrv12 I__3841 (
            .O(N__26612),
            .I(RAM_DATA_1Z0Z_10));
    InMux I__3840 (
            .O(N__26609),
            .I(N__26606));
    LocalMux I__3839 (
            .O(N__26606),
            .I(N__26603));
    Span12Mux_v I__3838 (
            .O(N__26603),
            .I(N__26600));
    Span12Mux_h I__3837 (
            .O(N__26600),
            .I(N__26597));
    Odrv12 I__3836 (
            .O(N__26597),
            .I(top_tour1_c));
    IoInMux I__3835 (
            .O(N__26594),
            .I(N__26591));
    LocalMux I__3834 (
            .O(N__26591),
            .I(N__26588));
    IoSpan4Mux I__3833 (
            .O(N__26588),
            .I(N__26585));
    Span4Mux_s2_h I__3832 (
            .O(N__26585),
            .I(N__26582));
    Sp12to4 I__3831 (
            .O(N__26582),
            .I(N__26579));
    Span12Mux_h I__3830 (
            .O(N__26579),
            .I(N__26576));
    Odrv12 I__3829 (
            .O(N__26576),
            .I(RAM_DATA_1Z0Z_11));
    InMux I__3828 (
            .O(N__26573),
            .I(N__26570));
    LocalMux I__3827 (
            .O(N__26570),
            .I(N__26567));
    Span4Mux_v I__3826 (
            .O(N__26567),
            .I(N__26564));
    Span4Mux_h I__3825 (
            .O(N__26564),
            .I(N__26559));
    InMux I__3824 (
            .O(N__26563),
            .I(N__26556));
    InMux I__3823 (
            .O(N__26562),
            .I(N__26553));
    Odrv4 I__3822 (
            .O(N__26559),
            .I(sTrigCounterZ0Z_0));
    LocalMux I__3821 (
            .O(N__26556),
            .I(sTrigCounterZ0Z_0));
    LocalMux I__3820 (
            .O(N__26553),
            .I(sTrigCounterZ0Z_0));
    IoInMux I__3819 (
            .O(N__26546),
            .I(N__26543));
    LocalMux I__3818 (
            .O(N__26543),
            .I(N__26540));
    IoSpan4Mux I__3817 (
            .O(N__26540),
            .I(N__26537));
    Span4Mux_s2_h I__3816 (
            .O(N__26537),
            .I(N__26534));
    Sp12to4 I__3815 (
            .O(N__26534),
            .I(N__26531));
    Span12Mux_h I__3814 (
            .O(N__26531),
            .I(N__26528));
    Odrv12 I__3813 (
            .O(N__26528),
            .I(RAM_DATA_1Z0Z_13));
    CEMux I__3812 (
            .O(N__26525),
            .I(N__26522));
    LocalMux I__3811 (
            .O(N__26522),
            .I(N__26519));
    Odrv12 I__3810 (
            .O(N__26519),
            .I(sAddress_RNIA6242_0Z0Z_0));
    InMux I__3809 (
            .O(N__26516),
            .I(N__26513));
    LocalMux I__3808 (
            .O(N__26513),
            .I(N__26510));
    Span4Mux_v I__3807 (
            .O(N__26510),
            .I(N__26507));
    Odrv4 I__3806 (
            .O(N__26507),
            .I(sEEPoffZ0Z_11));
    CascadeMux I__3805 (
            .O(N__26504),
            .I(N__26501));
    InMux I__3804 (
            .O(N__26501),
            .I(N__26498));
    LocalMux I__3803 (
            .O(N__26498),
            .I(N__26495));
    Odrv12 I__3802 (
            .O(N__26495),
            .I(sEEPoffZ0Z_12));
    InMux I__3801 (
            .O(N__26492),
            .I(N__26489));
    LocalMux I__3800 (
            .O(N__26489),
            .I(N__26486));
    Span4Mux_v I__3799 (
            .O(N__26486),
            .I(N__26483));
    Odrv4 I__3798 (
            .O(N__26483),
            .I(sEEPoffZ0Z_13));
    InMux I__3797 (
            .O(N__26480),
            .I(N__26477));
    LocalMux I__3796 (
            .O(N__26477),
            .I(N__26474));
    Odrv12 I__3795 (
            .O(N__26474),
            .I(sEEPoffZ0Z_14));
    CEMux I__3794 (
            .O(N__26471),
            .I(N__26468));
    LocalMux I__3793 (
            .O(N__26468),
            .I(N__26465));
    Span4Mux_v I__3792 (
            .O(N__26465),
            .I(N__26462));
    Span4Mux_h I__3791 (
            .O(N__26462),
            .I(N__26459));
    Odrv4 I__3790 (
            .O(N__26459),
            .I(sAddress_RNIA6242_1Z0Z_0));
    InMux I__3789 (
            .O(N__26456),
            .I(N__26453));
    LocalMux I__3788 (
            .O(N__26453),
            .I(sCounter_i_19));
    InMux I__3787 (
            .O(N__26450),
            .I(N__26447));
    LocalMux I__3786 (
            .O(N__26447),
            .I(sCounter_i_20));
    InMux I__3785 (
            .O(N__26444),
            .I(N__26441));
    LocalMux I__3784 (
            .O(N__26441),
            .I(sCounter_i_21));
    InMux I__3783 (
            .O(N__26438),
            .I(N__26435));
    LocalMux I__3782 (
            .O(N__26435),
            .I(sCounter_i_22));
    InMux I__3781 (
            .O(N__26432),
            .I(N__26429));
    LocalMux I__3780 (
            .O(N__26429),
            .I(sCounter_i_23));
    InMux I__3779 (
            .O(N__26426),
            .I(bfn_12_13_0_));
    IoInMux I__3778 (
            .O(N__26423),
            .I(N__26420));
    LocalMux I__3777 (
            .O(N__26420),
            .I(N__26417));
    IoSpan4Mux I__3776 (
            .O(N__26417),
            .I(N__26414));
    Span4Mux_s1_h I__3775 (
            .O(N__26414),
            .I(N__26411));
    Span4Mux_h I__3774 (
            .O(N__26411),
            .I(N__26408));
    Span4Mux_h I__3773 (
            .O(N__26408),
            .I(N__26405));
    Span4Mux_h I__3772 (
            .O(N__26405),
            .I(N__26402));
    Odrv4 I__3771 (
            .O(N__26402),
            .I(N_1683_i));
    InMux I__3770 (
            .O(N__26399),
            .I(N__26396));
    LocalMux I__3769 (
            .O(N__26396),
            .I(N__26393));
    Span4Mux_v I__3768 (
            .O(N__26393),
            .I(N__26390));
    Span4Mux_h I__3767 (
            .O(N__26390),
            .I(N__26386));
    CascadeMux I__3766 (
            .O(N__26389),
            .I(N__26383));
    Span4Mux_h I__3765 (
            .O(N__26386),
            .I(N__26380));
    InMux I__3764 (
            .O(N__26383),
            .I(N__26377));
    Odrv4 I__3763 (
            .O(N__26380),
            .I(sbuttonModeStatusZ0));
    LocalMux I__3762 (
            .O(N__26377),
            .I(sbuttonModeStatusZ0));
    InMux I__3761 (
            .O(N__26372),
            .I(N__26369));
    LocalMux I__3760 (
            .O(N__26369),
            .I(N__26366));
    Odrv4 I__3759 (
            .O(N__26366),
            .I(sbuttonModeStatus_0_sqmuxa_0));
    InMux I__3758 (
            .O(N__26363),
            .I(N__26360));
    LocalMux I__3757 (
            .O(N__26360),
            .I(sbuttonModeStatus_0_sqmuxa_18));
    InMux I__3756 (
            .O(N__26357),
            .I(N__26354));
    LocalMux I__3755 (
            .O(N__26354),
            .I(sCounter_i_16));
    InMux I__3754 (
            .O(N__26351),
            .I(N__26348));
    LocalMux I__3753 (
            .O(N__26348),
            .I(sCounter_i_17));
    InMux I__3752 (
            .O(N__26345),
            .I(N__26342));
    LocalMux I__3751 (
            .O(N__26342),
            .I(sCounter_i_18));
    InMux I__3750 (
            .O(N__26339),
            .I(N__26336));
    LocalMux I__3749 (
            .O(N__26336),
            .I(N__26333));
    Span4Mux_v I__3748 (
            .O(N__26333),
            .I(N__26330));
    Odrv4 I__3747 (
            .O(N__26330),
            .I(sEEPoffZ0Z_2));
    InMux I__3746 (
            .O(N__26327),
            .I(N__26324));
    LocalMux I__3745 (
            .O(N__26324),
            .I(N__26321));
    Span4Mux_v I__3744 (
            .O(N__26321),
            .I(N__26318));
    Odrv4 I__3743 (
            .O(N__26318),
            .I(sEEPoffZ0Z_3));
    InMux I__3742 (
            .O(N__26315),
            .I(N__26312));
    LocalMux I__3741 (
            .O(N__26312),
            .I(N__26309));
    Span4Mux_v I__3740 (
            .O(N__26309),
            .I(N__26306));
    Odrv4 I__3739 (
            .O(N__26306),
            .I(sEEPoffZ0Z_4));
    CascadeMux I__3738 (
            .O(N__26303),
            .I(N__26300));
    InMux I__3737 (
            .O(N__26300),
            .I(N__26297));
    LocalMux I__3736 (
            .O(N__26297),
            .I(N__26294));
    Span4Mux_v I__3735 (
            .O(N__26294),
            .I(N__26291));
    Odrv4 I__3734 (
            .O(N__26291),
            .I(sEEPoffZ0Z_5));
    InMux I__3733 (
            .O(N__26288),
            .I(N__26285));
    LocalMux I__3732 (
            .O(N__26285),
            .I(N__26282));
    Span4Mux_v I__3731 (
            .O(N__26282),
            .I(N__26279));
    Odrv4 I__3730 (
            .O(N__26279),
            .I(sEEPoffZ0Z_6));
    CascadeMux I__3729 (
            .O(N__26276),
            .I(N__26273));
    InMux I__3728 (
            .O(N__26273),
            .I(N__26270));
    LocalMux I__3727 (
            .O(N__26270),
            .I(N__26267));
    Span4Mux_v I__3726 (
            .O(N__26267),
            .I(N__26264));
    Odrv4 I__3725 (
            .O(N__26264),
            .I(sEEPoffZ0Z_7));
    InMux I__3724 (
            .O(N__26261),
            .I(N__26258));
    LocalMux I__3723 (
            .O(N__26258),
            .I(N__26255));
    Span4Mux_v I__3722 (
            .O(N__26255),
            .I(N__26252));
    Odrv4 I__3721 (
            .O(N__26252),
            .I(sEEPoffZ0Z_10));
    InMux I__3720 (
            .O(N__26249),
            .I(N__26246));
    LocalMux I__3719 (
            .O(N__26246),
            .I(N__26243));
    Odrv12 I__3718 (
            .O(N__26243),
            .I(sDAC_mem_39Z0Z_1));
    CEMux I__3717 (
            .O(N__26240),
            .I(N__26237));
    LocalMux I__3716 (
            .O(N__26237),
            .I(N__26234));
    Span4Mux_v I__3715 (
            .O(N__26234),
            .I(N__26231));
    Span4Mux_h I__3714 (
            .O(N__26231),
            .I(N__26228));
    Odrv4 I__3713 (
            .O(N__26228),
            .I(sDAC_mem_39_1_sqmuxa));
    CascadeMux I__3712 (
            .O(N__26225),
            .I(N__26222));
    InMux I__3711 (
            .O(N__26222),
            .I(N__26219));
    LocalMux I__3710 (
            .O(N__26219),
            .I(N__26216));
    Span4Mux_v I__3709 (
            .O(N__26216),
            .I(N__26213));
    Odrv4 I__3708 (
            .O(N__26213),
            .I(sEEPoffZ0Z_0));
    InMux I__3707 (
            .O(N__26210),
            .I(N__26207));
    LocalMux I__3706 (
            .O(N__26207),
            .I(N__26204));
    Span4Mux_v I__3705 (
            .O(N__26204),
            .I(N__26201));
    Odrv4 I__3704 (
            .O(N__26201),
            .I(sEEPoffZ0Z_1));
    InMux I__3703 (
            .O(N__26198),
            .I(N__26188));
    InMux I__3702 (
            .O(N__26197),
            .I(N__26188));
    InMux I__3701 (
            .O(N__26196),
            .I(N__26185));
    InMux I__3700 (
            .O(N__26195),
            .I(N__26179));
    InMux I__3699 (
            .O(N__26194),
            .I(N__26179));
    CascadeMux I__3698 (
            .O(N__26193),
            .I(N__26175));
    LocalMux I__3697 (
            .O(N__26188),
            .I(N__26171));
    LocalMux I__3696 (
            .O(N__26185),
            .I(N__26168));
    CascadeMux I__3695 (
            .O(N__26184),
            .I(N__26159));
    LocalMux I__3694 (
            .O(N__26179),
            .I(N__26156));
    InMux I__3693 (
            .O(N__26178),
            .I(N__26153));
    InMux I__3692 (
            .O(N__26175),
            .I(N__26148));
    InMux I__3691 (
            .O(N__26174),
            .I(N__26148));
    Span12Mux_s11_h I__3690 (
            .O(N__26171),
            .I(N__26145));
    Span4Mux_v I__3689 (
            .O(N__26168),
            .I(N__26142));
    InMux I__3688 (
            .O(N__26167),
            .I(N__26137));
    InMux I__3687 (
            .O(N__26166),
            .I(N__26137));
    InMux I__3686 (
            .O(N__26165),
            .I(N__26134));
    InMux I__3685 (
            .O(N__26164),
            .I(N__26131));
    InMux I__3684 (
            .O(N__26163),
            .I(N__26124));
    InMux I__3683 (
            .O(N__26162),
            .I(N__26124));
    InMux I__3682 (
            .O(N__26159),
            .I(N__26124));
    Span4Mux_v I__3681 (
            .O(N__26156),
            .I(N__26121));
    LocalMux I__3680 (
            .O(N__26153),
            .I(N__26118));
    LocalMux I__3679 (
            .O(N__26148),
            .I(sPointerZ0Z_1));
    Odrv12 I__3678 (
            .O(N__26145),
            .I(sPointerZ0Z_1));
    Odrv4 I__3677 (
            .O(N__26142),
            .I(sPointerZ0Z_1));
    LocalMux I__3676 (
            .O(N__26137),
            .I(sPointerZ0Z_1));
    LocalMux I__3675 (
            .O(N__26134),
            .I(sPointerZ0Z_1));
    LocalMux I__3674 (
            .O(N__26131),
            .I(sPointerZ0Z_1));
    LocalMux I__3673 (
            .O(N__26124),
            .I(sPointerZ0Z_1));
    Odrv4 I__3672 (
            .O(N__26121),
            .I(sPointerZ0Z_1));
    Odrv4 I__3671 (
            .O(N__26118),
            .I(sPointerZ0Z_1));
    InMux I__3670 (
            .O(N__26099),
            .I(N__26095));
    InMux I__3669 (
            .O(N__26098),
            .I(N__26092));
    LocalMux I__3668 (
            .O(N__26095),
            .I(N__26084));
    LocalMux I__3667 (
            .O(N__26092),
            .I(N__26081));
    InMux I__3666 (
            .O(N__26091),
            .I(N__26078));
    InMux I__3665 (
            .O(N__26090),
            .I(N__26073));
    InMux I__3664 (
            .O(N__26089),
            .I(N__26073));
    InMux I__3663 (
            .O(N__26088),
            .I(N__26068));
    InMux I__3662 (
            .O(N__26087),
            .I(N__26068));
    Span4Mux_h I__3661 (
            .O(N__26084),
            .I(N__26065));
    Span4Mux_v I__3660 (
            .O(N__26081),
            .I(N__26062));
    LocalMux I__3659 (
            .O(N__26078),
            .I(N__26059));
    LocalMux I__3658 (
            .O(N__26073),
            .I(sPointerZ0Z_0));
    LocalMux I__3657 (
            .O(N__26068),
            .I(sPointerZ0Z_0));
    Odrv4 I__3656 (
            .O(N__26065),
            .I(sPointerZ0Z_0));
    Odrv4 I__3655 (
            .O(N__26062),
            .I(sPointerZ0Z_0));
    Odrv4 I__3654 (
            .O(N__26059),
            .I(sPointerZ0Z_0));
    InMux I__3653 (
            .O(N__26048),
            .I(N__26045));
    LocalMux I__3652 (
            .O(N__26045),
            .I(N__26038));
    InMux I__3651 (
            .O(N__26044),
            .I(N__26031));
    InMux I__3650 (
            .O(N__26043),
            .I(N__26031));
    InMux I__3649 (
            .O(N__26042),
            .I(N__26031));
    InMux I__3648 (
            .O(N__26041),
            .I(N__26028));
    Span4Mux_v I__3647 (
            .O(N__26038),
            .I(N__26024));
    LocalMux I__3646 (
            .O(N__26031),
            .I(N__26019));
    LocalMux I__3645 (
            .O(N__26028),
            .I(N__26019));
    InMux I__3644 (
            .O(N__26027),
            .I(N__26016));
    Span4Mux_h I__3643 (
            .O(N__26024),
            .I(N__26009));
    Span4Mux_v I__3642 (
            .O(N__26019),
            .I(N__26009));
    LocalMux I__3641 (
            .O(N__26016),
            .I(N__26009));
    Odrv4 I__3640 (
            .O(N__26009),
            .I(spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1));
    InMux I__3639 (
            .O(N__26006),
            .I(N__26003));
    LocalMux I__3638 (
            .O(N__26003),
            .I(N__26000));
    Span4Mux_h I__3637 (
            .O(N__26000),
            .I(N__25997));
    Span4Mux_h I__3636 (
            .O(N__25997),
            .I(N__25994));
    Odrv4 I__3635 (
            .O(N__25994),
            .I(N_1624));
    InMux I__3634 (
            .O(N__25991),
            .I(N__25988));
    LocalMux I__3633 (
            .O(N__25988),
            .I(N__25985));
    Odrv4 I__3632 (
            .O(N__25985),
            .I(sDAC_mem_34Z0Z_3));
    CEMux I__3631 (
            .O(N__25982),
            .I(N__25979));
    LocalMux I__3630 (
            .O(N__25979),
            .I(N__25976));
    Span4Mux_h I__3629 (
            .O(N__25976),
            .I(N__25973));
    Odrv4 I__3628 (
            .O(N__25973),
            .I(sDAC_mem_34_1_sqmuxa));
    InMux I__3627 (
            .O(N__25970),
            .I(N__25967));
    LocalMux I__3626 (
            .O(N__25967),
            .I(sDAC_mem_7Z0Z_1));
    InMux I__3625 (
            .O(N__25964),
            .I(N__25961));
    LocalMux I__3624 (
            .O(N__25961),
            .I(N__25958));
    Span4Mux_v I__3623 (
            .O(N__25958),
            .I(N__25955));
    Odrv4 I__3622 (
            .O(N__25955),
            .I(un1_spointer11_2_0_0_a2_5));
    InMux I__3621 (
            .O(N__25952),
            .I(N__25949));
    LocalMux I__3620 (
            .O(N__25949),
            .I(N__25946));
    Span4Mux_h I__3619 (
            .O(N__25946),
            .I(N__25942));
    InMux I__3618 (
            .O(N__25945),
            .I(N__25939));
    Span4Mux_h I__3617 (
            .O(N__25942),
            .I(N__25936));
    LocalMux I__3616 (
            .O(N__25939),
            .I(N__25933));
    Odrv4 I__3615 (
            .O(N__25936),
            .I(N_183));
    Odrv12 I__3614 (
            .O(N__25933),
            .I(N_183));
    InMux I__3613 (
            .O(N__25928),
            .I(N__25925));
    LocalMux I__3612 (
            .O(N__25925),
            .I(sDAC_mem_8Z0Z_3));
    CascadeMux I__3611 (
            .O(N__25922),
            .I(sDAC_data_2_20_am_1_6_cascade_));
    InMux I__3610 (
            .O(N__25919),
            .I(N__25916));
    LocalMux I__3609 (
            .O(N__25916),
            .I(N__25913));
    Odrv4 I__3608 (
            .O(N__25913),
            .I(sDAC_mem_10Z0Z_3));
    InMux I__3607 (
            .O(N__25910),
            .I(N__25907));
    LocalMux I__3606 (
            .O(N__25907),
            .I(N__25904));
    Odrv12 I__3605 (
            .O(N__25904),
            .I(sDAC_mem_42Z0Z_3));
    CascadeMux I__3604 (
            .O(N__25901),
            .I(sDAC_data_RNO_17Z0Z_6_cascade_));
    InMux I__3603 (
            .O(N__25898),
            .I(N__25895));
    LocalMux I__3602 (
            .O(N__25895),
            .I(N__25892));
    Span4Mux_v I__3601 (
            .O(N__25892),
            .I(N__25889));
    Odrv4 I__3600 (
            .O(N__25889),
            .I(sDAC_mem_11Z0Z_3));
    CascadeMux I__3599 (
            .O(N__25886),
            .I(sDAC_data_RNO_8Z0Z_6_cascade_));
    InMux I__3598 (
            .O(N__25883),
            .I(N__25880));
    LocalMux I__3597 (
            .O(N__25880),
            .I(sDAC_data_RNO_7Z0Z_6));
    InMux I__3596 (
            .O(N__25877),
            .I(N__25874));
    LocalMux I__3595 (
            .O(N__25874),
            .I(sDAC_mem_2Z0Z_3));
    InMux I__3594 (
            .O(N__25871),
            .I(N__25868));
    LocalMux I__3593 (
            .O(N__25868),
            .I(N__25865));
    Span12Mux_s11_v I__3592 (
            .O(N__25865),
            .I(N__25862));
    Odrv12 I__3591 (
            .O(N__25862),
            .I(sDAC_mem_35Z0Z_3));
    CascadeMux I__3590 (
            .O(N__25859),
            .I(sDAC_data_2_6_bm_1_6_cascade_));
    InMux I__3589 (
            .O(N__25856),
            .I(N__25853));
    LocalMux I__3588 (
            .O(N__25853),
            .I(sDAC_mem_3Z0Z_3));
    InMux I__3587 (
            .O(N__25850),
            .I(N__25847));
    LocalMux I__3586 (
            .O(N__25847),
            .I(N__25844));
    Span4Mux_h I__3585 (
            .O(N__25844),
            .I(N__25841));
    Span4Mux_v I__3584 (
            .O(N__25841),
            .I(N__25838));
    Odrv4 I__3583 (
            .O(N__25838),
            .I(g0_4_0));
    InMux I__3582 (
            .O(N__25835),
            .I(bfn_11_20_0_));
    InMux I__3581 (
            .O(N__25832),
            .I(N__25829));
    LocalMux I__3580 (
            .O(N__25829),
            .I(N__25826));
    Sp12to4 I__3579 (
            .O(N__25826),
            .I(N__25823));
    Span12Mux_h I__3578 (
            .O(N__25823),
            .I(N__25820));
    Odrv12 I__3577 (
            .O(N__25820),
            .I(spi_sclk_ft_c));
    InMux I__3576 (
            .O(N__25817),
            .I(N__25814));
    LocalMux I__3575 (
            .O(N__25814),
            .I(N__25811));
    Span4Mux_v I__3574 (
            .O(N__25811),
            .I(N__25808));
    Sp12to4 I__3573 (
            .O(N__25808),
            .I(N__25805));
    Span12Mux_h I__3572 (
            .O(N__25805),
            .I(N__25802));
    Odrv12 I__3571 (
            .O(N__25802),
            .I(spi_sclk_rpi_c));
    IoInMux I__3570 (
            .O(N__25799),
            .I(N__25796));
    LocalMux I__3569 (
            .O(N__25796),
            .I(N__25793));
    Odrv12 I__3568 (
            .O(N__25793),
            .I(spi_sclk));
    InMux I__3567 (
            .O(N__25790),
            .I(N__25787));
    LocalMux I__3566 (
            .O(N__25787),
            .I(N__25784));
    Span4Mux_h I__3565 (
            .O(N__25784),
            .I(N__25781));
    Odrv4 I__3564 (
            .O(N__25781),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3 ));
    InMux I__3563 (
            .O(N__25778),
            .I(N__25775));
    LocalMux I__3562 (
            .O(N__25775),
            .I(N__25772));
    Span4Mux_h I__3561 (
            .O(N__25772),
            .I(N__25769));
    Odrv4 I__3560 (
            .O(N__25769),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_12 ));
    InMux I__3559 (
            .O(N__25766),
            .I(N__25763));
    LocalMux I__3558 (
            .O(N__25763),
            .I(N__25760));
    Span4Mux_h I__3557 (
            .O(N__25760),
            .I(N__25757));
    Odrv4 I__3556 (
            .O(N__25757),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12 ));
    InMux I__3555 (
            .O(N__25754),
            .I(N__25751));
    LocalMux I__3554 (
            .O(N__25751),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7 ));
    InMux I__3553 (
            .O(N__25748),
            .I(N__25745));
    LocalMux I__3552 (
            .O(N__25745),
            .I(N__25742));
    Odrv12 I__3551 (
            .O(N__25742),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9 ));
    InMux I__3550 (
            .O(N__25739),
            .I(N__25736));
    LocalMux I__3549 (
            .O(N__25736),
            .I(sEEDelayACQZ0Z_14));
    InMux I__3548 (
            .O(N__25733),
            .I(N__25730));
    LocalMux I__3547 (
            .O(N__25730),
            .I(sEEDelayACQ_i_14));
    InMux I__3546 (
            .O(N__25727),
            .I(N__25724));
    LocalMux I__3545 (
            .O(N__25724),
            .I(sEEDelayACQZ0Z_15));
    CascadeMux I__3544 (
            .O(N__25721),
            .I(N__25718));
    InMux I__3543 (
            .O(N__25718),
            .I(N__25715));
    LocalMux I__3542 (
            .O(N__25715),
            .I(sEEDelayACQ_i_15));
    InMux I__3541 (
            .O(N__25712),
            .I(N__25709));
    LocalMux I__3540 (
            .O(N__25709),
            .I(N__25706));
    Span4Mux_h I__3539 (
            .O(N__25706),
            .I(N__25703));
    Span4Mux_v I__3538 (
            .O(N__25703),
            .I(N__25700));
    Odrv4 I__3537 (
            .O(N__25700),
            .I(g1_i_a4_4));
    InMux I__3536 (
            .O(N__25697),
            .I(N__25694));
    LocalMux I__3535 (
            .O(N__25694),
            .I(sEEDelayACQZ0Z_6));
    InMux I__3534 (
            .O(N__25691),
            .I(N__25688));
    LocalMux I__3533 (
            .O(N__25688),
            .I(sEEDelayACQ_i_6));
    InMux I__3532 (
            .O(N__25685),
            .I(N__25682));
    LocalMux I__3531 (
            .O(N__25682),
            .I(sEEDelayACQZ0Z_7));
    CascadeMux I__3530 (
            .O(N__25679),
            .I(N__25676));
    InMux I__3529 (
            .O(N__25676),
            .I(N__25673));
    LocalMux I__3528 (
            .O(N__25673),
            .I(sEEDelayACQ_i_7));
    InMux I__3527 (
            .O(N__25670),
            .I(N__25667));
    LocalMux I__3526 (
            .O(N__25667),
            .I(sEEDelayACQZ0Z_8));
    InMux I__3525 (
            .O(N__25664),
            .I(N__25661));
    LocalMux I__3524 (
            .O(N__25661),
            .I(sEEDelayACQ_i_8));
    InMux I__3523 (
            .O(N__25658),
            .I(N__25655));
    LocalMux I__3522 (
            .O(N__25655),
            .I(sEEDelayACQZ0Z_9));
    InMux I__3521 (
            .O(N__25652),
            .I(N__25649));
    LocalMux I__3520 (
            .O(N__25649),
            .I(sEEDelayACQ_i_9));
    InMux I__3519 (
            .O(N__25646),
            .I(N__25643));
    LocalMux I__3518 (
            .O(N__25643),
            .I(sEEDelayACQZ0Z_10));
    InMux I__3517 (
            .O(N__25640),
            .I(N__25637));
    LocalMux I__3516 (
            .O(N__25637),
            .I(sEEDelayACQ_i_10));
    InMux I__3515 (
            .O(N__25634),
            .I(N__25631));
    LocalMux I__3514 (
            .O(N__25631),
            .I(sEEDelayACQZ0Z_11));
    InMux I__3513 (
            .O(N__25628),
            .I(N__25625));
    LocalMux I__3512 (
            .O(N__25625),
            .I(sEEDelayACQ_i_11));
    InMux I__3511 (
            .O(N__25622),
            .I(N__25619));
    LocalMux I__3510 (
            .O(N__25619),
            .I(sEEDelayACQZ0Z_12));
    InMux I__3509 (
            .O(N__25616),
            .I(N__25613));
    LocalMux I__3508 (
            .O(N__25613),
            .I(sEEDelayACQ_i_12));
    InMux I__3507 (
            .O(N__25610),
            .I(N__25607));
    LocalMux I__3506 (
            .O(N__25607),
            .I(sEEDelayACQZ0Z_13));
    InMux I__3505 (
            .O(N__25604),
            .I(N__25601));
    LocalMux I__3504 (
            .O(N__25601),
            .I(sEEDelayACQ_i_13));
    InMux I__3503 (
            .O(N__25598),
            .I(N__25595));
    LocalMux I__3502 (
            .O(N__25595),
            .I(sEEDelayACQZ0Z_0));
    InMux I__3501 (
            .O(N__25592),
            .I(N__25589));
    LocalMux I__3500 (
            .O(N__25589),
            .I(sEEDelayACQ_i_0));
    InMux I__3499 (
            .O(N__25586),
            .I(N__25583));
    LocalMux I__3498 (
            .O(N__25583),
            .I(sEEDelayACQZ0Z_1));
    InMux I__3497 (
            .O(N__25580),
            .I(N__25577));
    LocalMux I__3496 (
            .O(N__25577),
            .I(sEEDelayACQ_i_1));
    InMux I__3495 (
            .O(N__25574),
            .I(N__25571));
    LocalMux I__3494 (
            .O(N__25571),
            .I(sEEDelayACQZ0Z_2));
    InMux I__3493 (
            .O(N__25568),
            .I(N__25565));
    LocalMux I__3492 (
            .O(N__25565),
            .I(sEEDelayACQ_i_2));
    InMux I__3491 (
            .O(N__25562),
            .I(N__25559));
    LocalMux I__3490 (
            .O(N__25559),
            .I(sEEDelayACQZ0Z_3));
    CascadeMux I__3489 (
            .O(N__25556),
            .I(N__25553));
    InMux I__3488 (
            .O(N__25553),
            .I(N__25550));
    LocalMux I__3487 (
            .O(N__25550),
            .I(sEEDelayACQ_i_3));
    InMux I__3486 (
            .O(N__25547),
            .I(N__25544));
    LocalMux I__3485 (
            .O(N__25544),
            .I(sEEDelayACQZ0Z_4));
    InMux I__3484 (
            .O(N__25541),
            .I(N__25538));
    LocalMux I__3483 (
            .O(N__25538),
            .I(sEEDelayACQ_i_4));
    InMux I__3482 (
            .O(N__25535),
            .I(N__25532));
    LocalMux I__3481 (
            .O(N__25532),
            .I(sEEDelayACQZ0Z_5));
    InMux I__3480 (
            .O(N__25529),
            .I(N__25526));
    LocalMux I__3479 (
            .O(N__25526),
            .I(sEEDelayACQ_i_5));
    InMux I__3478 (
            .O(N__25523),
            .I(N__25517));
    InMux I__3477 (
            .O(N__25522),
            .I(N__25510));
    InMux I__3476 (
            .O(N__25521),
            .I(N__25510));
    InMux I__3475 (
            .O(N__25520),
            .I(N__25510));
    LocalMux I__3474 (
            .O(N__25517),
            .I(N__25505));
    LocalMux I__3473 (
            .O(N__25510),
            .I(N__25505));
    Span4Mux_h I__3472 (
            .O(N__25505),
            .I(N__25502));
    Span4Mux_v I__3471 (
            .O(N__25502),
            .I(N__25499));
    Odrv4 I__3470 (
            .O(N__25499),
            .I(un1_spointer11_5_0_2));
    CEMux I__3469 (
            .O(N__25496),
            .I(N__25493));
    LocalMux I__3468 (
            .O(N__25493),
            .I(sAddress_RNIA6242_3Z0Z_0));
    InMux I__3467 (
            .O(N__25490),
            .I(N__25486));
    InMux I__3466 (
            .O(N__25489),
            .I(N__25483));
    LocalMux I__3465 (
            .O(N__25486),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2 ));
    LocalMux I__3464 (
            .O(N__25483),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2 ));
    InMux I__3463 (
            .O(N__25478),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1 ));
    InMux I__3462 (
            .O(N__25475),
            .I(N__25471));
    InMux I__3461 (
            .O(N__25474),
            .I(N__25468));
    LocalMux I__3460 (
            .O(N__25471),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3 ));
    LocalMux I__3459 (
            .O(N__25468),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3 ));
    InMux I__3458 (
            .O(N__25463),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2 ));
    InMux I__3457 (
            .O(N__25460),
            .I(N__25457));
    LocalMux I__3456 (
            .O(N__25457),
            .I(N__25454));
    Span4Mux_h I__3455 (
            .O(N__25454),
            .I(N__25450));
    InMux I__3454 (
            .O(N__25453),
            .I(N__25447));
    Span4Mux_h I__3453 (
            .O(N__25450),
            .I(N__25444));
    LocalMux I__3452 (
            .O(N__25447),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4 ));
    Odrv4 I__3451 (
            .O(N__25444),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4 ));
    InMux I__3450 (
            .O(N__25439),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3 ));
    CascadeMux I__3449 (
            .O(N__25436),
            .I(N__25432));
    InMux I__3448 (
            .O(N__25435),
            .I(N__25429));
    InMux I__3447 (
            .O(N__25432),
            .I(N__25426));
    LocalMux I__3446 (
            .O(N__25429),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5 ));
    LocalMux I__3445 (
            .O(N__25426),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5 ));
    InMux I__3444 (
            .O(N__25421),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4 ));
    InMux I__3443 (
            .O(N__25418),
            .I(N__25414));
    InMux I__3442 (
            .O(N__25417),
            .I(N__25411));
    LocalMux I__3441 (
            .O(N__25414),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6 ));
    LocalMux I__3440 (
            .O(N__25411),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6 ));
    InMux I__3439 (
            .O(N__25406),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5 ));
    InMux I__3438 (
            .O(N__25403),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6 ));
    InMux I__3437 (
            .O(N__25400),
            .I(N__25396));
    InMux I__3436 (
            .O(N__25399),
            .I(N__25393));
    LocalMux I__3435 (
            .O(N__25396),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7 ));
    LocalMux I__3434 (
            .O(N__25393),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7 ));
    InMux I__3433 (
            .O(N__25388),
            .I(sCounter_cry_16));
    InMux I__3432 (
            .O(N__25385),
            .I(sCounter_cry_17));
    InMux I__3431 (
            .O(N__25382),
            .I(sCounter_cry_18));
    InMux I__3430 (
            .O(N__25379),
            .I(sCounter_cry_19));
    InMux I__3429 (
            .O(N__25376),
            .I(sCounter_cry_20));
    InMux I__3428 (
            .O(N__25373),
            .I(sCounter_cry_21));
    InMux I__3427 (
            .O(N__25370),
            .I(N__25340));
    InMux I__3426 (
            .O(N__25369),
            .I(N__25340));
    InMux I__3425 (
            .O(N__25368),
            .I(N__25340));
    InMux I__3424 (
            .O(N__25367),
            .I(N__25331));
    InMux I__3423 (
            .O(N__25366),
            .I(N__25331));
    InMux I__3422 (
            .O(N__25365),
            .I(N__25331));
    InMux I__3421 (
            .O(N__25364),
            .I(N__25331));
    InMux I__3420 (
            .O(N__25363),
            .I(N__25322));
    InMux I__3419 (
            .O(N__25362),
            .I(N__25322));
    InMux I__3418 (
            .O(N__25361),
            .I(N__25322));
    InMux I__3417 (
            .O(N__25360),
            .I(N__25322));
    InMux I__3416 (
            .O(N__25359),
            .I(N__25311));
    InMux I__3415 (
            .O(N__25358),
            .I(N__25311));
    InMux I__3414 (
            .O(N__25357),
            .I(N__25311));
    InMux I__3413 (
            .O(N__25356),
            .I(N__25311));
    InMux I__3412 (
            .O(N__25355),
            .I(N__25311));
    InMux I__3411 (
            .O(N__25354),
            .I(N__25302));
    InMux I__3410 (
            .O(N__25353),
            .I(N__25302));
    InMux I__3409 (
            .O(N__25352),
            .I(N__25302));
    InMux I__3408 (
            .O(N__25351),
            .I(N__25302));
    InMux I__3407 (
            .O(N__25350),
            .I(N__25293));
    InMux I__3406 (
            .O(N__25349),
            .I(N__25293));
    InMux I__3405 (
            .O(N__25348),
            .I(N__25293));
    InMux I__3404 (
            .O(N__25347),
            .I(N__25293));
    LocalMux I__3403 (
            .O(N__25340),
            .I(N__25288));
    LocalMux I__3402 (
            .O(N__25331),
            .I(N__25288));
    LocalMux I__3401 (
            .O(N__25322),
            .I(N__25281));
    LocalMux I__3400 (
            .O(N__25311),
            .I(N__25281));
    LocalMux I__3399 (
            .O(N__25302),
            .I(N__25281));
    LocalMux I__3398 (
            .O(N__25293),
            .I(LED_ACQ_c_i));
    Odrv4 I__3397 (
            .O(N__25288),
            .I(LED_ACQ_c_i));
    Odrv4 I__3396 (
            .O(N__25281),
            .I(LED_ACQ_c_i));
    InMux I__3395 (
            .O(N__25274),
            .I(sCounter_cry_22));
    InMux I__3394 (
            .O(N__25271),
            .I(N__25267));
    InMux I__3393 (
            .O(N__25270),
            .I(N__25264));
    LocalMux I__3392 (
            .O(N__25267),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0 ));
    LocalMux I__3391 (
            .O(N__25264),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0 ));
    InMux I__3390 (
            .O(N__25259),
            .I(bfn_11_13_0_));
    InMux I__3389 (
            .O(N__25256),
            .I(N__25252));
    InMux I__3388 (
            .O(N__25255),
            .I(N__25249));
    LocalMux I__3387 (
            .O(N__25252),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1 ));
    LocalMux I__3386 (
            .O(N__25249),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1 ));
    InMux I__3385 (
            .O(N__25244),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0 ));
    InMux I__3384 (
            .O(N__25241),
            .I(bfn_11_11_0_));
    InMux I__3383 (
            .O(N__25238),
            .I(sCounter_cry_8));
    InMux I__3382 (
            .O(N__25235),
            .I(sCounter_cry_9));
    InMux I__3381 (
            .O(N__25232),
            .I(sCounter_cry_10));
    InMux I__3380 (
            .O(N__25229),
            .I(sCounter_cry_11));
    InMux I__3379 (
            .O(N__25226),
            .I(sCounter_cry_12));
    InMux I__3378 (
            .O(N__25223),
            .I(sCounter_cry_13));
    InMux I__3377 (
            .O(N__25220),
            .I(sCounter_cry_14));
    InMux I__3376 (
            .O(N__25217),
            .I(bfn_11_12_0_));
    InMux I__3375 (
            .O(N__25214),
            .I(N__25210));
    InMux I__3374 (
            .O(N__25213),
            .I(N__25207));
    LocalMux I__3373 (
            .O(N__25210),
            .I(N__25203));
    LocalMux I__3372 (
            .O(N__25207),
            .I(N__25200));
    InMux I__3371 (
            .O(N__25206),
            .I(N__25197));
    Span4Mux_v I__3370 (
            .O(N__25203),
            .I(N__25194));
    Odrv4 I__3369 (
            .O(N__25200),
            .I(sTrigInternalZ0));
    LocalMux I__3368 (
            .O(N__25197),
            .I(sTrigInternalZ0));
    Odrv4 I__3367 (
            .O(N__25194),
            .I(sTrigInternalZ0));
    CascadeMux I__3366 (
            .O(N__25187),
            .I(N__25184));
    InMux I__3365 (
            .O(N__25184),
            .I(N__25180));
    InMux I__3364 (
            .O(N__25183),
            .I(N__25177));
    LocalMux I__3363 (
            .O(N__25180),
            .I(N__25174));
    LocalMux I__3362 (
            .O(N__25177),
            .I(N__25171));
    Sp12to4 I__3361 (
            .O(N__25174),
            .I(N__25168));
    Span4Mux_v I__3360 (
            .O(N__25171),
            .I(N__25165));
    Odrv12 I__3359 (
            .O(N__25168),
            .I(op_gt_op_gt_un13_striginternal_0));
    Odrv4 I__3358 (
            .O(N__25165),
            .I(op_gt_op_gt_un13_striginternal_0));
    InMux I__3357 (
            .O(N__25160),
            .I(N__25153));
    InMux I__3356 (
            .O(N__25159),
            .I(N__25153));
    InMux I__3355 (
            .O(N__25158),
            .I(N__25149));
    LocalMux I__3354 (
            .O(N__25153),
            .I(N__25146));
    InMux I__3353 (
            .O(N__25152),
            .I(N__25143));
    LocalMux I__3352 (
            .O(N__25149),
            .I(N__25138));
    Span4Mux_v I__3351 (
            .O(N__25146),
            .I(N__25138));
    LocalMux I__3350 (
            .O(N__25143),
            .I(un4_speriod_cry_23_THRU_CO));
    Odrv4 I__3349 (
            .O(N__25138),
            .I(un4_speriod_cry_23_THRU_CO));
    InMux I__3348 (
            .O(N__25133),
            .I(bfn_11_10_0_));
    InMux I__3347 (
            .O(N__25130),
            .I(sCounter_cry_0));
    InMux I__3346 (
            .O(N__25127),
            .I(sCounter_cry_1));
    InMux I__3345 (
            .O(N__25124),
            .I(sCounter_cry_2));
    InMux I__3344 (
            .O(N__25121),
            .I(sCounter_cry_3));
    InMux I__3343 (
            .O(N__25118),
            .I(sCounter_cry_4));
    InMux I__3342 (
            .O(N__25115),
            .I(sCounter_cry_5));
    InMux I__3341 (
            .O(N__25112),
            .I(sCounter_cry_6));
    InMux I__3340 (
            .O(N__25109),
            .I(N__25106));
    LocalMux I__3339 (
            .O(N__25106),
            .I(sEEPeriodZ0Z_19));
    InMux I__3338 (
            .O(N__25103),
            .I(N__25100));
    LocalMux I__3337 (
            .O(N__25100),
            .I(sEEPeriod_i_19));
    InMux I__3336 (
            .O(N__25097),
            .I(N__25094));
    LocalMux I__3335 (
            .O(N__25094),
            .I(sEEPeriodZ0Z_20));
    InMux I__3334 (
            .O(N__25091),
            .I(N__25088));
    LocalMux I__3333 (
            .O(N__25088),
            .I(sEEPeriod_i_20));
    InMux I__3332 (
            .O(N__25085),
            .I(N__25082));
    LocalMux I__3331 (
            .O(N__25082),
            .I(sEEPeriodZ0Z_21));
    InMux I__3330 (
            .O(N__25079),
            .I(N__25076));
    LocalMux I__3329 (
            .O(N__25076),
            .I(sEEPeriod_i_21));
    InMux I__3328 (
            .O(N__25073),
            .I(N__25070));
    LocalMux I__3327 (
            .O(N__25070),
            .I(sEEPeriodZ0Z_22));
    InMux I__3326 (
            .O(N__25067),
            .I(N__25064));
    LocalMux I__3325 (
            .O(N__25064),
            .I(sEEPeriod_i_22));
    InMux I__3324 (
            .O(N__25061),
            .I(N__25058));
    LocalMux I__3323 (
            .O(N__25058),
            .I(sEEPeriodZ0Z_23));
    InMux I__3322 (
            .O(N__25055),
            .I(N__25052));
    LocalMux I__3321 (
            .O(N__25052),
            .I(sEEPeriod_i_23));
    InMux I__3320 (
            .O(N__25049),
            .I(bfn_11_9_0_));
    CascadeMux I__3319 (
            .O(N__25046),
            .I(N__25043));
    InMux I__3318 (
            .O(N__25043),
            .I(N__25040));
    LocalMux I__3317 (
            .O(N__25040),
            .I(N__25037));
    Span4Mux_h I__3316 (
            .O(N__25037),
            .I(N__25034));
    Odrv4 I__3315 (
            .O(N__25034),
            .I(un1_spointer11_2_0_0_a2_6));
    InMux I__3314 (
            .O(N__25031),
            .I(N__25028));
    LocalMux I__3313 (
            .O(N__25028),
            .I(un1_spointer11_2_0_0_a2_1));
    InMux I__3312 (
            .O(N__25025),
            .I(N__25022));
    LocalMux I__3311 (
            .O(N__25022),
            .I(sEEPeriodZ0Z_11));
    InMux I__3310 (
            .O(N__25019),
            .I(N__25016));
    LocalMux I__3309 (
            .O(N__25016),
            .I(sEEPeriod_i_11));
    InMux I__3308 (
            .O(N__25013),
            .I(N__25010));
    LocalMux I__3307 (
            .O(N__25010),
            .I(sEEPeriodZ0Z_12));
    InMux I__3306 (
            .O(N__25007),
            .I(N__25004));
    LocalMux I__3305 (
            .O(N__25004),
            .I(sEEPeriod_i_12));
    InMux I__3304 (
            .O(N__25001),
            .I(N__24998));
    LocalMux I__3303 (
            .O(N__24998),
            .I(sEEPeriodZ0Z_13));
    InMux I__3302 (
            .O(N__24995),
            .I(N__24992));
    LocalMux I__3301 (
            .O(N__24992),
            .I(sEEPeriod_i_13));
    InMux I__3300 (
            .O(N__24989),
            .I(N__24986));
    LocalMux I__3299 (
            .O(N__24986),
            .I(sEEPeriodZ0Z_14));
    InMux I__3298 (
            .O(N__24983),
            .I(N__24980));
    LocalMux I__3297 (
            .O(N__24980),
            .I(sEEPeriod_i_14));
    InMux I__3296 (
            .O(N__24977),
            .I(N__24974));
    LocalMux I__3295 (
            .O(N__24974),
            .I(sEEPeriodZ0Z_15));
    InMux I__3294 (
            .O(N__24971),
            .I(N__24968));
    LocalMux I__3293 (
            .O(N__24968),
            .I(sEEPeriod_i_15));
    InMux I__3292 (
            .O(N__24965),
            .I(N__24962));
    LocalMux I__3291 (
            .O(N__24962),
            .I(sEEPeriodZ0Z_16));
    InMux I__3290 (
            .O(N__24959),
            .I(N__24956));
    LocalMux I__3289 (
            .O(N__24956),
            .I(sEEPeriod_i_16));
    InMux I__3288 (
            .O(N__24953),
            .I(N__24950));
    LocalMux I__3287 (
            .O(N__24950),
            .I(sEEPeriodZ0Z_17));
    InMux I__3286 (
            .O(N__24947),
            .I(N__24944));
    LocalMux I__3285 (
            .O(N__24944),
            .I(sEEPeriod_i_17));
    InMux I__3284 (
            .O(N__24941),
            .I(N__24938));
    LocalMux I__3283 (
            .O(N__24938),
            .I(sEEPeriodZ0Z_18));
    InMux I__3282 (
            .O(N__24935),
            .I(N__24932));
    LocalMux I__3281 (
            .O(N__24932),
            .I(sEEPeriod_i_18));
    InMux I__3280 (
            .O(N__24929),
            .I(N__24926));
    LocalMux I__3279 (
            .O(N__24926),
            .I(sEEPeriod_i_3));
    InMux I__3278 (
            .O(N__24923),
            .I(N__24920));
    LocalMux I__3277 (
            .O(N__24920),
            .I(sEEPeriodZ0Z_4));
    InMux I__3276 (
            .O(N__24917),
            .I(N__24914));
    LocalMux I__3275 (
            .O(N__24914),
            .I(sEEPeriod_i_4));
    InMux I__3274 (
            .O(N__24911),
            .I(N__24908));
    LocalMux I__3273 (
            .O(N__24908),
            .I(sEEPeriodZ0Z_5));
    InMux I__3272 (
            .O(N__24905),
            .I(N__24902));
    LocalMux I__3271 (
            .O(N__24902),
            .I(sEEPeriod_i_5));
    InMux I__3270 (
            .O(N__24899),
            .I(N__24896));
    LocalMux I__3269 (
            .O(N__24896),
            .I(sEEPeriodZ0Z_6));
    InMux I__3268 (
            .O(N__24893),
            .I(N__24890));
    LocalMux I__3267 (
            .O(N__24890),
            .I(sEEPeriod_i_6));
    InMux I__3266 (
            .O(N__24887),
            .I(N__24884));
    LocalMux I__3265 (
            .O(N__24884),
            .I(sEEPeriodZ0Z_7));
    CascadeMux I__3264 (
            .O(N__24881),
            .I(N__24878));
    InMux I__3263 (
            .O(N__24878),
            .I(N__24875));
    LocalMux I__3262 (
            .O(N__24875),
            .I(sEEPeriod_i_7));
    InMux I__3261 (
            .O(N__24872),
            .I(N__24869));
    LocalMux I__3260 (
            .O(N__24869),
            .I(sEEPeriodZ0Z_8));
    InMux I__3259 (
            .O(N__24866),
            .I(N__24863));
    LocalMux I__3258 (
            .O(N__24863),
            .I(sEEPeriod_i_8));
    InMux I__3257 (
            .O(N__24860),
            .I(N__24857));
    LocalMux I__3256 (
            .O(N__24857),
            .I(sEEPeriodZ0Z_9));
    InMux I__3255 (
            .O(N__24854),
            .I(N__24851));
    LocalMux I__3254 (
            .O(N__24851),
            .I(sEEPeriod_i_9));
    InMux I__3253 (
            .O(N__24848),
            .I(N__24845));
    LocalMux I__3252 (
            .O(N__24845),
            .I(sEEPeriodZ0Z_10));
    InMux I__3251 (
            .O(N__24842),
            .I(N__24839));
    LocalMux I__3250 (
            .O(N__24839),
            .I(sEEPeriod_i_10));
    CEMux I__3249 (
            .O(N__24836),
            .I(N__24833));
    LocalMux I__3248 (
            .O(N__24833),
            .I(N__24830));
    Span4Mux_v I__3247 (
            .O(N__24830),
            .I(N__24827));
    Odrv4 I__3246 (
            .O(N__24827),
            .I(sAddress_RNIETI62Z0Z_1));
    InMux I__3245 (
            .O(N__24824),
            .I(N__24821));
    LocalMux I__3244 (
            .O(N__24821),
            .I(sEEPeriodZ0Z_0));
    InMux I__3243 (
            .O(N__24818),
            .I(N__24815));
    LocalMux I__3242 (
            .O(N__24815),
            .I(sEEPeriod_i_0));
    InMux I__3241 (
            .O(N__24812),
            .I(N__24809));
    LocalMux I__3240 (
            .O(N__24809),
            .I(sEEPeriodZ0Z_1));
    InMux I__3239 (
            .O(N__24806),
            .I(N__24803));
    LocalMux I__3238 (
            .O(N__24803),
            .I(sEEPeriod_i_1));
    InMux I__3237 (
            .O(N__24800),
            .I(N__24797));
    LocalMux I__3236 (
            .O(N__24797),
            .I(sEEPeriodZ0Z_2));
    InMux I__3235 (
            .O(N__24794),
            .I(N__24791));
    LocalMux I__3234 (
            .O(N__24791),
            .I(sEEPeriod_i_2));
    InMux I__3233 (
            .O(N__24788),
            .I(N__24785));
    LocalMux I__3232 (
            .O(N__24785),
            .I(sEEPeriodZ0Z_3));
    InMux I__3231 (
            .O(N__24782),
            .I(N__24779));
    LocalMux I__3230 (
            .O(N__24779),
            .I(sDAC_dataZ0Z_0));
    InMux I__3229 (
            .O(N__24776),
            .I(N__24773));
    LocalMux I__3228 (
            .O(N__24773),
            .I(sDAC_dataZ0Z_1));
    InMux I__3227 (
            .O(N__24770),
            .I(N__24767));
    LocalMux I__3226 (
            .O(N__24767),
            .I(sDAC_dataZ0Z_11));
    InMux I__3225 (
            .O(N__24764),
            .I(N__24761));
    LocalMux I__3224 (
            .O(N__24761),
            .I(sDAC_dataZ0Z_12));
    InMux I__3223 (
            .O(N__24758),
            .I(N__24755));
    LocalMux I__3222 (
            .O(N__24755),
            .I(sDAC_dataZ0Z_13));
    InMux I__3221 (
            .O(N__24752),
            .I(N__24749));
    LocalMux I__3220 (
            .O(N__24749),
            .I(sDAC_dataZ0Z_14));
    InMux I__3219 (
            .O(N__24746),
            .I(N__24743));
    LocalMux I__3218 (
            .O(N__24743),
            .I(sDAC_dataZ0Z_15));
    CEMux I__3217 (
            .O(N__24740),
            .I(N__24737));
    LocalMux I__3216 (
            .O(N__24737),
            .I(N__24734));
    Span4Mux_v I__3215 (
            .O(N__24734),
            .I(N__24731));
    Span4Mux_v I__3214 (
            .O(N__24731),
            .I(N__24728));
    Odrv4 I__3213 (
            .O(N__24728),
            .I(sAddress_RNIA6242Z0Z_0));
    IoInMux I__3212 (
            .O(N__24725),
            .I(N__24722));
    LocalMux I__3211 (
            .O(N__24722),
            .I(N__24719));
    Span4Mux_s3_v I__3210 (
            .O(N__24719),
            .I(N__24716));
    Span4Mux_v I__3209 (
            .O(N__24716),
            .I(N__24713));
    Odrv4 I__3208 (
            .O(N__24713),
            .I(LED3_c_i));
    InMux I__3207 (
            .O(N__24710),
            .I(N__24707));
    LocalMux I__3206 (
            .O(N__24707),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15 ));
    InMux I__3205 (
            .O(N__24704),
            .I(N__24701));
    LocalMux I__3204 (
            .O(N__24701),
            .I(N__24697));
    InMux I__3203 (
            .O(N__24700),
            .I(N__24694));
    Span4Mux_h I__3202 (
            .O(N__24697),
            .I(N__24686));
    LocalMux I__3201 (
            .O(N__24694),
            .I(N__24686));
    InMux I__3200 (
            .O(N__24693),
            .I(N__24683));
    InMux I__3199 (
            .O(N__24692),
            .I(N__24677));
    InMux I__3198 (
            .O(N__24691),
            .I(N__24677));
    Span4Mux_h I__3197 (
            .O(N__24686),
            .I(N__24672));
    LocalMux I__3196 (
            .O(N__24683),
            .I(N__24672));
    InMux I__3195 (
            .O(N__24682),
            .I(N__24669));
    LocalMux I__3194 (
            .O(N__24677),
            .I(N__24664));
    Span4Mux_h I__3193 (
            .O(N__24672),
            .I(N__24659));
    LocalMux I__3192 (
            .O(N__24669),
            .I(N__24659));
    InMux I__3191 (
            .O(N__24668),
            .I(N__24656));
    InMux I__3190 (
            .O(N__24667),
            .I(N__24653));
    Span4Mux_h I__3189 (
            .O(N__24664),
            .I(N__24646));
    Span4Mux_v I__3188 (
            .O(N__24659),
            .I(N__24643));
    LocalMux I__3187 (
            .O(N__24656),
            .I(N__24638));
    LocalMux I__3186 (
            .O(N__24653),
            .I(N__24638));
    InMux I__3185 (
            .O(N__24652),
            .I(N__24633));
    InMux I__3184 (
            .O(N__24651),
            .I(N__24633));
    InMux I__3183 (
            .O(N__24650),
            .I(N__24630));
    InMux I__3182 (
            .O(N__24649),
            .I(N__24627));
    Odrv4 I__3181 (
            .O(N__24646),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ));
    Odrv4 I__3180 (
            .O(N__24643),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ));
    Odrv12 I__3179 (
            .O(N__24638),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ));
    LocalMux I__3178 (
            .O(N__24633),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ));
    LocalMux I__3177 (
            .O(N__24630),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ));
    LocalMux I__3176 (
            .O(N__24627),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ));
    InMux I__3175 (
            .O(N__24614),
            .I(N__24611));
    LocalMux I__3174 (
            .O(N__24611),
            .I(N__24608));
    Odrv12 I__3173 (
            .O(N__24608),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15 ));
    CEMux I__3172 (
            .O(N__24605),
            .I(N__24602));
    LocalMux I__3171 (
            .O(N__24602),
            .I(N__24599));
    Span4Mux_v I__3170 (
            .O(N__24599),
            .I(N__24596));
    Odrv4 I__3169 (
            .O(N__24596),
            .I(sAddress_RNIA6242_4Z0Z_0));
    CEMux I__3168 (
            .O(N__24593),
            .I(N__24590));
    LocalMux I__3167 (
            .O(N__24590),
            .I(N__24587));
    Span4Mux_v I__3166 (
            .O(N__24587),
            .I(N__24584));
    Span4Mux_h I__3165 (
            .O(N__24584),
            .I(N__24581));
    Odrv4 I__3164 (
            .O(N__24581),
            .I(sDAC_mem_31_1_sqmuxa));
    CascadeMux I__3163 (
            .O(N__24578),
            .I(\spi_slave_inst.un23_i_ssn_cascade_ ));
    InMux I__3162 (
            .O(N__24575),
            .I(N__24572));
    LocalMux I__3161 (
            .O(N__24572),
            .I(N__24569));
    Odrv4 I__3160 (
            .O(N__24569),
            .I(g0_10));
    InMux I__3159 (
            .O(N__24566),
            .I(N__24563));
    LocalMux I__3158 (
            .O(N__24563),
            .I(g0_10_0));
    CascadeMux I__3157 (
            .O(N__24560),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2_cascade_ ));
    InMux I__3156 (
            .O(N__24557),
            .I(N__24554));
    LocalMux I__3155 (
            .O(N__24554),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2 ));
    InMux I__3154 (
            .O(N__24551),
            .I(N__24547));
    InMux I__3153 (
            .O(N__24550),
            .I(N__24544));
    LocalMux I__3152 (
            .O(N__24547),
            .I(N__24538));
    LocalMux I__3151 (
            .O(N__24544),
            .I(N__24538));
    InMux I__3150 (
            .O(N__24543),
            .I(N__24535));
    Span4Mux_v I__3149 (
            .O(N__24538),
            .I(N__24530));
    LocalMux I__3148 (
            .O(N__24535),
            .I(N__24530));
    Span4Mux_h I__3147 (
            .O(N__24530),
            .I(N__24527));
    Span4Mux_h I__3146 (
            .O(N__24527),
            .I(N__24524));
    Odrv4 I__3145 (
            .O(N__24524),
            .I(\spi_master_inst.sclk_gen_u0.N_158_7 ));
    CascadeMux I__3144 (
            .O(N__24521),
            .I(N__24517));
    InMux I__3143 (
            .O(N__24520),
            .I(N__24514));
    InMux I__3142 (
            .O(N__24517),
            .I(N__24509));
    LocalMux I__3141 (
            .O(N__24514),
            .I(N__24506));
    CascadeMux I__3140 (
            .O(N__24513),
            .I(N__24503));
    CascadeMux I__3139 (
            .O(N__24512),
            .I(N__24500));
    LocalMux I__3138 (
            .O(N__24509),
            .I(N__24496));
    Span4Mux_v I__3137 (
            .O(N__24506),
            .I(N__24492));
    InMux I__3136 (
            .O(N__24503),
            .I(N__24489));
    InMux I__3135 (
            .O(N__24500),
            .I(N__24486));
    InMux I__3134 (
            .O(N__24499),
            .I(N__24483));
    Span4Mux_h I__3133 (
            .O(N__24496),
            .I(N__24480));
    InMux I__3132 (
            .O(N__24495),
            .I(N__24477));
    Span4Mux_h I__3131 (
            .O(N__24492),
            .I(N__24474));
    LocalMux I__3130 (
            .O(N__24489),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ));
    LocalMux I__3129 (
            .O(N__24486),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ));
    LocalMux I__3128 (
            .O(N__24483),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ));
    Odrv4 I__3127 (
            .O(N__24480),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ));
    LocalMux I__3126 (
            .O(N__24477),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ));
    Odrv4 I__3125 (
            .O(N__24474),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ));
    InMux I__3124 (
            .O(N__24461),
            .I(N__24456));
    InMux I__3123 (
            .O(N__24460),
            .I(N__24451));
    InMux I__3122 (
            .O(N__24459),
            .I(N__24448));
    LocalMux I__3121 (
            .O(N__24456),
            .I(N__24445));
    InMux I__3120 (
            .O(N__24455),
            .I(N__24442));
    InMux I__3119 (
            .O(N__24454),
            .I(N__24439));
    LocalMux I__3118 (
            .O(N__24451),
            .I(N__24434));
    LocalMux I__3117 (
            .O(N__24448),
            .I(N__24434));
    Span4Mux_h I__3116 (
            .O(N__24445),
            .I(N__24431));
    LocalMux I__3115 (
            .O(N__24442),
            .I(N__24428));
    LocalMux I__3114 (
            .O(N__24439),
            .I(N__24425));
    Span4Mux_h I__3113 (
            .O(N__24434),
            .I(N__24422));
    Span4Mux_h I__3112 (
            .O(N__24431),
            .I(N__24419));
    Span4Mux_v I__3111 (
            .O(N__24428),
            .I(N__24416));
    Span4Mux_v I__3110 (
            .O(N__24425),
            .I(N__24413));
    Span4Mux_h I__3109 (
            .O(N__24422),
            .I(N__24410));
    Span4Mux_v I__3108 (
            .O(N__24419),
            .I(N__24407));
    Span4Mux_v I__3107 (
            .O(N__24416),
            .I(N__24404));
    Span4Mux_h I__3106 (
            .O(N__24413),
            .I(N__24399));
    Span4Mux_v I__3105 (
            .O(N__24410),
            .I(N__24399));
    Odrv4 I__3104 (
            .O(N__24407),
            .I(\spi_master_inst.sclk_gen_u0.spi_start_iZ0 ));
    Odrv4 I__3103 (
            .O(N__24404),
            .I(\spi_master_inst.sclk_gen_u0.spi_start_iZ0 ));
    Odrv4 I__3102 (
            .O(N__24399),
            .I(\spi_master_inst.sclk_gen_u0.spi_start_iZ0 ));
    CascadeMux I__3101 (
            .O(N__24392),
            .I(\spi_master_inst.sclk_gen_u0.N_158_7_cascade_ ));
    InMux I__3100 (
            .O(N__24389),
            .I(N__24382));
    InMux I__3099 (
            .O(N__24388),
            .I(N__24379));
    CascadeMux I__3098 (
            .O(N__24387),
            .I(N__24375));
    InMux I__3097 (
            .O(N__24386),
            .I(N__24372));
    InMux I__3096 (
            .O(N__24385),
            .I(N__24369));
    LocalMux I__3095 (
            .O(N__24382),
            .I(N__24366));
    LocalMux I__3094 (
            .O(N__24379),
            .I(N__24363));
    InMux I__3093 (
            .O(N__24378),
            .I(N__24360));
    InMux I__3092 (
            .O(N__24375),
            .I(N__24357));
    LocalMux I__3091 (
            .O(N__24372),
            .I(N__24354));
    LocalMux I__3090 (
            .O(N__24369),
            .I(N__24349));
    Span4Mux_v I__3089 (
            .O(N__24366),
            .I(N__24349));
    Span12Mux_h I__3088 (
            .O(N__24363),
            .I(N__24346));
    LocalMux I__3087 (
            .O(N__24360),
            .I(N__24339));
    LocalMux I__3086 (
            .O(N__24357),
            .I(N__24339));
    Span4Mux_h I__3085 (
            .O(N__24354),
            .I(N__24339));
    Odrv4 I__3084 (
            .O(N__24349),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ));
    Odrv12 I__3083 (
            .O(N__24346),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ));
    Odrv4 I__3082 (
            .O(N__24339),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ));
    InMux I__3081 (
            .O(N__24332),
            .I(N__24329));
    LocalMux I__3080 (
            .O(N__24329),
            .I(N__24326));
    Span4Mux_h I__3079 (
            .O(N__24326),
            .I(N__24323));
    Span4Mux_v I__3078 (
            .O(N__24323),
            .I(N__24320));
    Span4Mux_h I__3077 (
            .O(N__24320),
            .I(N__24317));
    Odrv4 I__3076 (
            .O(N__24317),
            .I(\spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0 ));
    InMux I__3075 (
            .O(N__24314),
            .I(N__24311));
    LocalMux I__3074 (
            .O(N__24311),
            .I(g2_6));
    InMux I__3073 (
            .O(N__24308),
            .I(N__24305));
    LocalMux I__3072 (
            .O(N__24305),
            .I(N__24301));
    InMux I__3071 (
            .O(N__24304),
            .I(N__24298));
    Span4Mux_h I__3070 (
            .O(N__24301),
            .I(N__24295));
    LocalMux I__3069 (
            .O(N__24298),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4 ));
    Odrv4 I__3068 (
            .O(N__24295),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4 ));
    InMux I__3067 (
            .O(N__24290),
            .I(N__24287));
    LocalMux I__3066 (
            .O(N__24287),
            .I(N__24283));
    InMux I__3065 (
            .O(N__24286),
            .I(N__24280));
    Span4Mux_h I__3064 (
            .O(N__24283),
            .I(N__24277));
    LocalMux I__3063 (
            .O(N__24280),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3 ));
    Odrv4 I__3062 (
            .O(N__24277),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3 ));
    InMux I__3061 (
            .O(N__24272),
            .I(N__24269));
    LocalMux I__3060 (
            .O(N__24269),
            .I(N__24266));
    Span4Mux_v I__3059 (
            .O(N__24266),
            .I(N__24263));
    Span4Mux_h I__3058 (
            .O(N__24263),
            .I(N__24260));
    Odrv4 I__3057 (
            .O(N__24260),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_i6_3 ));
    InMux I__3056 (
            .O(N__24257),
            .I(N__24251));
    InMux I__3055 (
            .O(N__24256),
            .I(N__24248));
    InMux I__3054 (
            .O(N__24255),
            .I(N__24243));
    InMux I__3053 (
            .O(N__24254),
            .I(N__24243));
    LocalMux I__3052 (
            .O(N__24251),
            .I(N__24240));
    LocalMux I__3051 (
            .O(N__24248),
            .I(N__24235));
    LocalMux I__3050 (
            .O(N__24243),
            .I(N__24235));
    Span4Mux_h I__3049 (
            .O(N__24240),
            .I(N__24232));
    Span12Mux_h I__3048 (
            .O(N__24235),
            .I(N__24227));
    Sp12to4 I__3047 (
            .O(N__24232),
            .I(N__24227));
    Odrv12 I__3046 (
            .O(N__24227),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_i6 ));
    CascadeMux I__3045 (
            .O(N__24224),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_ ));
    CascadeMux I__3044 (
            .O(N__24221),
            .I(N__24217));
    InMux I__3043 (
            .O(N__24220),
            .I(N__24214));
    InMux I__3042 (
            .O(N__24217),
            .I(N__24211));
    LocalMux I__3041 (
            .O(N__24214),
            .I(N__24206));
    LocalMux I__3040 (
            .O(N__24211),
            .I(N__24206));
    Span4Mux_h I__3039 (
            .O(N__24206),
            .I(N__24203));
    Odrv4 I__3038 (
            .O(N__24203),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_3 ));
    CascadeMux I__3037 (
            .O(N__24200),
            .I(\spi_slave_inst.un23_i_ssn_3_cascade_ ));
    InMux I__3036 (
            .O(N__24197),
            .I(N__24194));
    LocalMux I__3035 (
            .O(N__24194),
            .I(N__24191));
    Span4Mux_v I__3034 (
            .O(N__24191),
            .I(N__24188));
    Odrv4 I__3033 (
            .O(N__24188),
            .I(un21_trig_prev_21_5));
    CascadeMux I__3032 (
            .O(N__24185),
            .I(op_gt_op_gt_un13_striginternallto23_5_cascade_));
    InMux I__3031 (
            .O(N__24182),
            .I(N__24179));
    LocalMux I__3030 (
            .O(N__24179),
            .I(N__24176));
    Odrv12 I__3029 (
            .O(N__24176),
            .I(un1_reset_rpi_inv_2_0_o2_2));
    InMux I__3028 (
            .O(N__24173),
            .I(N__24170));
    LocalMux I__3027 (
            .O(N__24170),
            .I(g0_13_0));
    InMux I__3026 (
            .O(N__24167),
            .I(N__24164));
    LocalMux I__3025 (
            .O(N__24164),
            .I(un21_trig_prev_21_4));
    InMux I__3024 (
            .O(N__24161),
            .I(N__24158));
    LocalMux I__3023 (
            .O(N__24158),
            .I(g0_6));
    CascadeMux I__3022 (
            .O(N__24155),
            .I(N__24152));
    InMux I__3021 (
            .O(N__24152),
            .I(N__24149));
    LocalMux I__3020 (
            .O(N__24149),
            .I(N__24146));
    Odrv4 I__3019 (
            .O(N__24146),
            .I(N_99));
    InMux I__3018 (
            .O(N__24143),
            .I(N__24140));
    LocalMux I__3017 (
            .O(N__24140),
            .I(op_gt_op_gt_un13_striginternallto23_3));
    CascadeMux I__3016 (
            .O(N__24137),
            .I(N__24133));
    InMux I__3015 (
            .O(N__24136),
            .I(N__24130));
    InMux I__3014 (
            .O(N__24133),
            .I(N__24127));
    LocalMux I__3013 (
            .O(N__24130),
            .I(N__24124));
    LocalMux I__3012 (
            .O(N__24127),
            .I(N_831_16));
    Odrv4 I__3011 (
            .O(N__24124),
            .I(N_831_16));
    InMux I__3010 (
            .O(N__24119),
            .I(N__24116));
    LocalMux I__3009 (
            .O(N__24116),
            .I(op_gt_op_gt_un13_striginternallto23_6));
    CEMux I__3008 (
            .O(N__24113),
            .I(N__24110));
    LocalMux I__3007 (
            .O(N__24110),
            .I(sDAC_mem_15_1_sqmuxa));
    CEMux I__3006 (
            .O(N__24107),
            .I(N__24104));
    LocalMux I__3005 (
            .O(N__24104),
            .I(N__24101));
    Span4Mux_v I__3004 (
            .O(N__24101),
            .I(N__24098));
    Span4Mux_h I__3003 (
            .O(N__24098),
            .I(N__24095));
    Odrv4 I__3002 (
            .O(N__24095),
            .I(sAddress_RNI9IH12_1Z0Z_2));
    CEMux I__3001 (
            .O(N__24092),
            .I(N__24089));
    LocalMux I__3000 (
            .O(N__24089),
            .I(N__24086));
    Span4Mux_v I__2999 (
            .O(N__24086),
            .I(N__24083));
    Span4Mux_h I__2998 (
            .O(N__24083),
            .I(N__24080));
    Odrv4 I__2997 (
            .O(N__24080),
            .I(sDAC_mem_14_1_sqmuxa));
    CEMux I__2996 (
            .O(N__24077),
            .I(N__24074));
    LocalMux I__2995 (
            .O(N__24074),
            .I(N__24071));
    Span4Mux_h I__2994 (
            .O(N__24071),
            .I(N__24068));
    Span4Mux_h I__2993 (
            .O(N__24068),
            .I(N__24065));
    Odrv4 I__2992 (
            .O(N__24065),
            .I(sAddress_RNI9IH12Z0Z_0));
    CEMux I__2991 (
            .O(N__24062),
            .I(N__24059));
    LocalMux I__2990 (
            .O(N__24059),
            .I(N__24056));
    Odrv4 I__2989 (
            .O(N__24056),
            .I(sDAC_mem_42_1_sqmuxa));
    InMux I__2988 (
            .O(N__24053),
            .I(N__24050));
    LocalMux I__2987 (
            .O(N__24050),
            .I(N__24047));
    Span4Mux_h I__2986 (
            .O(N__24047),
            .I(N__24044));
    Odrv4 I__2985 (
            .O(N__24044),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_11 ));
    InMux I__2984 (
            .O(N__24041),
            .I(N__24038));
    LocalMux I__2983 (
            .O(N__24038),
            .I(N__24035));
    Odrv4 I__2982 (
            .O(N__24035),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_13 ));
    InMux I__2981 (
            .O(N__24032),
            .I(N__24029));
    LocalMux I__2980 (
            .O(N__24029),
            .I(N__24026));
    Odrv4 I__2979 (
            .O(N__24026),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_14 ));
    InMux I__2978 (
            .O(N__24023),
            .I(N__24020));
    LocalMux I__2977 (
            .O(N__24020),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_15 ));
    InMux I__2976 (
            .O(N__24017),
            .I(bfn_9_20_0_));
    IoInMux I__2975 (
            .O(N__24014),
            .I(N__24011));
    LocalMux I__2974 (
            .O(N__24011),
            .I(N__24008));
    Span12Mux_s0_h I__2973 (
            .O(N__24008),
            .I(N__24005));
    Span12Mux_h I__2972 (
            .O(N__24005),
            .I(N__24002));
    Odrv12 I__2971 (
            .O(N__24002),
            .I(pon_obuf_RNOZ0));
    InMux I__2970 (
            .O(N__23999),
            .I(N__23996));
    LocalMux I__2969 (
            .O(N__23996),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10 ));
    InMux I__2968 (
            .O(N__23993),
            .I(N__23990));
    LocalMux I__2967 (
            .O(N__23990),
            .I(N__23987));
    Odrv12 I__2966 (
            .O(N__23987),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_0 ));
    InMux I__2965 (
            .O(N__23984),
            .I(N__23981));
    LocalMux I__2964 (
            .O(N__23981),
            .I(N__23978));
    Odrv12 I__2963 (
            .O(N__23978),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_1 ));
    InMux I__2962 (
            .O(N__23975),
            .I(N__23972));
    LocalMux I__2961 (
            .O(N__23972),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_10 ));
    InMux I__2960 (
            .O(N__23969),
            .I(N__23966));
    LocalMux I__2959 (
            .O(N__23966),
            .I(sEEPonZ0Z_4));
    InMux I__2958 (
            .O(N__23963),
            .I(N__23960));
    LocalMux I__2957 (
            .O(N__23960),
            .I(sEEPon_i_4));
    InMux I__2956 (
            .O(N__23957),
            .I(N__23954));
    LocalMux I__2955 (
            .O(N__23954),
            .I(sEEPonZ0Z_5));
    InMux I__2954 (
            .O(N__23951),
            .I(N__23948));
    LocalMux I__2953 (
            .O(N__23948),
            .I(sEEPon_i_5));
    InMux I__2952 (
            .O(N__23945),
            .I(N__23942));
    LocalMux I__2951 (
            .O(N__23942),
            .I(sEEPonZ0Z_6));
    InMux I__2950 (
            .O(N__23939),
            .I(N__23936));
    LocalMux I__2949 (
            .O(N__23936),
            .I(sEEPon_i_6));
    InMux I__2948 (
            .O(N__23933),
            .I(N__23930));
    LocalMux I__2947 (
            .O(N__23930),
            .I(sEEPonZ0Z_7));
    InMux I__2946 (
            .O(N__23927),
            .I(N__23924));
    LocalMux I__2945 (
            .O(N__23924),
            .I(sEEPon_i_7));
    CEMux I__2944 (
            .O(N__23921),
            .I(N__23918));
    LocalMux I__2943 (
            .O(N__23918),
            .I(N__23915));
    Sp12to4 I__2942 (
            .O(N__23915),
            .I(N__23912));
    Odrv12 I__2941 (
            .O(N__23912),
            .I(sDAC_mem_30_1_sqmuxa));
    InMux I__2940 (
            .O(N__23909),
            .I(N__23906));
    LocalMux I__2939 (
            .O(N__23906),
            .I(sEEPonZ0Z_0));
    CascadeMux I__2938 (
            .O(N__23903),
            .I(N__23900));
    InMux I__2937 (
            .O(N__23900),
            .I(N__23897));
    LocalMux I__2936 (
            .O(N__23897),
            .I(sEEPon_i_0));
    InMux I__2935 (
            .O(N__23894),
            .I(N__23891));
    LocalMux I__2934 (
            .O(N__23891),
            .I(sEEPonZ0Z_1));
    InMux I__2933 (
            .O(N__23888),
            .I(N__23885));
    LocalMux I__2932 (
            .O(N__23885),
            .I(sEEPon_i_1));
    InMux I__2931 (
            .O(N__23882),
            .I(N__23879));
    LocalMux I__2930 (
            .O(N__23879),
            .I(sEEPonZ0Z_2));
    InMux I__2929 (
            .O(N__23876),
            .I(N__23873));
    LocalMux I__2928 (
            .O(N__23873),
            .I(sEEPon_i_2));
    InMux I__2927 (
            .O(N__23870),
            .I(N__23867));
    LocalMux I__2926 (
            .O(N__23867),
            .I(sEEPonZ0Z_3));
    InMux I__2925 (
            .O(N__23864),
            .I(N__23861));
    LocalMux I__2924 (
            .O(N__23861),
            .I(sEEPon_i_3));
    CascadeMux I__2923 (
            .O(N__23858),
            .I(N__23855));
    InMux I__2922 (
            .O(N__23855),
            .I(N__23852));
    LocalMux I__2921 (
            .O(N__23852),
            .I(g0_13_1));
    CascadeMux I__2920 (
            .O(N__23849),
            .I(N__23846));
    InMux I__2919 (
            .O(N__23846),
            .I(N__23843));
    LocalMux I__2918 (
            .O(N__23843),
            .I(g0_17_0));
    InMux I__2917 (
            .O(N__23840),
            .I(N__23837));
    LocalMux I__2916 (
            .O(N__23837),
            .I(N__23831));
    InMux I__2915 (
            .O(N__23836),
            .I(N__23828));
    CascadeMux I__2914 (
            .O(N__23835),
            .I(N__23825));
    CascadeMux I__2913 (
            .O(N__23834),
            .I(N__23820));
    Span4Mux_v I__2912 (
            .O(N__23831),
            .I(N__23817));
    LocalMux I__2911 (
            .O(N__23828),
            .I(N__23814));
    InMux I__2910 (
            .O(N__23825),
            .I(N__23805));
    InMux I__2909 (
            .O(N__23824),
            .I(N__23805));
    InMux I__2908 (
            .O(N__23823),
            .I(N__23805));
    InMux I__2907 (
            .O(N__23820),
            .I(N__23805));
    Odrv4 I__2906 (
            .O(N__23817),
            .I(N_326));
    Odrv12 I__2905 (
            .O(N__23814),
            .I(N_326));
    LocalMux I__2904 (
            .O(N__23805),
            .I(N_326));
    InMux I__2903 (
            .O(N__23798),
            .I(N__23795));
    LocalMux I__2902 (
            .O(N__23795),
            .I(g0_16_0));
    InMux I__2901 (
            .O(N__23792),
            .I(N__23789));
    LocalMux I__2900 (
            .O(N__23789),
            .I(g1_i_a4_6));
    CascadeMux I__2899 (
            .O(N__23786),
            .I(g1_i_a4_5_cascade_));
    InMux I__2898 (
            .O(N__23783),
            .I(N__23780));
    LocalMux I__2897 (
            .O(N__23780),
            .I(N__23777));
    Odrv4 I__2896 (
            .O(N__23777),
            .I(un1_reset_rpi_inv_2_0_o2_5));
    CascadeMux I__2895 (
            .O(N__23774),
            .I(g1_i_a4_9_cascade_));
    InMux I__2894 (
            .O(N__23771),
            .I(N__23768));
    LocalMux I__2893 (
            .O(N__23768),
            .I(N__23765));
    Odrv4 I__2892 (
            .O(N__23765),
            .I(sEETrigInternal_prev_RNIH3OJZ0Z1));
    CascadeMux I__2891 (
            .O(N__23762),
            .I(N__23759));
    InMux I__2890 (
            .O(N__23759),
            .I(N__23756));
    LocalMux I__2889 (
            .O(N__23756),
            .I(N__23753));
    Span4Mux_h I__2888 (
            .O(N__23753),
            .I(N__23750));
    Odrv4 I__2887 (
            .O(N__23750),
            .I(g0_0_1));
    InMux I__2886 (
            .O(N__23747),
            .I(N__23744));
    LocalMux I__2885 (
            .O(N__23744),
            .I(g0_16));
    CascadeMux I__2884 (
            .O(N__23741),
            .I(N__23738));
    InMux I__2883 (
            .O(N__23738),
            .I(N__23735));
    LocalMux I__2882 (
            .O(N__23735),
            .I(N__23732));
    Span4Mux_v I__2881 (
            .O(N__23732),
            .I(N__23729));
    Odrv4 I__2880 (
            .O(N__23729),
            .I(g0_11));
    InMux I__2879 (
            .O(N__23726),
            .I(N__23723));
    LocalMux I__2878 (
            .O(N__23723),
            .I(g0_14));
    InMux I__2877 (
            .O(N__23720),
            .I(N__23715));
    InMux I__2876 (
            .O(N__23719),
            .I(N__23712));
    InMux I__2875 (
            .O(N__23718),
            .I(N__23708));
    LocalMux I__2874 (
            .O(N__23715),
            .I(N__23699));
    LocalMux I__2873 (
            .O(N__23712),
            .I(N__23699));
    InMux I__2872 (
            .O(N__23711),
            .I(N__23696));
    LocalMux I__2871 (
            .O(N__23708),
            .I(N__23693));
    InMux I__2870 (
            .O(N__23707),
            .I(N__23688));
    InMux I__2869 (
            .O(N__23706),
            .I(N__23688));
    InMux I__2868 (
            .O(N__23705),
            .I(N__23683));
    InMux I__2867 (
            .O(N__23704),
            .I(N__23683));
    Sp12to4 I__2866 (
            .O(N__23699),
            .I(N__23678));
    LocalMux I__2865 (
            .O(N__23696),
            .I(N__23678));
    Span4Mux_v I__2864 (
            .O(N__23693),
            .I(N__23675));
    LocalMux I__2863 (
            .O(N__23688),
            .I(sEETrigInternalZ0));
    LocalMux I__2862 (
            .O(N__23683),
            .I(sEETrigInternalZ0));
    Odrv12 I__2861 (
            .O(N__23678),
            .I(sEETrigInternalZ0));
    Odrv4 I__2860 (
            .O(N__23675),
            .I(sEETrigInternalZ0));
    InMux I__2859 (
            .O(N__23666),
            .I(N__23663));
    LocalMux I__2858 (
            .O(N__23663),
            .I(N__23660));
    Odrv4 I__2857 (
            .O(N__23660),
            .I(g3_0));
    CascadeMux I__2856 (
            .O(N__23657),
            .I(N__23652));
    InMux I__2855 (
            .O(N__23656),
            .I(N__23649));
    InMux I__2854 (
            .O(N__23655),
            .I(N__23646));
    InMux I__2853 (
            .O(N__23652),
            .I(N__23642));
    LocalMux I__2852 (
            .O(N__23649),
            .I(N__23637));
    LocalMux I__2851 (
            .O(N__23646),
            .I(N__23637));
    InMux I__2850 (
            .O(N__23645),
            .I(N__23634));
    LocalMux I__2849 (
            .O(N__23642),
            .I(N__23631));
    Sp12to4 I__2848 (
            .O(N__23637),
            .I(N__23628));
    LocalMux I__2847 (
            .O(N__23634),
            .I(N__23623));
    Span4Mux_h I__2846 (
            .O(N__23631),
            .I(N__23623));
    Odrv12 I__2845 (
            .O(N__23628),
            .I(sEETrigInternal_prevZ0));
    Odrv4 I__2844 (
            .O(N__23623),
            .I(sEETrigInternal_prevZ0));
    IoInMux I__2843 (
            .O(N__23618),
            .I(N__23615));
    LocalMux I__2842 (
            .O(N__23615),
            .I(N__23612));
    Span4Mux_s1_h I__2841 (
            .O(N__23612),
            .I(N__23609));
    Span4Mux_h I__2840 (
            .O(N__23609),
            .I(N__23603));
    InMux I__2839 (
            .O(N__23608),
            .I(N__23598));
    InMux I__2838 (
            .O(N__23607),
            .I(N__23598));
    InMux I__2837 (
            .O(N__23606),
            .I(N__23595));
    Sp12to4 I__2836 (
            .O(N__23603),
            .I(N__23592));
    LocalMux I__2835 (
            .O(N__23598),
            .I(N__23589));
    LocalMux I__2834 (
            .O(N__23595),
            .I(N__23586));
    Span12Mux_v I__2833 (
            .O(N__23592),
            .I(N__23583));
    Span4Mux_h I__2832 (
            .O(N__23589),
            .I(N__23580));
    Span4Mux_h I__2831 (
            .O(N__23586),
            .I(N__23577));
    Odrv12 I__2830 (
            .O(N__23583),
            .I(LED_MODE_c));
    Odrv4 I__2829 (
            .O(N__23580),
            .I(LED_MODE_c));
    Odrv4 I__2828 (
            .O(N__23577),
            .I(LED_MODE_c));
    CascadeMux I__2827 (
            .O(N__23570),
            .I(N_831_16_cascade_));
    InMux I__2826 (
            .O(N__23567),
            .I(N__23562));
    CascadeMux I__2825 (
            .O(N__23566),
            .I(N__23558));
    CascadeMux I__2824 (
            .O(N__23565),
            .I(N__23555));
    LocalMux I__2823 (
            .O(N__23562),
            .I(N__23551));
    InMux I__2822 (
            .O(N__23561),
            .I(N__23547));
    InMux I__2821 (
            .O(N__23558),
            .I(N__23542));
    InMux I__2820 (
            .O(N__23555),
            .I(N__23542));
    InMux I__2819 (
            .O(N__23554),
            .I(N__23539));
    Span4Mux_h I__2818 (
            .O(N__23551),
            .I(N__23536));
    InMux I__2817 (
            .O(N__23550),
            .I(N__23533));
    LocalMux I__2816 (
            .O(N__23547),
            .I(N__23528));
    LocalMux I__2815 (
            .O(N__23542),
            .I(N__23528));
    LocalMux I__2814 (
            .O(N__23539),
            .I(N_319));
    Odrv4 I__2813 (
            .O(N__23536),
            .I(N_319));
    LocalMux I__2812 (
            .O(N__23533),
            .I(N_319));
    Odrv4 I__2811 (
            .O(N__23528),
            .I(N_319));
    CascadeMux I__2810 (
            .O(N__23519),
            .I(g0_13_cascade_));
    CascadeMux I__2809 (
            .O(N__23516),
            .I(N__23513));
    InMux I__2808 (
            .O(N__23513),
            .I(N__23510));
    LocalMux I__2807 (
            .O(N__23510),
            .I(g0_1_0));
    InMux I__2806 (
            .O(N__23507),
            .I(N__23504));
    LocalMux I__2805 (
            .O(N__23504),
            .I(g0_15_0));
    CascadeMux I__2804 (
            .O(N__23501),
            .I(sAddress_RNIAM2A_0Z0Z_1_cascade_));
    CascadeMux I__2803 (
            .O(N__23498),
            .I(N_445_cascade_));
    CascadeMux I__2802 (
            .O(N__23495),
            .I(N__23491));
    InMux I__2801 (
            .O(N__23494),
            .I(N__23485));
    InMux I__2800 (
            .O(N__23491),
            .I(N__23485));
    InMux I__2799 (
            .O(N__23490),
            .I(N__23482));
    LocalMux I__2798 (
            .O(N__23485),
            .I(N__23479));
    LocalMux I__2797 (
            .O(N__23482),
            .I(sAddress_RNI6VH7_5Z0Z_1));
    Odrv4 I__2796 (
            .O(N__23479),
            .I(sAddress_RNI6VH7_5Z0Z_1));
    InMux I__2795 (
            .O(N__23474),
            .I(N__23471));
    LocalMux I__2794 (
            .O(N__23471),
            .I(N_445));
    CascadeMux I__2793 (
            .O(N__23468),
            .I(N__23465));
    InMux I__2792 (
            .O(N__23465),
            .I(N__23458));
    InMux I__2791 (
            .O(N__23464),
            .I(N__23455));
    InMux I__2790 (
            .O(N__23463),
            .I(N__23452));
    InMux I__2789 (
            .O(N__23462),
            .I(N__23449));
    InMux I__2788 (
            .O(N__23461),
            .I(N__23446));
    LocalMux I__2787 (
            .O(N__23458),
            .I(N__23434));
    LocalMux I__2786 (
            .O(N__23455),
            .I(N__23434));
    LocalMux I__2785 (
            .O(N__23452),
            .I(N__23434));
    LocalMux I__2784 (
            .O(N__23449),
            .I(N__23434));
    LocalMux I__2783 (
            .O(N__23446),
            .I(N__23434));
    InMux I__2782 (
            .O(N__23445),
            .I(N__23431));
    Span4Mux_v I__2781 (
            .O(N__23434),
            .I(N__23428));
    LocalMux I__2780 (
            .O(N__23431),
            .I(N_316));
    Odrv4 I__2779 (
            .O(N__23428),
            .I(N_316));
    CEMux I__2778 (
            .O(N__23423),
            .I(N__23419));
    CEMux I__2777 (
            .O(N__23422),
            .I(N__23414));
    LocalMux I__2776 (
            .O(N__23419),
            .I(N__23410));
    CEMux I__2775 (
            .O(N__23418),
            .I(N__23406));
    CEMux I__2774 (
            .O(N__23417),
            .I(N__23403));
    LocalMux I__2773 (
            .O(N__23414),
            .I(N__23400));
    CEMux I__2772 (
            .O(N__23413),
            .I(N__23397));
    Span4Mux_v I__2771 (
            .O(N__23410),
            .I(N__23394));
    CEMux I__2770 (
            .O(N__23409),
            .I(N__23391));
    LocalMux I__2769 (
            .O(N__23406),
            .I(N__23388));
    LocalMux I__2768 (
            .O(N__23403),
            .I(N__23385));
    Span4Mux_h I__2767 (
            .O(N__23400),
            .I(N__23382));
    LocalMux I__2766 (
            .O(N__23397),
            .I(N__23379));
    Span4Mux_h I__2765 (
            .O(N__23394),
            .I(N__23374));
    LocalMux I__2764 (
            .O(N__23391),
            .I(N__23374));
    Span4Mux_v I__2763 (
            .O(N__23388),
            .I(N__23371));
    Span4Mux_h I__2762 (
            .O(N__23385),
            .I(N__23368));
    Span4Mux_h I__2761 (
            .O(N__23382),
            .I(N__23365));
    Span4Mux_v I__2760 (
            .O(N__23379),
            .I(N__23362));
    Span4Mux_h I__2759 (
            .O(N__23374),
            .I(N__23359));
    Span4Mux_h I__2758 (
            .O(N__23371),
            .I(N__23354));
    Span4Mux_h I__2757 (
            .O(N__23368),
            .I(N__23354));
    Odrv4 I__2756 (
            .O(N__23365),
            .I(un1_spointer11_0));
    Odrv4 I__2755 (
            .O(N__23362),
            .I(un1_spointer11_0));
    Odrv4 I__2754 (
            .O(N__23359),
            .I(un1_spointer11_0));
    Odrv4 I__2753 (
            .O(N__23354),
            .I(un1_spointer11_0));
    InMux I__2752 (
            .O(N__23345),
            .I(N__23341));
    InMux I__2751 (
            .O(N__23344),
            .I(N__23337));
    LocalMux I__2750 (
            .O(N__23341),
            .I(N__23334));
    InMux I__2749 (
            .O(N__23340),
            .I(N__23331));
    LocalMux I__2748 (
            .O(N__23337),
            .I(N__23328));
    Span4Mux_h I__2747 (
            .O(N__23334),
            .I(N__23325));
    LocalMux I__2746 (
            .O(N__23331),
            .I(sAddress_RNI6VH7_2Z0Z_1));
    Odrv4 I__2745 (
            .O(N__23328),
            .I(sAddress_RNI6VH7_2Z0Z_1));
    Odrv4 I__2744 (
            .O(N__23325),
            .I(sAddress_RNI6VH7_2Z0Z_1));
    IoInMux I__2743 (
            .O(N__23318),
            .I(N__23315));
    LocalMux I__2742 (
            .O(N__23315),
            .I(N__23312));
    Span12Mux_s0_h I__2741 (
            .O(N__23312),
            .I(N__23309));
    Span12Mux_v I__2740 (
            .O(N__23309),
            .I(N__23306));
    Span12Mux_h I__2739 (
            .O(N__23306),
            .I(N__23303));
    Odrv12 I__2738 (
            .O(N__23303),
            .I(LED_ACQ_obuf_RNOZ0));
    InMux I__2737 (
            .O(N__23300),
            .I(N__23295));
    CascadeMux I__2736 (
            .O(N__23299),
            .I(N__23290));
    CascadeMux I__2735 (
            .O(N__23298),
            .I(N__23287));
    LocalMux I__2734 (
            .O(N__23295),
            .I(N__23284));
    InMux I__2733 (
            .O(N__23294),
            .I(N__23281));
    InMux I__2732 (
            .O(N__23293),
            .I(N__23274));
    InMux I__2731 (
            .O(N__23290),
            .I(N__23274));
    InMux I__2730 (
            .O(N__23287),
            .I(N__23274));
    Odrv4 I__2729 (
            .O(N__23284),
            .I(sAddress_RNI6VH7_3Z0Z_1));
    LocalMux I__2728 (
            .O(N__23281),
            .I(sAddress_RNI6VH7_3Z0Z_1));
    LocalMux I__2727 (
            .O(N__23274),
            .I(sAddress_RNI6VH7_3Z0Z_1));
    CascadeMux I__2726 (
            .O(N__23267),
            .I(sAddress_RNI6VH7_3Z0Z_1_cascade_));
    CEMux I__2725 (
            .O(N__23264),
            .I(N__23261));
    LocalMux I__2724 (
            .O(N__23261),
            .I(N__23258));
    Span4Mux_h I__2723 (
            .O(N__23258),
            .I(N__23255));
    Span4Mux_h I__2722 (
            .O(N__23255),
            .I(N__23252));
    Odrv4 I__2721 (
            .O(N__23252),
            .I(sDAC_mem_10_1_sqmuxa));
    CascadeMux I__2720 (
            .O(N__23249),
            .I(N_326_cascade_));
    CEMux I__2719 (
            .O(N__23246),
            .I(N__23243));
    LocalMux I__2718 (
            .O(N__23243),
            .I(N__23240));
    Span4Mux_v I__2717 (
            .O(N__23240),
            .I(N__23237));
    Odrv4 I__2716 (
            .O(N__23237),
            .I(sDAC_mem_38_1_sqmuxa));
    InMux I__2715 (
            .O(N__23234),
            .I(N__23231));
    LocalMux I__2714 (
            .O(N__23231),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4 ));
    InMux I__2713 (
            .O(N__23228),
            .I(N__23225));
    LocalMux I__2712 (
            .O(N__23225),
            .I(N__23222));
    Odrv12 I__2711 (
            .O(N__23222),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12 ));
    InMux I__2710 (
            .O(N__23219),
            .I(N__23216));
    LocalMux I__2709 (
            .O(N__23216),
            .I(N__23213));
    Span4Mux_h I__2708 (
            .O(N__23213),
            .I(N__23210));
    Odrv4 I__2707 (
            .O(N__23210),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10 ));
    CEMux I__2706 (
            .O(N__23207),
            .I(N__23204));
    LocalMux I__2705 (
            .O(N__23204),
            .I(N__23201));
    Span4Mux_v I__2704 (
            .O(N__23201),
            .I(N__23198));
    Odrv4 I__2703 (
            .O(N__23198),
            .I(sEEPon_1_sqmuxa));
    InMux I__2702 (
            .O(N__23195),
            .I(N__23192));
    LocalMux I__2701 (
            .O(N__23192),
            .I(\spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0 ));
    InMux I__2700 (
            .O(N__23189),
            .I(N__23183));
    InMux I__2699 (
            .O(N__23188),
            .I(N__23183));
    LocalMux I__2698 (
            .O(N__23183),
            .I(\spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0 ));
    InMux I__2697 (
            .O(N__23180),
            .I(N__23177));
    LocalMux I__2696 (
            .O(N__23177),
            .I(N__23174));
    Span4Mux_h I__2695 (
            .O(N__23174),
            .I(N__23171));
    Span4Mux_v I__2694 (
            .O(N__23171),
            .I(N__23167));
    InMux I__2693 (
            .O(N__23170),
            .I(N__23164));
    Odrv4 I__2692 (
            .O(N__23167),
            .I(\spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0 ));
    LocalMux I__2691 (
            .O(N__23164),
            .I(\spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0 ));
    InMux I__2690 (
            .O(N__23159),
            .I(N__23156));
    LocalMux I__2689 (
            .O(N__23156),
            .I(\spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0 ));
    CEMux I__2688 (
            .O(N__23153),
            .I(N__23150));
    LocalMux I__2687 (
            .O(N__23150),
            .I(N__23146));
    CEMux I__2686 (
            .O(N__23149),
            .I(N__23143));
    Span4Mux_h I__2685 (
            .O(N__23146),
            .I(N__23140));
    LocalMux I__2684 (
            .O(N__23143),
            .I(N__23137));
    Odrv4 I__2683 (
            .O(N__23140),
            .I(sDAC_mem_29_1_sqmuxa));
    Odrv12 I__2682 (
            .O(N__23137),
            .I(sDAC_mem_29_1_sqmuxa));
    InMux I__2681 (
            .O(N__23132),
            .I(un1_sTrigCounter_cry_11));
    InMux I__2680 (
            .O(N__23129),
            .I(N__23125));
    InMux I__2679 (
            .O(N__23128),
            .I(N__23122));
    LocalMux I__2678 (
            .O(N__23125),
            .I(sTrigCounterZ0Z_13));
    LocalMux I__2677 (
            .O(N__23122),
            .I(sTrigCounterZ0Z_13));
    InMux I__2676 (
            .O(N__23117),
            .I(un1_sTrigCounter_cry_12));
    InMux I__2675 (
            .O(N__23114),
            .I(N__23110));
    InMux I__2674 (
            .O(N__23113),
            .I(N__23107));
    LocalMux I__2673 (
            .O(N__23110),
            .I(sTrigCounterZ0Z_14));
    LocalMux I__2672 (
            .O(N__23107),
            .I(sTrigCounterZ0Z_14));
    InMux I__2671 (
            .O(N__23102),
            .I(un1_sTrigCounter_cry_13));
    InMux I__2670 (
            .O(N__23099),
            .I(un1_sTrigCounter_cry_14));
    InMux I__2669 (
            .O(N__23096),
            .I(N__23092));
    InMux I__2668 (
            .O(N__23095),
            .I(N__23089));
    LocalMux I__2667 (
            .O(N__23092),
            .I(sTrigCounterZ0Z_15));
    LocalMux I__2666 (
            .O(N__23089),
            .I(sTrigCounterZ0Z_15));
    SRMux I__2665 (
            .O(N__23084),
            .I(N__23080));
    SRMux I__2664 (
            .O(N__23083),
            .I(N__23077));
    LocalMux I__2663 (
            .O(N__23080),
            .I(N_82_i));
    LocalMux I__2662 (
            .O(N__23077),
            .I(N_82_i));
    InMux I__2661 (
            .O(N__23072),
            .I(N__23068));
    InMux I__2660 (
            .O(N__23071),
            .I(N__23065));
    LocalMux I__2659 (
            .O(N__23068),
            .I(sTrigCounterZ0Z_4));
    LocalMux I__2658 (
            .O(N__23065),
            .I(sTrigCounterZ0Z_4));
    InMux I__2657 (
            .O(N__23060),
            .I(un1_sTrigCounter_cry_3));
    InMux I__2656 (
            .O(N__23057),
            .I(N__23053));
    InMux I__2655 (
            .O(N__23056),
            .I(N__23050));
    LocalMux I__2654 (
            .O(N__23053),
            .I(sTrigCounterZ0Z_5));
    LocalMux I__2653 (
            .O(N__23050),
            .I(sTrigCounterZ0Z_5));
    InMux I__2652 (
            .O(N__23045),
            .I(un1_sTrigCounter_cry_4));
    InMux I__2651 (
            .O(N__23042),
            .I(N__23038));
    InMux I__2650 (
            .O(N__23041),
            .I(N__23035));
    LocalMux I__2649 (
            .O(N__23038),
            .I(sTrigCounterZ0Z_6));
    LocalMux I__2648 (
            .O(N__23035),
            .I(sTrigCounterZ0Z_6));
    InMux I__2647 (
            .O(N__23030),
            .I(un1_sTrigCounter_cry_5));
    InMux I__2646 (
            .O(N__23027),
            .I(N__23023));
    InMux I__2645 (
            .O(N__23026),
            .I(N__23020));
    LocalMux I__2644 (
            .O(N__23023),
            .I(sTrigCounterZ0Z_7));
    LocalMux I__2643 (
            .O(N__23020),
            .I(sTrigCounterZ0Z_7));
    InMux I__2642 (
            .O(N__23015),
            .I(un1_sTrigCounter_cry_6));
    InMux I__2641 (
            .O(N__23012),
            .I(N__23008));
    InMux I__2640 (
            .O(N__23011),
            .I(N__23005));
    LocalMux I__2639 (
            .O(N__23008),
            .I(sTrigCounterZ0Z_8));
    LocalMux I__2638 (
            .O(N__23005),
            .I(sTrigCounterZ0Z_8));
    InMux I__2637 (
            .O(N__23000),
            .I(bfn_8_14_0_));
    InMux I__2636 (
            .O(N__22997),
            .I(N__22993));
    InMux I__2635 (
            .O(N__22996),
            .I(N__22990));
    LocalMux I__2634 (
            .O(N__22993),
            .I(sTrigCounterZ0Z_9));
    LocalMux I__2633 (
            .O(N__22990),
            .I(sTrigCounterZ0Z_9));
    InMux I__2632 (
            .O(N__22985),
            .I(un1_sTrigCounter_cry_8));
    InMux I__2631 (
            .O(N__22982),
            .I(N__22978));
    InMux I__2630 (
            .O(N__22981),
            .I(N__22975));
    LocalMux I__2629 (
            .O(N__22978),
            .I(sTrigCounterZ0Z_10));
    LocalMux I__2628 (
            .O(N__22975),
            .I(sTrigCounterZ0Z_10));
    InMux I__2627 (
            .O(N__22970),
            .I(un1_sTrigCounter_cry_9));
    InMux I__2626 (
            .O(N__22967),
            .I(N__22963));
    InMux I__2625 (
            .O(N__22966),
            .I(N__22960));
    LocalMux I__2624 (
            .O(N__22963),
            .I(sTrigCounterZ0Z_11));
    LocalMux I__2623 (
            .O(N__22960),
            .I(sTrigCounterZ0Z_11));
    InMux I__2622 (
            .O(N__22955),
            .I(un1_sTrigCounter_cry_10));
    InMux I__2621 (
            .O(N__22952),
            .I(N__22948));
    InMux I__2620 (
            .O(N__22951),
            .I(N__22945));
    LocalMux I__2619 (
            .O(N__22948),
            .I(sTrigCounterZ0Z_12));
    LocalMux I__2618 (
            .O(N__22945),
            .I(sTrigCounterZ0Z_12));
    InMux I__2617 (
            .O(N__22940),
            .I(N__22931));
    InMux I__2616 (
            .O(N__22939),
            .I(N__22931));
    InMux I__2615 (
            .O(N__22938),
            .I(N__22931));
    LocalMux I__2614 (
            .O(N__22931),
            .I(N__22928));
    Odrv4 I__2613 (
            .O(N__22928),
            .I(un10_trig_prev_cry_15_THRU_CO));
    InMux I__2612 (
            .O(N__22925),
            .I(N__22922));
    LocalMux I__2611 (
            .O(N__22922),
            .I(N_178));
    InMux I__2610 (
            .O(N__22919),
            .I(N__22916));
    LocalMux I__2609 (
            .O(N__22916),
            .I(N__22913));
    Span4Mux_h I__2608 (
            .O(N__22913),
            .I(N__22910));
    Odrv4 I__2607 (
            .O(N__22910),
            .I(un1_scounter_i_0));
    CascadeMux I__2606 (
            .O(N__22907),
            .I(N_178_cascade_));
    InMux I__2605 (
            .O(N__22904),
            .I(N__22901));
    LocalMux I__2604 (
            .O(N__22901),
            .I(N_96));
    CascadeMux I__2603 (
            .O(N__22898),
            .I(N_77_cascade_));
    CascadeMux I__2602 (
            .O(N__22895),
            .I(N__22890));
    CascadeMux I__2601 (
            .O(N__22894),
            .I(N__22887));
    InMux I__2600 (
            .O(N__22893),
            .I(N__22880));
    InMux I__2599 (
            .O(N__22890),
            .I(N__22880));
    InMux I__2598 (
            .O(N__22887),
            .I(N__22880));
    LocalMux I__2597 (
            .O(N__22880),
            .I(sPeriod_prevZ0));
    CascadeMux I__2596 (
            .O(N__22877),
            .I(N__22873));
    InMux I__2595 (
            .O(N__22876),
            .I(N__22870));
    InMux I__2594 (
            .O(N__22873),
            .I(N__22867));
    LocalMux I__2593 (
            .O(N__22870),
            .I(un1_reset_rpi_inv_2_0));
    LocalMux I__2592 (
            .O(N__22867),
            .I(un1_reset_rpi_inv_2_0));
    InMux I__2591 (
            .O(N__22862),
            .I(un1_sTrigCounter_cry_0));
    InMux I__2590 (
            .O(N__22859),
            .I(N__22855));
    InMux I__2589 (
            .O(N__22858),
            .I(N__22852));
    LocalMux I__2588 (
            .O(N__22855),
            .I(sTrigCounterZ0Z_2));
    LocalMux I__2587 (
            .O(N__22852),
            .I(sTrigCounterZ0Z_2));
    InMux I__2586 (
            .O(N__22847),
            .I(un1_sTrigCounter_cry_1));
    InMux I__2585 (
            .O(N__22844),
            .I(N__22840));
    InMux I__2584 (
            .O(N__22843),
            .I(N__22837));
    LocalMux I__2583 (
            .O(N__22840),
            .I(sTrigCounterZ0Z_3));
    LocalMux I__2582 (
            .O(N__22837),
            .I(sTrigCounterZ0Z_3));
    InMux I__2581 (
            .O(N__22832),
            .I(un1_sTrigCounter_cry_2));
    InMux I__2580 (
            .O(N__22829),
            .I(N__22824));
    InMux I__2579 (
            .O(N__22828),
            .I(N__22821));
    InMux I__2578 (
            .O(N__22827),
            .I(N__22818));
    LocalMux I__2577 (
            .O(N__22824),
            .I(N__22813));
    LocalMux I__2576 (
            .O(N__22821),
            .I(N__22813));
    LocalMux I__2575 (
            .O(N__22818),
            .I(N__22810));
    Span4Mux_v I__2574 (
            .O(N__22813),
            .I(N__22807));
    Span12Mux_v I__2573 (
            .O(N__22810),
            .I(N__22802));
    Sp12to4 I__2572 (
            .O(N__22807),
            .I(N__22802));
    Odrv12 I__2571 (
            .O(N__22802),
            .I(trig_rpi_c));
    InMux I__2570 (
            .O(N__22799),
            .I(N__22795));
    InMux I__2569 (
            .O(N__22798),
            .I(N__22792));
    LocalMux I__2568 (
            .O(N__22795),
            .I(N__22789));
    LocalMux I__2567 (
            .O(N__22792),
            .I(N__22786));
    Span4Mux_v I__2566 (
            .O(N__22789),
            .I(N__22782));
    Span4Mux_v I__2565 (
            .O(N__22786),
            .I(N__22779));
    InMux I__2564 (
            .O(N__22785),
            .I(N__22776));
    Sp12to4 I__2563 (
            .O(N__22782),
            .I(N__22769));
    Sp12to4 I__2562 (
            .O(N__22779),
            .I(N__22769));
    LocalMux I__2561 (
            .O(N__22776),
            .I(N__22769));
    Odrv12 I__2560 (
            .O(N__22769),
            .I(trig_ext_c));
    InMux I__2559 (
            .O(N__22766),
            .I(N__22763));
    LocalMux I__2558 (
            .O(N__22763),
            .I(N__22759));
    CascadeMux I__2557 (
            .O(N__22762),
            .I(N__22755));
    Span4Mux_v I__2556 (
            .O(N__22759),
            .I(N__22752));
    InMux I__2555 (
            .O(N__22758),
            .I(N__22749));
    InMux I__2554 (
            .O(N__22755),
            .I(N__22746));
    Sp12to4 I__2553 (
            .O(N__22752),
            .I(N__22739));
    LocalMux I__2552 (
            .O(N__22749),
            .I(N__22739));
    LocalMux I__2551 (
            .O(N__22746),
            .I(N__22739));
    Span12Mux_h I__2550 (
            .O(N__22739),
            .I(N__22736));
    Span12Mux_v I__2549 (
            .O(N__22736),
            .I(N__22733));
    Span12Mux_h I__2548 (
            .O(N__22733),
            .I(N__22730));
    Odrv12 I__2547 (
            .O(N__22730),
            .I(trig_ft_c));
    InMux I__2546 (
            .O(N__22727),
            .I(N__22723));
    InMux I__2545 (
            .O(N__22726),
            .I(N__22720));
    LocalMux I__2544 (
            .O(N__22723),
            .I(N__22717));
    LocalMux I__2543 (
            .O(N__22720),
            .I(N__22711));
    Span4Mux_v I__2542 (
            .O(N__22717),
            .I(N__22711));
    InMux I__2541 (
            .O(N__22716),
            .I(N__22708));
    Odrv4 I__2540 (
            .O(N__22711),
            .I(trig_prevZ0));
    LocalMux I__2539 (
            .O(N__22708),
            .I(trig_prevZ0));
    CascadeMux I__2538 (
            .O(N__22703),
            .I(g3_0_cascade_));
    CascadeMux I__2537 (
            .O(N__22700),
            .I(sAddress_RNI70I7Z0Z_1_cascade_));
    InMux I__2536 (
            .O(N__22697),
            .I(N__22694));
    LocalMux I__2535 (
            .O(N__22694),
            .I(g1_i_a4_0_0));
    InMux I__2534 (
            .O(N__22691),
            .I(N__22688));
    LocalMux I__2533 (
            .O(N__22688),
            .I(N_8_mux));
    CascadeMux I__2532 (
            .O(N__22685),
            .I(N_319_cascade_));
    CEMux I__2531 (
            .O(N__22682),
            .I(N__22679));
    LocalMux I__2530 (
            .O(N__22679),
            .I(N__22676));
    Span4Mux_v I__2529 (
            .O(N__22676),
            .I(N__22673));
    Odrv4 I__2528 (
            .O(N__22673),
            .I(sAddress_RNI9IH12_2Z0Z_1));
    InMux I__2527 (
            .O(N__22670),
            .I(N__22667));
    LocalMux I__2526 (
            .O(N__22667),
            .I(N__22664));
    Span4Mux_v I__2525 (
            .O(N__22664),
            .I(N__22659));
    InMux I__2524 (
            .O(N__22663),
            .I(N__22656));
    InMux I__2523 (
            .O(N__22662),
            .I(N__22653));
    Odrv4 I__2522 (
            .O(N__22659),
            .I(\spi_slave_inst.rx_done_reg2_iZ0 ));
    LocalMux I__2521 (
            .O(N__22656),
            .I(\spi_slave_inst.rx_done_reg2_iZ0 ));
    LocalMux I__2520 (
            .O(N__22653),
            .I(\spi_slave_inst.rx_done_reg2_iZ0 ));
    CascadeMux I__2519 (
            .O(N__22646),
            .I(N__22643));
    InMux I__2518 (
            .O(N__22643),
            .I(N__22640));
    LocalMux I__2517 (
            .O(N__22640),
            .I(N__22637));
    Odrv4 I__2516 (
            .O(N__22637),
            .I(\spi_slave_inst.rx_done_reg3_iZ0 ));
    InMux I__2515 (
            .O(N__22634),
            .I(N__22631));
    LocalMux I__2514 (
            .O(N__22631),
            .I(N__22628));
    Odrv4 I__2513 (
            .O(N__22628),
            .I(\spi_slave_inst.rx_ready_i_RNOZ0Z_0 ));
    CascadeMux I__2512 (
            .O(N__22625),
            .I(sPointer_RNI5LBD1Z0Z_0_cascade_));
    InMux I__2511 (
            .O(N__22622),
            .I(N__22616));
    InMux I__2510 (
            .O(N__22621),
            .I(N__22616));
    LocalMux I__2509 (
            .O(N__22616),
            .I(sDAC_mem_17_1_sqmuxa_0_a2_0_a2_1_0));
    InMux I__2508 (
            .O(N__22613),
            .I(N__22604));
    InMux I__2507 (
            .O(N__22612),
            .I(N__22604));
    InMux I__2506 (
            .O(N__22611),
            .I(N__22599));
    InMux I__2505 (
            .O(N__22610),
            .I(N__22599));
    InMux I__2504 (
            .O(N__22609),
            .I(N__22596));
    LocalMux I__2503 (
            .O(N__22604),
            .I(sAddressZ0Z_4));
    LocalMux I__2502 (
            .O(N__22599),
            .I(sAddressZ0Z_4));
    LocalMux I__2501 (
            .O(N__22596),
            .I(sAddressZ0Z_4));
    CascadeMux I__2500 (
            .O(N__22589),
            .I(sAddress_RNIP2UK1Z0Z_4_cascade_));
    InMux I__2499 (
            .O(N__22586),
            .I(N__22583));
    LocalMux I__2498 (
            .O(N__22583),
            .I(N__22580));
    Span4Mux_v I__2497 (
            .O(N__22580),
            .I(N__22577));
    Span4Mux_v I__2496 (
            .O(N__22577),
            .I(N__22573));
    InMux I__2495 (
            .O(N__22576),
            .I(N__22570));
    Odrv4 I__2494 (
            .O(N__22573),
            .I(\spi_slave_inst.rx_done_neg_sclk_iZ0 ));
    LocalMux I__2493 (
            .O(N__22570),
            .I(\spi_slave_inst.rx_done_neg_sclk_iZ0 ));
    CEMux I__2492 (
            .O(N__22565),
            .I(N__22562));
    LocalMux I__2491 (
            .O(N__22562),
            .I(N__22559));
    Odrv12 I__2490 (
            .O(N__22559),
            .I(\spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541 ));
    InMux I__2489 (
            .O(N__22556),
            .I(N__22550));
    InMux I__2488 (
            .O(N__22555),
            .I(N__22550));
    LocalMux I__2487 (
            .O(N__22550),
            .I(\spi_slave_inst.rx_done_reg1_iZ0 ));
    CascadeMux I__2486 (
            .O(N__22547),
            .I(N_344_cascade_));
    CEMux I__2485 (
            .O(N__22544),
            .I(N__22541));
    LocalMux I__2484 (
            .O(N__22541),
            .I(N__22538));
    Span4Mux_h I__2483 (
            .O(N__22538),
            .I(N__22535));
    Odrv4 I__2482 (
            .O(N__22535),
            .I(sDAC_mem_35_1_sqmuxa));
    InMux I__2481 (
            .O(N__22532),
            .I(N__22529));
    LocalMux I__2480 (
            .O(N__22529),
            .I(sEESingleCont_RNOZ0Z_0));
    InMux I__2479 (
            .O(N__22526),
            .I(N__22523));
    LocalMux I__2478 (
            .O(N__22523),
            .I(N__22519));
    InMux I__2477 (
            .O(N__22522),
            .I(N__22516));
    Span4Mux_v I__2476 (
            .O(N__22519),
            .I(N__22513));
    LocalMux I__2475 (
            .O(N__22516),
            .I(sEESingleContZ0));
    Odrv4 I__2474 (
            .O(N__22513),
            .I(sEESingleContZ0));
    InMux I__2473 (
            .O(N__22508),
            .I(N__22505));
    LocalMux I__2472 (
            .O(N__22505),
            .I(N_1631));
    CascadeMux I__2471 (
            .O(N__22502),
            .I(N__22499));
    InMux I__2470 (
            .O(N__22499),
            .I(N__22496));
    LocalMux I__2469 (
            .O(N__22496),
            .I(sEETrigInternal_3_iv_0_0_i_0));
    CEMux I__2468 (
            .O(N__22493),
            .I(N__22490));
    LocalMux I__2467 (
            .O(N__22490),
            .I(N__22487));
    Odrv12 I__2466 (
            .O(N__22487),
            .I(sDAC_mem_11_1_sqmuxa));
    InMux I__2465 (
            .O(N__22484),
            .I(N__22481));
    LocalMux I__2464 (
            .O(N__22481),
            .I(N__22477));
    InMux I__2463 (
            .O(N__22480),
            .I(N__22474));
    Odrv4 I__2462 (
            .O(N__22477),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0 ));
    LocalMux I__2461 (
            .O(N__22474),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0 ));
    InMux I__2460 (
            .O(N__22469),
            .I(N__22466));
    LocalMux I__2459 (
            .O(N__22466),
            .I(N__22462));
    InMux I__2458 (
            .O(N__22465),
            .I(N__22459));
    Span4Mux_v I__2457 (
            .O(N__22462),
            .I(N__22454));
    LocalMux I__2456 (
            .O(N__22459),
            .I(N__22454));
    Odrv4 I__2455 (
            .O(N__22454),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1 ));
    InMux I__2454 (
            .O(N__22451),
            .I(N__22447));
    InMux I__2453 (
            .O(N__22450),
            .I(N__22444));
    LocalMux I__2452 (
            .O(N__22447),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2 ));
    LocalMux I__2451 (
            .O(N__22444),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2 ));
    InMux I__2450 (
            .O(N__22439),
            .I(N__22435));
    InMux I__2449 (
            .O(N__22438),
            .I(N__22432));
    LocalMux I__2448 (
            .O(N__22435),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3 ));
    LocalMux I__2447 (
            .O(N__22432),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3 ));
    InMux I__2446 (
            .O(N__22427),
            .I(N__22423));
    InMux I__2445 (
            .O(N__22426),
            .I(N__22420));
    LocalMux I__2444 (
            .O(N__22423),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4 ));
    LocalMux I__2443 (
            .O(N__22420),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4 ));
    InMux I__2442 (
            .O(N__22415),
            .I(N__22411));
    InMux I__2441 (
            .O(N__22414),
            .I(N__22408));
    LocalMux I__2440 (
            .O(N__22411),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5 ));
    LocalMux I__2439 (
            .O(N__22408),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5 ));
    InMux I__2438 (
            .O(N__22403),
            .I(N__22399));
    InMux I__2437 (
            .O(N__22402),
            .I(N__22396));
    LocalMux I__2436 (
            .O(N__22399),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6 ));
    LocalMux I__2435 (
            .O(N__22396),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6 ));
    InMux I__2434 (
            .O(N__22391),
            .I(N__22388));
    LocalMux I__2433 (
            .O(N__22388),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7 ));
    CascadeMux I__2432 (
            .O(N__22385),
            .I(N__22382));
    InMux I__2431 (
            .O(N__22382),
            .I(N__22378));
    CascadeMux I__2430 (
            .O(N__22381),
            .I(N__22375));
    LocalMux I__2429 (
            .O(N__22378),
            .I(N__22372));
    InMux I__2428 (
            .O(N__22375),
            .I(N__22369));
    Odrv4 I__2427 (
            .O(N__22372),
            .I(un3_trig_0));
    LocalMux I__2426 (
            .O(N__22369),
            .I(un3_trig_0));
    CascadeMux I__2425 (
            .O(N__22364),
            .I(N__22361));
    InMux I__2424 (
            .O(N__22361),
            .I(N__22358));
    LocalMux I__2423 (
            .O(N__22358),
            .I(sEEADC_freqZ0Z_5));
    InMux I__2422 (
            .O(N__22355),
            .I(N__22352));
    LocalMux I__2421 (
            .O(N__22352),
            .I(N__22349));
    Span4Mux_v I__2420 (
            .O(N__22349),
            .I(N__22346));
    Sp12to4 I__2419 (
            .O(N__22346),
            .I(N__22343));
    Span12Mux_h I__2418 (
            .O(N__22343),
            .I(N__22340));
    Odrv12 I__2417 (
            .O(N__22340),
            .I(spi_mosi_rpi_c));
    InMux I__2416 (
            .O(N__22337),
            .I(N__22334));
    LocalMux I__2415 (
            .O(N__22334),
            .I(N__22331));
    Span4Mux_v I__2414 (
            .O(N__22331),
            .I(N__22328));
    Span4Mux_h I__2413 (
            .O(N__22328),
            .I(N__22325));
    Sp12to4 I__2412 (
            .O(N__22325),
            .I(N__22322));
    Span12Mux_h I__2411 (
            .O(N__22322),
            .I(N__22319));
    Odrv12 I__2410 (
            .O(N__22319),
            .I(spi_mosi_ft_c));
    InMux I__2409 (
            .O(N__22316),
            .I(N__22313));
    LocalMux I__2408 (
            .O(N__22313),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11 ));
    CascadeMux I__2407 (
            .O(N__22310),
            .I(N__22307));
    InMux I__2406 (
            .O(N__22307),
            .I(N__22304));
    LocalMux I__2405 (
            .O(N__22304),
            .I(un10_trig_prev_14));
    InMux I__2404 (
            .O(N__22301),
            .I(N__22298));
    LocalMux I__2403 (
            .O(N__22298),
            .I(sTrigCounter_i_14));
    CascadeMux I__2402 (
            .O(N__22295),
            .I(N__22292));
    InMux I__2401 (
            .O(N__22292),
            .I(N__22289));
    LocalMux I__2400 (
            .O(N__22289),
            .I(un10_trig_prev_15));
    InMux I__2399 (
            .O(N__22286),
            .I(N__22283));
    LocalMux I__2398 (
            .O(N__22283),
            .I(sTrigCounter_i_15));
    InMux I__2397 (
            .O(N__22280),
            .I(bfn_7_14_0_));
    InMux I__2396 (
            .O(N__22277),
            .I(N__22274));
    LocalMux I__2395 (
            .O(N__22274),
            .I(N_173));
    InMux I__2394 (
            .O(N__22271),
            .I(N__22268));
    LocalMux I__2393 (
            .O(N__22268),
            .I(sEEADC_freqZ0Z_4));
    CascadeMux I__2392 (
            .O(N__22265),
            .I(N__22262));
    InMux I__2391 (
            .O(N__22262),
            .I(N__22259));
    LocalMux I__2390 (
            .O(N__22259),
            .I(un10_trig_prev_6));
    InMux I__2389 (
            .O(N__22256),
            .I(N__22253));
    LocalMux I__2388 (
            .O(N__22253),
            .I(sTrigCounter_i_6));
    CascadeMux I__2387 (
            .O(N__22250),
            .I(N__22247));
    InMux I__2386 (
            .O(N__22247),
            .I(N__22244));
    LocalMux I__2385 (
            .O(N__22244),
            .I(un10_trig_prev_7));
    InMux I__2384 (
            .O(N__22241),
            .I(N__22238));
    LocalMux I__2383 (
            .O(N__22238),
            .I(sTrigCounter_i_7));
    CascadeMux I__2382 (
            .O(N__22235),
            .I(N__22232));
    InMux I__2381 (
            .O(N__22232),
            .I(N__22229));
    LocalMux I__2380 (
            .O(N__22229),
            .I(un10_trig_prev_8));
    InMux I__2379 (
            .O(N__22226),
            .I(N__22223));
    LocalMux I__2378 (
            .O(N__22223),
            .I(sTrigCounter_i_8));
    CascadeMux I__2377 (
            .O(N__22220),
            .I(N__22217));
    InMux I__2376 (
            .O(N__22217),
            .I(N__22214));
    LocalMux I__2375 (
            .O(N__22214),
            .I(un10_trig_prev_9));
    InMux I__2374 (
            .O(N__22211),
            .I(N__22208));
    LocalMux I__2373 (
            .O(N__22208),
            .I(sTrigCounter_i_9));
    CascadeMux I__2372 (
            .O(N__22205),
            .I(N__22202));
    InMux I__2371 (
            .O(N__22202),
            .I(N__22199));
    LocalMux I__2370 (
            .O(N__22199),
            .I(un10_trig_prev_10));
    InMux I__2369 (
            .O(N__22196),
            .I(N__22193));
    LocalMux I__2368 (
            .O(N__22193),
            .I(sTrigCounter_i_10));
    CascadeMux I__2367 (
            .O(N__22190),
            .I(N__22187));
    InMux I__2366 (
            .O(N__22187),
            .I(N__22184));
    LocalMux I__2365 (
            .O(N__22184),
            .I(un10_trig_prev_11));
    InMux I__2364 (
            .O(N__22181),
            .I(N__22178));
    LocalMux I__2363 (
            .O(N__22178),
            .I(sTrigCounter_i_11));
    CascadeMux I__2362 (
            .O(N__22175),
            .I(N__22172));
    InMux I__2361 (
            .O(N__22172),
            .I(N__22169));
    LocalMux I__2360 (
            .O(N__22169),
            .I(un10_trig_prev_12));
    InMux I__2359 (
            .O(N__22166),
            .I(N__22163));
    LocalMux I__2358 (
            .O(N__22163),
            .I(sTrigCounter_i_12));
    CascadeMux I__2357 (
            .O(N__22160),
            .I(N__22157));
    InMux I__2356 (
            .O(N__22157),
            .I(N__22154));
    LocalMux I__2355 (
            .O(N__22154),
            .I(un10_trig_prev_13));
    InMux I__2354 (
            .O(N__22151),
            .I(N__22148));
    LocalMux I__2353 (
            .O(N__22148),
            .I(sTrigCounter_i_13));
    CascadeMux I__2352 (
            .O(N__22145),
            .I(N__22141));
    InMux I__2351 (
            .O(N__22144),
            .I(N__22138));
    InMux I__2350 (
            .O(N__22141),
            .I(N__22135));
    LocalMux I__2349 (
            .O(N__22138),
            .I(un8_trig_prev_0));
    LocalMux I__2348 (
            .O(N__22135),
            .I(un8_trig_prev_0));
    CascadeMux I__2347 (
            .O(N__22130),
            .I(N__22127));
    InMux I__2346 (
            .O(N__22127),
            .I(N__22124));
    LocalMux I__2345 (
            .O(N__22124),
            .I(un10_trig_prev_0));
    InMux I__2344 (
            .O(N__22121),
            .I(N__22118));
    LocalMux I__2343 (
            .O(N__22118),
            .I(sTrigCounter_i_0));
    CascadeMux I__2342 (
            .O(N__22115),
            .I(N__22112));
    InMux I__2341 (
            .O(N__22112),
            .I(N__22109));
    LocalMux I__2340 (
            .O(N__22109),
            .I(un10_trig_prev_1));
    InMux I__2339 (
            .O(N__22106),
            .I(N__22103));
    LocalMux I__2338 (
            .O(N__22103),
            .I(sTrigCounter_i_1));
    CascadeMux I__2337 (
            .O(N__22100),
            .I(N__22097));
    InMux I__2336 (
            .O(N__22097),
            .I(N__22094));
    LocalMux I__2335 (
            .O(N__22094),
            .I(un10_trig_prev_2));
    InMux I__2334 (
            .O(N__22091),
            .I(N__22088));
    LocalMux I__2333 (
            .O(N__22088),
            .I(sTrigCounter_i_2));
    CascadeMux I__2332 (
            .O(N__22085),
            .I(N__22082));
    InMux I__2331 (
            .O(N__22082),
            .I(N__22079));
    LocalMux I__2330 (
            .O(N__22079),
            .I(un10_trig_prev_3));
    InMux I__2329 (
            .O(N__22076),
            .I(N__22073));
    LocalMux I__2328 (
            .O(N__22073),
            .I(sTrigCounter_i_3));
    CascadeMux I__2327 (
            .O(N__22070),
            .I(N__22067));
    InMux I__2326 (
            .O(N__22067),
            .I(N__22064));
    LocalMux I__2325 (
            .O(N__22064),
            .I(un10_trig_prev_4));
    InMux I__2324 (
            .O(N__22061),
            .I(N__22058));
    LocalMux I__2323 (
            .O(N__22058),
            .I(sTrigCounter_i_4));
    CascadeMux I__2322 (
            .O(N__22055),
            .I(N__22052));
    InMux I__2321 (
            .O(N__22052),
            .I(N__22049));
    LocalMux I__2320 (
            .O(N__22049),
            .I(un10_trig_prev_5));
    InMux I__2319 (
            .O(N__22046),
            .I(N__22043));
    LocalMux I__2318 (
            .O(N__22043),
            .I(sTrigCounter_i_5));
    InMux I__2317 (
            .O(N__22040),
            .I(N__22036));
    InMux I__2316 (
            .O(N__22039),
            .I(N__22033));
    LocalMux I__2315 (
            .O(N__22036),
            .I(N__22030));
    LocalMux I__2314 (
            .O(N__22033),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2 ));
    Odrv4 I__2313 (
            .O(N__22030),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2 ));
    InMux I__2312 (
            .O(N__22025),
            .I(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1 ));
    InMux I__2311 (
            .O(N__22022),
            .I(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2 ));
    InMux I__2310 (
            .O(N__22019),
            .I(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3 ));
    InMux I__2309 (
            .O(N__22016),
            .I(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4 ));
    InMux I__2308 (
            .O(N__22013),
            .I(N__22009));
    InMux I__2307 (
            .O(N__22012),
            .I(N__22006));
    LocalMux I__2306 (
            .O(N__22009),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5 ));
    LocalMux I__2305 (
            .O(N__22006),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5 ));
    InMux I__2304 (
            .O(N__22001),
            .I(N__21998));
    LocalMux I__2303 (
            .O(N__21998),
            .I(N__21995));
    Span4Mux_h I__2302 (
            .O(N__21995),
            .I(N__21988));
    InMux I__2301 (
            .O(N__21994),
            .I(N__21983));
    InMux I__2300 (
            .O(N__21993),
            .I(N__21983));
    InMux I__2299 (
            .O(N__21992),
            .I(N__21978));
    InMux I__2298 (
            .O(N__21991),
            .I(N__21978));
    Odrv4 I__2297 (
            .O(N__21988),
            .I(spi_mosi_ready));
    LocalMux I__2296 (
            .O(N__21983),
            .I(spi_mosi_ready));
    LocalMux I__2295 (
            .O(N__21978),
            .I(spi_mosi_ready));
    InMux I__2294 (
            .O(N__21971),
            .I(N__21967));
    InMux I__2293 (
            .O(N__21970),
            .I(N__21964));
    LocalMux I__2292 (
            .O(N__21967),
            .I(spi_mosi_ready_prevZ0));
    LocalMux I__2291 (
            .O(N__21964),
            .I(spi_mosi_ready_prevZ0));
    InMux I__2290 (
            .O(N__21959),
            .I(N__21955));
    InMux I__2289 (
            .O(N__21958),
            .I(N__21952));
    LocalMux I__2288 (
            .O(N__21955),
            .I(spi_mosi_ready_prevZ0Z2));
    LocalMux I__2287 (
            .O(N__21952),
            .I(spi_mosi_ready_prevZ0Z2));
    CascadeMux I__2286 (
            .O(N__21947),
            .I(N__21944));
    InMux I__2285 (
            .O(N__21944),
            .I(N__21941));
    LocalMux I__2284 (
            .O(N__21941),
            .I(spi_mosi_ready_prevZ0Z3));
    CascadeMux I__2283 (
            .O(N__21938),
            .I(N_346_i_cascade_));
    CascadeMux I__2282 (
            .O(N__21935),
            .I(un1_spointer11_8_0_0_a2_1_cascade_));
    CEMux I__2281 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__2280 (
            .O(N__21929),
            .I(N__21926));
    Span4Mux_v I__2279 (
            .O(N__21926),
            .I(N__21923));
    Odrv4 I__2278 (
            .O(N__21923),
            .I(sAddress_RNI7G5E2Z0Z_6));
    InMux I__2277 (
            .O(N__21920),
            .I(N__21910));
    InMux I__2276 (
            .O(N__21919),
            .I(N__21910));
    InMux I__2275 (
            .O(N__21918),
            .I(N__21910));
    CascadeMux I__2274 (
            .O(N__21917),
            .I(N__21907));
    LocalMux I__2273 (
            .O(N__21910),
            .I(N__21904));
    InMux I__2272 (
            .O(N__21907),
            .I(N__21901));
    Span4Mux_v I__2271 (
            .O(N__21904),
            .I(N__21896));
    LocalMux I__2270 (
            .O(N__21901),
            .I(N__21896));
    Span4Mux_h I__2269 (
            .O(N__21896),
            .I(N__21893));
    Odrv4 I__2268 (
            .O(N__21893),
            .I(sAddressZ0Z_7));
    InMux I__2267 (
            .O(N__21890),
            .I(N__21881));
    InMux I__2266 (
            .O(N__21889),
            .I(N__21881));
    InMux I__2265 (
            .O(N__21888),
            .I(N__21881));
    LocalMux I__2264 (
            .O(N__21881),
            .I(N__21877));
    InMux I__2263 (
            .O(N__21880),
            .I(N__21874));
    Span4Mux_v I__2262 (
            .O(N__21877),
            .I(N__21869));
    LocalMux I__2261 (
            .O(N__21874),
            .I(N__21869));
    Span4Mux_h I__2260 (
            .O(N__21869),
            .I(N__21866));
    Odrv4 I__2259 (
            .O(N__21866),
            .I(sAddressZ0Z_6));
    CascadeMux I__2258 (
            .O(N__21863),
            .I(N__21860));
    InMux I__2257 (
            .O(N__21860),
            .I(N__21856));
    InMux I__2256 (
            .O(N__21859),
            .I(N__21853));
    LocalMux I__2255 (
            .O(N__21856),
            .I(N__21850));
    LocalMux I__2254 (
            .O(N__21853),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0 ));
    Odrv4 I__2253 (
            .O(N__21850),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0 ));
    InMux I__2252 (
            .O(N__21845),
            .I(N__21841));
    InMux I__2251 (
            .O(N__21844),
            .I(N__21838));
    LocalMux I__2250 (
            .O(N__21841),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1 ));
    LocalMux I__2249 (
            .O(N__21838),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1 ));
    InMux I__2248 (
            .O(N__21833),
            .I(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0 ));
    CascadeMux I__2247 (
            .O(N__21830),
            .I(N_316_cascade_));
    CascadeMux I__2246 (
            .O(N__21827),
            .I(N_317_cascade_));
    CascadeMux I__2245 (
            .O(N__21824),
            .I(sAddress_RNI8U0V1Z0Z_1_cascade_));
    InMux I__2244 (
            .O(N__21821),
            .I(N__21818));
    LocalMux I__2243 (
            .O(N__21818),
            .I(sAddress_RNI8U0V1Z0Z_1));
    CascadeMux I__2242 (
            .O(N__21815),
            .I(N_454_cascade_));
    CascadeMux I__2241 (
            .O(N__21812),
            .I(N__21809));
    InMux I__2240 (
            .O(N__21809),
            .I(N__21806));
    LocalMux I__2239 (
            .O(N__21806),
            .I(sEETrigCounterZ0Z_9));
    InMux I__2238 (
            .O(N__21803),
            .I(N__21800));
    LocalMux I__2237 (
            .O(N__21800),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11 ));
    InMux I__2236 (
            .O(N__21797),
            .I(N__21794));
    LocalMux I__2235 (
            .O(N__21794),
            .I(N__21791));
    Span4Mux_v I__2234 (
            .O(N__21791),
            .I(N__21788));
    Odrv4 I__2233 (
            .O(N__21788),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1 ));
    InMux I__2232 (
            .O(N__21785),
            .I(N__21782));
    LocalMux I__2231 (
            .O(N__21782),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5 ));
    InMux I__2230 (
            .O(N__21779),
            .I(N__21776));
    LocalMux I__2229 (
            .O(N__21776),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13 ));
    InMux I__2228 (
            .O(N__21773),
            .I(N__21770));
    LocalMux I__2227 (
            .O(N__21770),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14 ));
    InMux I__2226 (
            .O(N__21767),
            .I(N__21764));
    LocalMux I__2225 (
            .O(N__21764),
            .I(N__21761));
    Odrv4 I__2224 (
            .O(N__21761),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0 ));
    InMux I__2223 (
            .O(N__21758),
            .I(N__21755));
    LocalMux I__2222 (
            .O(N__21755),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_6 ));
    InMux I__2221 (
            .O(N__21752),
            .I(N__21749));
    LocalMux I__2220 (
            .O(N__21749),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_5 ));
    InMux I__2219 (
            .O(N__21746),
            .I(un8_trig_prev_0_cry_13));
    InMux I__2218 (
            .O(N__21743),
            .I(un8_trig_prev_0_cry_14));
    CascadeMux I__2217 (
            .O(N__21740),
            .I(N__21737));
    InMux I__2216 (
            .O(N__21737),
            .I(N__21734));
    LocalMux I__2215 (
            .O(N__21734),
            .I(sEETrigCounterZ0Z_10));
    CascadeMux I__2214 (
            .O(N__21731),
            .I(N__21728));
    InMux I__2213 (
            .O(N__21728),
            .I(N__21725));
    LocalMux I__2212 (
            .O(N__21725),
            .I(sEETrigCounterZ0Z_11));
    CascadeMux I__2211 (
            .O(N__21722),
            .I(N__21719));
    InMux I__2210 (
            .O(N__21719),
            .I(N__21716));
    LocalMux I__2209 (
            .O(N__21716),
            .I(sEETrigCounterZ0Z_12));
    CascadeMux I__2208 (
            .O(N__21713),
            .I(N__21710));
    InMux I__2207 (
            .O(N__21710),
            .I(N__21707));
    LocalMux I__2206 (
            .O(N__21707),
            .I(sEETrigCounterZ0Z_13));
    CascadeMux I__2205 (
            .O(N__21704),
            .I(N__21701));
    InMux I__2204 (
            .O(N__21701),
            .I(N__21698));
    LocalMux I__2203 (
            .O(N__21698),
            .I(sEETrigCounterZ0Z_14));
    InMux I__2202 (
            .O(N__21695),
            .I(N__21692));
    LocalMux I__2201 (
            .O(N__21692),
            .I(sEETrigCounterZ0Z_15));
    CascadeMux I__2200 (
            .O(N__21689),
            .I(N__21686));
    InMux I__2199 (
            .O(N__21686),
            .I(N__21683));
    LocalMux I__2198 (
            .O(N__21683),
            .I(sEETrigCounterZ0Z_8));
    CascadeMux I__2197 (
            .O(N__21680),
            .I(N__21677));
    InMux I__2196 (
            .O(N__21677),
            .I(N__21674));
    LocalMux I__2195 (
            .O(N__21674),
            .I(sEETrigCounterZ0Z_5));
    InMux I__2194 (
            .O(N__21671),
            .I(un8_trig_prev_0_cry_4));
    CascadeMux I__2193 (
            .O(N__21668),
            .I(N__21665));
    InMux I__2192 (
            .O(N__21665),
            .I(N__21662));
    LocalMux I__2191 (
            .O(N__21662),
            .I(sEETrigCounterZ0Z_6));
    InMux I__2190 (
            .O(N__21659),
            .I(un8_trig_prev_0_cry_5));
    CascadeMux I__2189 (
            .O(N__21656),
            .I(N__21653));
    InMux I__2188 (
            .O(N__21653),
            .I(N__21650));
    LocalMux I__2187 (
            .O(N__21650),
            .I(sEETrigCounterZ0Z_7));
    InMux I__2186 (
            .O(N__21647),
            .I(un8_trig_prev_0_cry_6));
    InMux I__2185 (
            .O(N__21644),
            .I(bfn_6_13_0_));
    InMux I__2184 (
            .O(N__21641),
            .I(un8_trig_prev_0_cry_8));
    InMux I__2183 (
            .O(N__21638),
            .I(un8_trig_prev_0_cry_9));
    InMux I__2182 (
            .O(N__21635),
            .I(un8_trig_prev_0_cry_10));
    InMux I__2181 (
            .O(N__21632),
            .I(un8_trig_prev_0_cry_11));
    InMux I__2180 (
            .O(N__21629),
            .I(un8_trig_prev_0_cry_12));
    CascadeMux I__2179 (
            .O(N__21626),
            .I(N__21623));
    InMux I__2178 (
            .O(N__21623),
            .I(N__21620));
    LocalMux I__2177 (
            .O(N__21620),
            .I(sEETrigCounterZ0Z_1));
    InMux I__2176 (
            .O(N__21617),
            .I(un8_trig_prev_0_cry_0));
    CascadeMux I__2175 (
            .O(N__21614),
            .I(N__21611));
    InMux I__2174 (
            .O(N__21611),
            .I(N__21608));
    LocalMux I__2173 (
            .O(N__21608),
            .I(sEETrigCounterZ0Z_2));
    InMux I__2172 (
            .O(N__21605),
            .I(un8_trig_prev_0_cry_1));
    CascadeMux I__2171 (
            .O(N__21602),
            .I(N__21599));
    InMux I__2170 (
            .O(N__21599),
            .I(N__21596));
    LocalMux I__2169 (
            .O(N__21596),
            .I(sEETrigCounterZ0Z_3));
    InMux I__2168 (
            .O(N__21593),
            .I(un8_trig_prev_0_cry_2));
    CascadeMux I__2167 (
            .O(N__21590),
            .I(N__21587));
    InMux I__2166 (
            .O(N__21587),
            .I(N__21584));
    LocalMux I__2165 (
            .O(N__21584),
            .I(sEETrigCounterZ0Z_4));
    InMux I__2164 (
            .O(N__21581),
            .I(un8_trig_prev_0_cry_3));
    InMux I__2163 (
            .O(N__21578),
            .I(N__21574));
    CascadeMux I__2162 (
            .O(N__21577),
            .I(N__21571));
    LocalMux I__2161 (
            .O(N__21574),
            .I(N__21567));
    InMux I__2160 (
            .O(N__21571),
            .I(N__21564));
    InMux I__2159 (
            .O(N__21570),
            .I(N__21560));
    Span4Mux_v I__2158 (
            .O(N__21567),
            .I(N__21555));
    LocalMux I__2157 (
            .O(N__21564),
            .I(N__21555));
    InMux I__2156 (
            .O(N__21563),
            .I(N__21552));
    LocalMux I__2155 (
            .O(N__21560),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0 ));
    Odrv4 I__2154 (
            .O(N__21555),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0 ));
    LocalMux I__2153 (
            .O(N__21552),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0 ));
    InMux I__2152 (
            .O(N__21545),
            .I(N__21541));
    InMux I__2151 (
            .O(N__21544),
            .I(N__21538));
    LocalMux I__2150 (
            .O(N__21541),
            .I(N__21535));
    LocalMux I__2149 (
            .O(N__21538),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5 ));
    Odrv12 I__2148 (
            .O(N__21535),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5 ));
    CascadeMux I__2147 (
            .O(N__21530),
            .I(N__21527));
    InMux I__2146 (
            .O(N__21527),
            .I(N__21523));
    InMux I__2145 (
            .O(N__21526),
            .I(N__21520));
    LocalMux I__2144 (
            .O(N__21523),
            .I(N__21517));
    LocalMux I__2143 (
            .O(N__21520),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4 ));
    Odrv12 I__2142 (
            .O(N__21517),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4 ));
    InMux I__2141 (
            .O(N__21512),
            .I(N__21508));
    InMux I__2140 (
            .O(N__21511),
            .I(N__21505));
    LocalMux I__2139 (
            .O(N__21508),
            .I(N__21498));
    LocalMux I__2138 (
            .O(N__21505),
            .I(N__21498));
    InMux I__2137 (
            .O(N__21504),
            .I(N__21495));
    InMux I__2136 (
            .O(N__21503),
            .I(N__21491));
    Span4Mux_v I__2135 (
            .O(N__21498),
            .I(N__21486));
    LocalMux I__2134 (
            .O(N__21495),
            .I(N__21486));
    InMux I__2133 (
            .O(N__21494),
            .I(N__21483));
    LocalMux I__2132 (
            .O(N__21491),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1 ));
    Odrv4 I__2131 (
            .O(N__21486),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1 ));
    LocalMux I__2130 (
            .O(N__21483),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1 ));
    InMux I__2129 (
            .O(N__21476),
            .I(N__21472));
    InMux I__2128 (
            .O(N__21475),
            .I(N__21469));
    LocalMux I__2127 (
            .O(N__21472),
            .I(N__21466));
    LocalMux I__2126 (
            .O(N__21469),
            .I(N__21463));
    Odrv4 I__2125 (
            .O(N__21466),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3 ));
    Odrv4 I__2124 (
            .O(N__21463),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3 ));
    InMux I__2123 (
            .O(N__21458),
            .I(N__21454));
    InMux I__2122 (
            .O(N__21457),
            .I(N__21451));
    LocalMux I__2121 (
            .O(N__21454),
            .I(spi_mosi_ready64_prevZ0Z2));
    LocalMux I__2120 (
            .O(N__21451),
            .I(spi_mosi_ready64_prevZ0Z2));
    InMux I__2119 (
            .O(N__21446),
            .I(N__21442));
    InMux I__2118 (
            .O(N__21445),
            .I(N__21439));
    LocalMux I__2117 (
            .O(N__21442),
            .I(spi_mosi_ready64_prevZ0));
    LocalMux I__2116 (
            .O(N__21439),
            .I(spi_mosi_ready64_prevZ0));
    CascadeMux I__2115 (
            .O(N__21434),
            .I(N__21431));
    InMux I__2114 (
            .O(N__21431),
            .I(N__21428));
    LocalMux I__2113 (
            .O(N__21428),
            .I(spi_mosi_ready64_prevZ0Z3));
    CascadeMux I__2112 (
            .O(N__21425),
            .I(spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_));
    InMux I__2111 (
            .O(N__21422),
            .I(N__21418));
    InMux I__2110 (
            .O(N__21421),
            .I(N__21412));
    LocalMux I__2109 (
            .O(N__21418),
            .I(N__21409));
    InMux I__2108 (
            .O(N__21417),
            .I(N__21406));
    InMux I__2107 (
            .O(N__21416),
            .I(N__21403));
    CascadeMux I__2106 (
            .O(N__21415),
            .I(N__21397));
    LocalMux I__2105 (
            .O(N__21412),
            .I(N__21394));
    Span4Mux_h I__2104 (
            .O(N__21409),
            .I(N__21387));
    LocalMux I__2103 (
            .O(N__21406),
            .I(N__21387));
    LocalMux I__2102 (
            .O(N__21403),
            .I(N__21387));
    InMux I__2101 (
            .O(N__21402),
            .I(N__21384));
    InMux I__2100 (
            .O(N__21401),
            .I(N__21379));
    InMux I__2099 (
            .O(N__21400),
            .I(N__21379));
    InMux I__2098 (
            .O(N__21397),
            .I(N__21376));
    Odrv12 I__2097 (
            .O(N__21394),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ));
    Odrv4 I__2096 (
            .O(N__21387),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ));
    LocalMux I__2095 (
            .O(N__21384),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ));
    LocalMux I__2094 (
            .O(N__21379),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ));
    LocalMux I__2093 (
            .O(N__21376),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ));
    InMux I__2092 (
            .O(N__21365),
            .I(N__21362));
    LocalMux I__2091 (
            .O(N__21362),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO ));
    InMux I__2090 (
            .O(N__21359),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1 ));
    InMux I__2089 (
            .O(N__21356),
            .I(N__21353));
    LocalMux I__2088 (
            .O(N__21353),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO ));
    InMux I__2087 (
            .O(N__21350),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2 ));
    InMux I__2086 (
            .O(N__21347),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3 ));
    InMux I__2085 (
            .O(N__21344),
            .I(bfn_6_8_0_));
    InMux I__2084 (
            .O(N__21341),
            .I(N__21338));
    LocalMux I__2083 (
            .O(N__21338),
            .I(N__21335));
    Odrv4 I__2082 (
            .O(N__21335),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO ));
    CascadeMux I__2081 (
            .O(N__21332),
            .I(N__21328));
    InMux I__2080 (
            .O(N__21331),
            .I(N__21321));
    InMux I__2079 (
            .O(N__21328),
            .I(N__21321));
    InMux I__2078 (
            .O(N__21327),
            .I(N__21316));
    InMux I__2077 (
            .O(N__21326),
            .I(N__21316));
    LocalMux I__2076 (
            .O(N__21321),
            .I(N__21313));
    LocalMux I__2075 (
            .O(N__21316),
            .I(N__21310));
    Odrv4 I__2074 (
            .O(N__21313),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6 ));
    Odrv4 I__2073 (
            .O(N__21310),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6 ));
    CascadeMux I__2072 (
            .O(N__21305),
            .I(N__21301));
    CascadeMux I__2071 (
            .O(N__21304),
            .I(N__21298));
    InMux I__2070 (
            .O(N__21301),
            .I(N__21291));
    InMux I__2069 (
            .O(N__21298),
            .I(N__21291));
    CEMux I__2068 (
            .O(N__21297),
            .I(N__21288));
    CascadeMux I__2067 (
            .O(N__21296),
            .I(N__21285));
    LocalMux I__2066 (
            .O(N__21291),
            .I(N__21277));
    LocalMux I__2065 (
            .O(N__21288),
            .I(N__21277));
    InMux I__2064 (
            .O(N__21285),
            .I(N__21274));
    InMux I__2063 (
            .O(N__21284),
            .I(N__21269));
    InMux I__2062 (
            .O(N__21283),
            .I(N__21269));
    InMux I__2061 (
            .O(N__21282),
            .I(N__21266));
    Span4Mux_v I__2060 (
            .O(N__21277),
            .I(N__21263));
    LocalMux I__2059 (
            .O(N__21274),
            .I(\spi_master_inst.o_sclk_RNIH6AC ));
    LocalMux I__2058 (
            .O(N__21269),
            .I(\spi_master_inst.o_sclk_RNIH6AC ));
    LocalMux I__2057 (
            .O(N__21266),
            .I(\spi_master_inst.o_sclk_RNIH6AC ));
    Odrv4 I__2056 (
            .O(N__21263),
            .I(\spi_master_inst.o_sclk_RNIH6AC ));
    InMux I__2055 (
            .O(N__21254),
            .I(N__21250));
    InMux I__2054 (
            .O(N__21253),
            .I(N__21247));
    LocalMux I__2053 (
            .O(N__21250),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2 ));
    LocalMux I__2052 (
            .O(N__21247),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2 ));
    InMux I__2051 (
            .O(N__21242),
            .I(N__21239));
    LocalMux I__2050 (
            .O(N__21239),
            .I(\spi_master_inst.spi_data_path_u1.N_1411 ));
    InMux I__2049 (
            .O(N__21236),
            .I(N__21233));
    LocalMux I__2048 (
            .O(N__21233),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13 ));
    InMux I__2047 (
            .O(N__21230),
            .I(N__21227));
    LocalMux I__2046 (
            .O(N__21227),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14 ));
    InMux I__2045 (
            .O(N__21224),
            .I(N__21221));
    LocalMux I__2044 (
            .O(N__21221),
            .I(\spi_master_inst.spi_data_path_u1.N_1418 ));
    InMux I__2043 (
            .O(N__21218),
            .I(N__21215));
    LocalMux I__2042 (
            .O(N__21215),
            .I(N__21212));
    Odrv4 I__2041 (
            .O(N__21212),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6 ));
    InMux I__2040 (
            .O(N__21209),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0 ));
    InMux I__2039 (
            .O(N__21206),
            .I(N__21202));
    InMux I__2038 (
            .O(N__21205),
            .I(N__21199));
    LocalMux I__2037 (
            .O(N__21202),
            .I(N__21194));
    LocalMux I__2036 (
            .O(N__21199),
            .I(N__21194));
    Odrv4 I__2035 (
            .O(N__21194),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6 ));
    InMux I__2034 (
            .O(N__21191),
            .I(N__21187));
    InMux I__2033 (
            .O(N__21190),
            .I(N__21184));
    LocalMux I__2032 (
            .O(N__21187),
            .I(N__21181));
    LocalMux I__2031 (
            .O(N__21184),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5 ));
    Odrv4 I__2030 (
            .O(N__21181),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5 ));
    CascadeMux I__2029 (
            .O(N__21176),
            .I(N__21173));
    InMux I__2028 (
            .O(N__21173),
            .I(N__21169));
    InMux I__2027 (
            .O(N__21172),
            .I(N__21166));
    LocalMux I__2026 (
            .O(N__21169),
            .I(N__21163));
    LocalMux I__2025 (
            .O(N__21166),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7 ));
    Odrv4 I__2024 (
            .O(N__21163),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7 ));
    InMux I__2023 (
            .O(N__21158),
            .I(N__21154));
    InMux I__2022 (
            .O(N__21157),
            .I(N__21151));
    LocalMux I__2021 (
            .O(N__21154),
            .I(N__21148));
    LocalMux I__2020 (
            .O(N__21151),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4 ));
    Odrv4 I__2019 (
            .O(N__21148),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4 ));
    InMux I__2018 (
            .O(N__21143),
            .I(N__21140));
    LocalMux I__2017 (
            .O(N__21140),
            .I(N__21136));
    InMux I__2016 (
            .O(N__21139),
            .I(N__21133));
    Span4Mux_h I__2015 (
            .O(N__21136),
            .I(N__21130));
    LocalMux I__2014 (
            .O(N__21133),
            .I(N__21127));
    Odrv4 I__2013 (
            .O(N__21130),
            .I(\spi_master_inst.sclk_gen_u0.N_1737 ));
    Odrv12 I__2012 (
            .O(N__21127),
            .I(\spi_master_inst.sclk_gen_u0.N_1737 ));
    InMux I__2011 (
            .O(N__21122),
            .I(N__21119));
    LocalMux I__2010 (
            .O(N__21119),
            .I(N__21116));
    Span4Mux_h I__2009 (
            .O(N__21116),
            .I(N__21113));
    Odrv4 I__2008 (
            .O(N__21113),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4 ));
    CascadeMux I__2007 (
            .O(N__21110),
            .I(\spi_master_inst.sclk_gen_u0.N_1737_cascade_ ));
    InMux I__2006 (
            .O(N__21107),
            .I(N__21104));
    LocalMux I__2005 (
            .O(N__21104),
            .I(N__21100));
    InMux I__2004 (
            .O(N__21103),
            .I(N__21097));
    Span4Mux_h I__2003 (
            .O(N__21100),
            .I(N__21094));
    LocalMux I__2002 (
            .O(N__21097),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0 ));
    Odrv4 I__2001 (
            .O(N__21094),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0 ));
    InMux I__2000 (
            .O(N__21089),
            .I(N__21083));
    InMux I__1999 (
            .O(N__21088),
            .I(N__21083));
    LocalMux I__1998 (
            .O(N__21083),
            .I(N__21080));
    Odrv12 I__1997 (
            .O(N__21080),
            .I(\spi_master_inst.sclk_gen_u0.N_1540 ));
    InMux I__1996 (
            .O(N__21077),
            .I(N__21073));
    InMux I__1995 (
            .O(N__21076),
            .I(N__21070));
    LocalMux I__1994 (
            .O(N__21073),
            .I(N__21067));
    LocalMux I__1993 (
            .O(N__21070),
            .I(N__21059));
    Span12Mux_s8_h I__1992 (
            .O(N__21067),
            .I(N__21059));
    InMux I__1991 (
            .O(N__21066),
            .I(N__21056));
    InMux I__1990 (
            .O(N__21065),
            .I(N__21051));
    InMux I__1989 (
            .O(N__21064),
            .I(N__21051));
    Odrv12 I__1988 (
            .O(N__21059),
            .I(\spi_master_inst.ss_start_i ));
    LocalMux I__1987 (
            .O(N__21056),
            .I(\spi_master_inst.ss_start_i ));
    LocalMux I__1986 (
            .O(N__21051),
            .I(\spi_master_inst.ss_start_i ));
    CascadeMux I__1985 (
            .O(N__21044),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_ ));
    CascadeMux I__1984 (
            .O(N__21041),
            .I(\spi_master_inst.spi_data_path_u1.N_1421_cascade_ ));
    InMux I__1983 (
            .O(N__21038),
            .I(N__21035));
    LocalMux I__1982 (
            .O(N__21035),
            .I(\spi_master_inst.spi_data_path_u1.N_1422 ));
    InMux I__1981 (
            .O(N__21032),
            .I(N__21029));
    LocalMux I__1980 (
            .O(N__21029),
            .I(N__21024));
    InMux I__1979 (
            .O(N__21028),
            .I(N__21021));
    InMux I__1978 (
            .O(N__21027),
            .I(N__21018));
    Odrv4 I__1977 (
            .O(N__21024),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2 ));
    LocalMux I__1976 (
            .O(N__21021),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2 ));
    LocalMux I__1975 (
            .O(N__21018),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2 ));
    InMux I__1974 (
            .O(N__21011),
            .I(N__21007));
    InMux I__1973 (
            .O(N__21010),
            .I(N__21003));
    LocalMux I__1972 (
            .O(N__21007),
            .I(N__21000));
    InMux I__1971 (
            .O(N__21006),
            .I(N__20997));
    LocalMux I__1970 (
            .O(N__21003),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5 ));
    Odrv4 I__1969 (
            .O(N__21000),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5 ));
    LocalMux I__1968 (
            .O(N__20997),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5 ));
    CascadeMux I__1967 (
            .O(N__20990),
            .I(N__20987));
    InMux I__1966 (
            .O(N__20987),
            .I(N__20984));
    LocalMux I__1965 (
            .O(N__20984),
            .I(N__20979));
    InMux I__1964 (
            .O(N__20983),
            .I(N__20976));
    InMux I__1963 (
            .O(N__20982),
            .I(N__20973));
    Odrv4 I__1962 (
            .O(N__20979),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3 ));
    LocalMux I__1961 (
            .O(N__20976),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3 ));
    LocalMux I__1960 (
            .O(N__20973),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3 ));
    InMux I__1959 (
            .O(N__20966),
            .I(N__20962));
    InMux I__1958 (
            .O(N__20965),
            .I(N__20958));
    LocalMux I__1957 (
            .O(N__20962),
            .I(N__20955));
    InMux I__1956 (
            .O(N__20961),
            .I(N__20952));
    LocalMux I__1955 (
            .O(N__20958),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4 ));
    Odrv4 I__1954 (
            .O(N__20955),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4 ));
    LocalMux I__1953 (
            .O(N__20952),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4 ));
    InMux I__1952 (
            .O(N__20945),
            .I(N__20942));
    LocalMux I__1951 (
            .O(N__20942),
            .I(\spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1 ));
    InMux I__1950 (
            .O(N__20939),
            .I(N__20936));
    LocalMux I__1949 (
            .O(N__20936),
            .I(N__20932));
    CascadeMux I__1948 (
            .O(N__20935),
            .I(N__20928));
    Span4Mux_h I__1947 (
            .O(N__20932),
            .I(N__20925));
    InMux I__1946 (
            .O(N__20931),
            .I(N__20922));
    InMux I__1945 (
            .O(N__20928),
            .I(N__20919));
    Odrv4 I__1944 (
            .O(N__20925),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7 ));
    LocalMux I__1943 (
            .O(N__20922),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7 ));
    LocalMux I__1942 (
            .O(N__20919),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7 ));
    InMux I__1941 (
            .O(N__20912),
            .I(N__20909));
    LocalMux I__1940 (
            .O(N__20909),
            .I(N__20906));
    Span4Mux_h I__1939 (
            .O(N__20906),
            .I(N__20901));
    InMux I__1938 (
            .O(N__20905),
            .I(N__20898));
    InMux I__1937 (
            .O(N__20904),
            .I(N__20895));
    Odrv4 I__1936 (
            .O(N__20901),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6 ));
    LocalMux I__1935 (
            .O(N__20898),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6 ));
    LocalMux I__1934 (
            .O(N__20895),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6 ));
    IoInMux I__1933 (
            .O(N__20888),
            .I(N__20885));
    LocalMux I__1932 (
            .O(N__20885),
            .I(N__20882));
    Span4Mux_s2_v I__1931 (
            .O(N__20882),
            .I(N__20879));
    Sp12to4 I__1930 (
            .O(N__20879),
            .I(N__20876));
    Span12Mux_s8_h I__1929 (
            .O(N__20876),
            .I(N__20872));
    InMux I__1928 (
            .O(N__20875),
            .I(N__20869));
    Odrv12 I__1927 (
            .O(N__20872),
            .I(DAC_sclk_c));
    LocalMux I__1926 (
            .O(N__20869),
            .I(DAC_sclk_c));
    CascadeMux I__1925 (
            .O(N__20864),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_cascade_ ));
    InMux I__1924 (
            .O(N__20861),
            .I(N__20857));
    InMux I__1923 (
            .O(N__20860),
            .I(N__20854));
    LocalMux I__1922 (
            .O(N__20857),
            .I(\spi_master_inst.sclk_gen_u0.N_36 ));
    LocalMux I__1921 (
            .O(N__20854),
            .I(\spi_master_inst.sclk_gen_u0.N_36 ));
    InMux I__1920 (
            .O(N__20849),
            .I(N__20846));
    LocalMux I__1919 (
            .O(N__20846),
            .I(\spi_master_inst.sclk_gen_u0.N_5 ));
    InMux I__1918 (
            .O(N__20843),
            .I(N__20839));
    InMux I__1917 (
            .O(N__20842),
            .I(N__20835));
    LocalMux I__1916 (
            .O(N__20839),
            .I(N__20832));
    InMux I__1915 (
            .O(N__20838),
            .I(N__20829));
    LocalMux I__1914 (
            .O(N__20835),
            .I(\spi_master_inst.sclk_gen_u0.N_150_0 ));
    Odrv4 I__1913 (
            .O(N__20832),
            .I(\spi_master_inst.sclk_gen_u0.N_150_0 ));
    LocalMux I__1912 (
            .O(N__20829),
            .I(\spi_master_inst.sclk_gen_u0.N_150_0 ));
    InMux I__1911 (
            .O(N__20822),
            .I(N__20819));
    LocalMux I__1910 (
            .O(N__20819),
            .I(\spi_master_inst.sclk_gen_u0.N_48 ));
    CascadeMux I__1909 (
            .O(N__20816),
            .I(\spi_master_inst.spi_data_path_u1.N_1414_cascade_ ));
    CascadeMux I__1908 (
            .O(N__20813),
            .I(\spi_master_inst.spi_data_path_u1.N_1415_cascade_ ));
    IoInMux I__1907 (
            .O(N__20810),
            .I(N__20807));
    LocalMux I__1906 (
            .O(N__20807),
            .I(N__20804));
    IoSpan4Mux I__1905 (
            .O(N__20804),
            .I(N__20801));
    Span4Mux_s3_v I__1904 (
            .O(N__20801),
            .I(N__20798));
    Span4Mux_v I__1903 (
            .O(N__20798),
            .I(N__20795));
    Odrv4 I__1902 (
            .O(N__20795),
            .I(DAC_mosi_c));
    InMux I__1901 (
            .O(N__20792),
            .I(N__20789));
    LocalMux I__1900 (
            .O(N__20789),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1 ));
    InMux I__1899 (
            .O(N__20786),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_4 ));
    InMux I__1898 (
            .O(N__20783),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_5 ));
    InMux I__1897 (
            .O(N__20780),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_6 ));
    InMux I__1896 (
            .O(N__20777),
            .I(N__20774));
    LocalMux I__1895 (
            .O(N__20774),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3 ));
    InMux I__1894 (
            .O(N__20771),
            .I(N__20766));
    InMux I__1893 (
            .O(N__20770),
            .I(N__20763));
    InMux I__1892 (
            .O(N__20769),
            .I(N__20760));
    LocalMux I__1891 (
            .O(N__20766),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3 ));
    LocalMux I__1890 (
            .O(N__20763),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3 ));
    LocalMux I__1889 (
            .O(N__20760),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3 ));
    InMux I__1888 (
            .O(N__20753),
            .I(N__20747));
    InMux I__1887 (
            .O(N__20752),
            .I(N__20744));
    InMux I__1886 (
            .O(N__20751),
            .I(N__20739));
    InMux I__1885 (
            .O(N__20750),
            .I(N__20739));
    LocalMux I__1884 (
            .O(N__20747),
            .I(\spi_master_inst.sclk_gen_u0.N_1531 ));
    LocalMux I__1883 (
            .O(N__20744),
            .I(\spi_master_inst.sclk_gen_u0.N_1531 ));
    LocalMux I__1882 (
            .O(N__20739),
            .I(\spi_master_inst.sclk_gen_u0.N_1531 ));
    InMux I__1881 (
            .O(N__20732),
            .I(N__20728));
    InMux I__1880 (
            .O(N__20731),
            .I(N__20725));
    LocalMux I__1879 (
            .O(N__20728),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_start_iZ0 ));
    LocalMux I__1878 (
            .O(N__20725),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_start_iZ0 ));
    InMux I__1877 (
            .O(N__20720),
            .I(N__20711));
    InMux I__1876 (
            .O(N__20719),
            .I(N__20711));
    InMux I__1875 (
            .O(N__20718),
            .I(N__20711));
    LocalMux I__1874 (
            .O(N__20711),
            .I(N__20703));
    InMux I__1873 (
            .O(N__20710),
            .I(N__20692));
    InMux I__1872 (
            .O(N__20709),
            .I(N__20692));
    InMux I__1871 (
            .O(N__20708),
            .I(N__20692));
    InMux I__1870 (
            .O(N__20707),
            .I(N__20692));
    InMux I__1869 (
            .O(N__20706),
            .I(N__20692));
    Odrv4 I__1868 (
            .O(N__20703),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_start_i_i ));
    LocalMux I__1867 (
            .O(N__20692),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_start_i_i ));
    InMux I__1866 (
            .O(N__20687),
            .I(N__20682));
    InMux I__1865 (
            .O(N__20686),
            .I(N__20677));
    InMux I__1864 (
            .O(N__20685),
            .I(N__20677));
    LocalMux I__1863 (
            .O(N__20682),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0 ));
    LocalMux I__1862 (
            .O(N__20677),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0 ));
    InMux I__1861 (
            .O(N__20672),
            .I(N__20667));
    InMux I__1860 (
            .O(N__20671),
            .I(N__20664));
    InMux I__1859 (
            .O(N__20670),
            .I(N__20661));
    LocalMux I__1858 (
            .O(N__20667),
            .I(N__20658));
    LocalMux I__1857 (
            .O(N__20664),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1 ));
    LocalMux I__1856 (
            .O(N__20661),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1 ));
    Odrv4 I__1855 (
            .O(N__20658),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1 ));
    CascadeMux I__1854 (
            .O(N__20651),
            .I(N__20646));
    CascadeMux I__1853 (
            .O(N__20650),
            .I(N__20643));
    InMux I__1852 (
            .O(N__20649),
            .I(N__20640));
    InMux I__1851 (
            .O(N__20646),
            .I(N__20637));
    InMux I__1850 (
            .O(N__20643),
            .I(N__20634));
    LocalMux I__1849 (
            .O(N__20640),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3 ));
    LocalMux I__1848 (
            .O(N__20637),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3 ));
    LocalMux I__1847 (
            .O(N__20634),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3 ));
    InMux I__1846 (
            .O(N__20627),
            .I(N__20622));
    InMux I__1845 (
            .O(N__20626),
            .I(N__20619));
    InMux I__1844 (
            .O(N__20625),
            .I(N__20616));
    LocalMux I__1843 (
            .O(N__20622),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2 ));
    LocalMux I__1842 (
            .O(N__20619),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2 ));
    LocalMux I__1841 (
            .O(N__20616),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2 ));
    CascadeMux I__1840 (
            .O(N__20609),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_ ));
    CascadeMux I__1839 (
            .O(N__20606),
            .I(\spi_master_inst.sclk_gen_u0.N_48_cascade_ ));
    InMux I__1838 (
            .O(N__20603),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6 ));
    InMux I__1837 (
            .O(N__20600),
            .I(N__20597));
    LocalMux I__1836 (
            .O(N__20597),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_s_1 ));
    InMux I__1835 (
            .O(N__20594),
            .I(N__20590));
    InMux I__1834 (
            .O(N__20593),
            .I(N__20587));
    LocalMux I__1833 (
            .O(N__20590),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1 ));
    LocalMux I__1832 (
            .O(N__20587),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1 ));
    CascadeMux I__1831 (
            .O(N__20582),
            .I(N__20579));
    InMux I__1830 (
            .O(N__20579),
            .I(N__20572));
    InMux I__1829 (
            .O(N__20578),
            .I(N__20572));
    InMux I__1828 (
            .O(N__20577),
            .I(N__20568));
    LocalMux I__1827 (
            .O(N__20572),
            .I(N__20565));
    InMux I__1826 (
            .O(N__20571),
            .I(N__20562));
    LocalMux I__1825 (
            .O(N__20568),
            .I(N__20559));
    Odrv4 I__1824 (
            .O(N__20565),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0 ));
    LocalMux I__1823 (
            .O(N__20562),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0 ));
    Odrv12 I__1822 (
            .O(N__20559),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0 ));
    InMux I__1821 (
            .O(N__20552),
            .I(N__20549));
    LocalMux I__1820 (
            .O(N__20549),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_s_0 ));
    CascadeMux I__1819 (
            .O(N__20546),
            .I(N__20542));
    InMux I__1818 (
            .O(N__20545),
            .I(N__20533));
    InMux I__1817 (
            .O(N__20542),
            .I(N__20530));
    InMux I__1816 (
            .O(N__20541),
            .I(N__20523));
    InMux I__1815 (
            .O(N__20540),
            .I(N__20523));
    InMux I__1814 (
            .O(N__20539),
            .I(N__20523));
    InMux I__1813 (
            .O(N__20538),
            .I(N__20516));
    InMux I__1812 (
            .O(N__20537),
            .I(N__20516));
    InMux I__1811 (
            .O(N__20536),
            .I(N__20516));
    LocalMux I__1810 (
            .O(N__20533),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i ));
    LocalMux I__1809 (
            .O(N__20530),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i ));
    LocalMux I__1808 (
            .O(N__20523),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i ));
    LocalMux I__1807 (
            .O(N__20516),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i ));
    InMux I__1806 (
            .O(N__20507),
            .I(N__20500));
    InMux I__1805 (
            .O(N__20506),
            .I(N__20500));
    InMux I__1804 (
            .O(N__20505),
            .I(N__20497));
    LocalMux I__1803 (
            .O(N__20500),
            .I(\spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i ));
    LocalMux I__1802 (
            .O(N__20497),
            .I(\spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i ));
    InMux I__1801 (
            .O(N__20492),
            .I(N__20489));
    LocalMux I__1800 (
            .O(N__20489),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0 ));
    InMux I__1799 (
            .O(N__20486),
            .I(bfn_3_8_0_));
    InMux I__1798 (
            .O(N__20483),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_0 ));
    InMux I__1797 (
            .O(N__20480),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_1 ));
    InMux I__1796 (
            .O(N__20477),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_2 ));
    InMux I__1795 (
            .O(N__20474),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_3 ));
    IoInMux I__1794 (
            .O(N__20471),
            .I(N__20468));
    LocalMux I__1793 (
            .O(N__20468),
            .I(N__20465));
    Span4Mux_s3_v I__1792 (
            .O(N__20465),
            .I(N__20462));
    Span4Mux_h I__1791 (
            .O(N__20462),
            .I(N__20459));
    Odrv4 I__1790 (
            .O(N__20459),
            .I(DAC_cs_c));
    InMux I__1789 (
            .O(N__20456),
            .I(bfn_3_6_0_));
    InMux I__1788 (
            .O(N__20453),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0 ));
    InMux I__1787 (
            .O(N__20450),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1 ));
    InMux I__1786 (
            .O(N__20447),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2 ));
    InMux I__1785 (
            .O(N__20444),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3 ));
    InMux I__1784 (
            .O(N__20441),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4 ));
    InMux I__1783 (
            .O(N__20438),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5 ));
    CascadeMux I__1782 (
            .O(N__20435),
            .I(\spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1_cascade_ ));
    CascadeMux I__1781 (
            .O(N__20432),
            .I(\spi_master_inst.sclk_gen_u0.N_1531_cascade_ ));
    CascadeMux I__1780 (
            .O(N__20429),
            .I(N__20426));
    InMux I__1779 (
            .O(N__20426),
            .I(N__20417));
    InMux I__1778 (
            .O(N__20425),
            .I(N__20417));
    InMux I__1777 (
            .O(N__20424),
            .I(N__20417));
    LocalMux I__1776 (
            .O(N__20417),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1 ));
    InMux I__1775 (
            .O(N__20414),
            .I(N__20411));
    LocalMux I__1774 (
            .O(N__20411),
            .I(N__20408));
    Span12Mux_h I__1773 (
            .O(N__20408),
            .I(N__20405));
    Span12Mux_v I__1772 (
            .O(N__20405),
            .I(N__20402));
    Odrv12 I__1771 (
            .O(N__20402),
            .I(button_mode_c));
    IoInMux I__1770 (
            .O(N__20399),
            .I(N__20396));
    LocalMux I__1769 (
            .O(N__20396),
            .I(N__20393));
    Odrv12 I__1768 (
            .O(N__20393),
            .I(button_mode_ibuf_RNIN5KZ0Z7));
    InMux I__1767 (
            .O(N__20390),
            .I(sRAM_pointer_write_cry_10));
    InMux I__1766 (
            .O(N__20387),
            .I(sRAM_pointer_write_cry_11));
    InMux I__1765 (
            .O(N__20384),
            .I(sRAM_pointer_write_cry_12));
    InMux I__1764 (
            .O(N__20381),
            .I(sRAM_pointer_write_cry_13));
    InMux I__1763 (
            .O(N__20378),
            .I(sRAM_pointer_write_cry_14));
    InMux I__1762 (
            .O(N__20375),
            .I(bfn_1_13_0_));
    InMux I__1761 (
            .O(N__20372),
            .I(sRAM_pointer_write_cry_16));
    InMux I__1760 (
            .O(N__20369),
            .I(sRAM_pointer_write_cry_17));
    CEMux I__1759 (
            .O(N__20366),
            .I(N__20357));
    CEMux I__1758 (
            .O(N__20365),
            .I(N__20357));
    CEMux I__1757 (
            .O(N__20364),
            .I(N__20357));
    GlobalMux I__1756 (
            .O(N__20357),
            .I(N__20354));
    gio2CtrlBuf I__1755 (
            .O(N__20354),
            .I(N_1487_g));
    InMux I__1754 (
            .O(N__20351),
            .I(sRAM_pointer_write_cry_1));
    InMux I__1753 (
            .O(N__20348),
            .I(sRAM_pointer_write_cry_2));
    InMux I__1752 (
            .O(N__20345),
            .I(sRAM_pointer_write_cry_3));
    InMux I__1751 (
            .O(N__20342),
            .I(sRAM_pointer_write_cry_4));
    InMux I__1750 (
            .O(N__20339),
            .I(sRAM_pointer_write_cry_5));
    InMux I__1749 (
            .O(N__20336),
            .I(sRAM_pointer_write_cry_6));
    InMux I__1748 (
            .O(N__20333),
            .I(bfn_1_12_0_));
    InMux I__1747 (
            .O(N__20330),
            .I(sRAM_pointer_write_cry_8));
    InMux I__1746 (
            .O(N__20327),
            .I(sRAM_pointer_write_cry_9));
    InMux I__1745 (
            .O(N__20324),
            .I(bfn_1_11_0_));
    InMux I__1744 (
            .O(N__20321),
            .I(sRAM_pointer_write_cry_0));
    IoInMux I__1743 (
            .O(N__20318),
            .I(N__20315));
    LocalMux I__1742 (
            .O(N__20315),
            .I(N__20312));
    Span4Mux_s0_h I__1741 (
            .O(N__20312),
            .I(N__20309));
    Span4Mux_h I__1740 (
            .O(N__20309),
            .I(N__20306));
    Sp12to4 I__1739 (
            .O(N__20306),
            .I(N__20303));
    Span12Mux_v I__1738 (
            .O(N__20303),
            .I(N__20300));
    Span12Mux_h I__1737 (
            .O(N__20300),
            .I(N__20297));
    Odrv12 I__1736 (
            .O(N__20297),
            .I(\pll128M2_inst.pll_clk128 ));
    IoInMux I__1735 (
            .O(N__20294),
            .I(N__20291));
    LocalMux I__1734 (
            .O(N__20291),
            .I(N__20288));
    Span4Mux_s2_h I__1733 (
            .O(N__20288),
            .I(N__20285));
    Span4Mux_v I__1732 (
            .O(N__20285),
            .I(N__20282));
    Sp12to4 I__1731 (
            .O(N__20282),
            .I(N__20279));
    Span12Mux_s11_h I__1730 (
            .O(N__20279),
            .I(N__20276));
    Span12Mux_h I__1729 (
            .O(N__20276),
            .I(N__20273));
    Odrv12 I__1728 (
            .O(N__20273),
            .I(cs_rpi2flash_c));
    IoInMux I__1727 (
            .O(N__20270),
            .I(N__20267));
    LocalMux I__1726 (
            .O(N__20267),
            .I(N__20264));
    Span4Mux_s3_v I__1725 (
            .O(N__20264),
            .I(N__20261));
    Sp12to4 I__1724 (
            .O(N__20261),
            .I(N__20258));
    Span12Mux_h I__1723 (
            .O(N__20258),
            .I(N__20255));
    Span12Mux_v I__1722 (
            .O(N__20255),
            .I(N__20252));
    Odrv12 I__1721 (
            .O(N__20252),
            .I(clk_c));
    IoInMux I__1720 (
            .O(N__20249),
            .I(N__20246));
    LocalMux I__1719 (
            .O(N__20246),
            .I(N__20243));
    Odrv4 I__1718 (
            .O(N__20243),
            .I(\pll128M2_inst.pll_clk64_0 ));
    INV \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C  (
            .O(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .I(N__48262));
    INV \INVspi_slave_inst.rx_done_neg_sclk_iC  (
            .O(\INVspi_slave_inst.rx_done_neg_sclk_iC_net ),
            .I(N__48265));
    INV \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C  (
            .O(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .I(N__48261));
    defparam IN_MUX_bfv_6_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_12_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(un8_trig_prev_0_cry_7),
            .carryinitout(bfn_6_13_0_));
    defparam IN_MUX_bfv_20_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_10_0_));
    defparam IN_MUX_bfv_20_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_11_0_ (
            .carryinitin(un2_scounterdac_cry_8),
            .carryinitout(bfn_20_11_0_));
    defparam IN_MUX_bfv_13_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_14_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(un1_sacqtime_cry_7),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(un1_sacqtime_cry_15),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(un1_sacqtime_cry_23),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_16_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_14_0_ (
            .carryinitin(un1_button_debounce_counter_cry_8),
            .carryinitout(bfn_16_14_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(un1_button_debounce_counter_cry_16),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO ),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(un7_spon_cry_7),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(un7_spon_cry_15),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(un7_spon_cry_23),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(un5_sdacdyn_cry_7),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(un5_sdacdyn_cry_15),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(un5_sdacdyn_cry_23),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(un4_spoff_cry_7),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(un4_spoff_cry_15),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(un4_spoff_cry_23),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(un4_speriod_cry_7),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(un4_speriod_cry_15),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(un4_speriod_cry_23),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(un4_sacqtime_cry_7),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(un4_sacqtime_cry_15),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(un4_sacqtime_cry_23),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(un1_spoff_cry_7),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(un1_spoff_cry_15),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(un1_spoff_cry_23),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(un10_trig_prev_cry_7),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(un10_trig_prev_cry_15),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_22_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_7_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_3_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_6_0_));
    defparam IN_MUX_bfv_3_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_8_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(un1_sTrigCounter_cry_7),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(sRAM_pointer_write_cry_7),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(sRAM_pointer_write_cry_15),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(sRAM_pointer_read_cry_7),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(sRAM_pointer_read_cry_15),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(sCounter_cry_7),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(sCounter_cry_15),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_15_0_));
    ICE_GB reset_rpi_ibuf_RNIIUT3_0 (
            .USERSIGNALTOGLOBALBUFFER(N__24725),
            .GLOBALBUFFEROUTPUT(LED3_c_i_g));
    ICE_GB un4_sacqtime_cry_23_c_RNI2CQM_0 (
            .USERSIGNALTOGLOBALBUFFER(N__26744),
            .GLOBALBUFFEROUTPUT(N_1487_g));
    ICE_GB \pll128M2_inst.PLLOUTCOREB_derived_clock_RNI5L14  (
            .USERSIGNALTOGLOBALBUFFER(N__20249),
            .GLOBALBUFFEROUTPUT(pll_clk64_0_g));
    ICE_GB spi_sclk_inferred_clock_RNIH8F3 (
            .USERSIGNALTOGLOBALBUFFER(N__25799),
            .GLOBALBUFFEROUTPUT(spi_sclk_g));
    ICE_GB sSPI_MSB0LSB1_RNILL2C1_0 (
            .USERSIGNALTOGLOBALBUFFER(N__39191),
            .GLOBALBUFFEROUTPUT(N_28_g));
    ICE_GB sCounterDAC_RNIBR1C_0_5 (
            .USERSIGNALTOGLOBALBUFFER(N__48179),
            .GLOBALBUFFEROUTPUT(op_eq_scounterdac10_g));
    ICE_GB \pll128M2_inst.PLLOUTCOREA_derived_clock_RNI4765  (
            .USERSIGNALTOGLOBALBUFFER(N__20318),
            .GLOBALBUFFEROUTPUT(pll_clk128_g));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB button_mode_ibuf_RNIN5K7_0 (
            .USERSIGNALTOGLOBALBUFFER(N__20399),
            .GLOBALBUFFEROUTPUT(N_3154_g));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam sRAM_pointer_write_0_LC_1_11_0.C_ON=1'b1;
    defparam sRAM_pointer_write_0_LC_1_11_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_0_LC_1_11_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_0_LC_1_11_0 (
            .in0(N__39407),
            .in1(N__35872),
            .in2(_gnd_net_),
            .in3(N__20324),
            .lcout(sRAM_pointer_writeZ0Z_0),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(sRAM_pointer_write_cry_0),
            .clk(N__52346),
            .ce(N__20364),
            .sr(N__51801));
    defparam sRAM_pointer_write_1_LC_1_11_1.C_ON=1'b1;
    defparam sRAM_pointer_write_1_LC_1_11_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_1_LC_1_11_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_1_LC_1_11_1 (
            .in0(N__39399),
            .in1(N__36058),
            .in2(_gnd_net_),
            .in3(N__20321),
            .lcout(sRAM_pointer_writeZ0Z_1),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_0),
            .carryout(sRAM_pointer_write_cry_1),
            .clk(N__52346),
            .ce(N__20364),
            .sr(N__51801));
    defparam sRAM_pointer_write_2_LC_1_11_2.C_ON=1'b1;
    defparam sRAM_pointer_write_2_LC_1_11_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_2_LC_1_11_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_2_LC_1_11_2 (
            .in0(N__39408),
            .in1(N__36100),
            .in2(_gnd_net_),
            .in3(N__20351),
            .lcout(sRAM_pointer_writeZ0Z_2),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_1),
            .carryout(sRAM_pointer_write_cry_2),
            .clk(N__52346),
            .ce(N__20364),
            .sr(N__51801));
    defparam sRAM_pointer_write_3_LC_1_11_3.C_ON=1'b1;
    defparam sRAM_pointer_write_3_LC_1_11_3.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_3_LC_1_11_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_3_LC_1_11_3 (
            .in0(N__39400),
            .in1(N__43510),
            .in2(_gnd_net_),
            .in3(N__20348),
            .lcout(sRAM_pointer_writeZ0Z_3),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_2),
            .carryout(sRAM_pointer_write_cry_3),
            .clk(N__52346),
            .ce(N__20364),
            .sr(N__51801));
    defparam sRAM_pointer_write_4_LC_1_11_4.C_ON=1'b1;
    defparam sRAM_pointer_write_4_LC_1_11_4.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_4_LC_1_11_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_4_LC_1_11_4 (
            .in0(N__39409),
            .in1(N__43573),
            .in2(_gnd_net_),
            .in3(N__20345),
            .lcout(sRAM_pointer_writeZ0Z_4),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_3),
            .carryout(sRAM_pointer_write_cry_4),
            .clk(N__52346),
            .ce(N__20364),
            .sr(N__51801));
    defparam sRAM_pointer_write_5_LC_1_11_5.C_ON=1'b1;
    defparam sRAM_pointer_write_5_LC_1_11_5.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_5_LC_1_11_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_5_LC_1_11_5 (
            .in0(N__39401),
            .in1(N__35227),
            .in2(_gnd_net_),
            .in3(N__20342),
            .lcout(sRAM_pointer_writeZ0Z_5),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_4),
            .carryout(sRAM_pointer_write_cry_5),
            .clk(N__52346),
            .ce(N__20364),
            .sr(N__51801));
    defparam sRAM_pointer_write_6_LC_1_11_6.C_ON=1'b1;
    defparam sRAM_pointer_write_6_LC_1_11_6.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_6_LC_1_11_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_6_LC_1_11_6 (
            .in0(N__39410),
            .in1(N__36001),
            .in2(_gnd_net_),
            .in3(N__20339),
            .lcout(sRAM_pointer_writeZ0Z_6),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_5),
            .carryout(sRAM_pointer_write_cry_6),
            .clk(N__52346),
            .ce(N__20364),
            .sr(N__51801));
    defparam sRAM_pointer_write_7_LC_1_11_7.C_ON=1'b1;
    defparam sRAM_pointer_write_7_LC_1_11_7.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_7_LC_1_11_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_7_LC_1_11_7 (
            .in0(N__39402),
            .in1(N__36181),
            .in2(_gnd_net_),
            .in3(N__20336),
            .lcout(sRAM_pointer_writeZ0Z_7),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_6),
            .carryout(sRAM_pointer_write_cry_7),
            .clk(N__52346),
            .ce(N__20364),
            .sr(N__51801));
    defparam sRAM_pointer_write_8_LC_1_12_0.C_ON=1'b1;
    defparam sRAM_pointer_write_8_LC_1_12_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_8_LC_1_12_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_8_LC_1_12_0 (
            .in0(N__39406),
            .in1(N__43645),
            .in2(_gnd_net_),
            .in3(N__20333),
            .lcout(sRAM_pointer_writeZ0Z_8),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(sRAM_pointer_write_cry_8),
            .clk(N__52348),
            .ce(N__20365),
            .sr(N__51788));
    defparam sRAM_pointer_write_9_LC_1_12_1.C_ON=1'b1;
    defparam sRAM_pointer_write_9_LC_1_12_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_9_LC_1_12_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_9_LC_1_12_1 (
            .in0(N__39359),
            .in1(N__36250),
            .in2(_gnd_net_),
            .in3(N__20330),
            .lcout(sRAM_pointer_writeZ0Z_9),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_8),
            .carryout(sRAM_pointer_write_cry_9),
            .clk(N__52348),
            .ce(N__20365),
            .sr(N__51788));
    defparam sRAM_pointer_write_10_LC_1_12_2.C_ON=1'b1;
    defparam sRAM_pointer_write_10_LC_1_12_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_10_LC_1_12_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_10_LC_1_12_2 (
            .in0(N__39403),
            .in1(N__35809),
            .in2(_gnd_net_),
            .in3(N__20327),
            .lcout(sRAM_pointer_writeZ0Z_10),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_9),
            .carryout(sRAM_pointer_write_cry_10),
            .clk(N__52348),
            .ce(N__20365),
            .sr(N__51788));
    defparam sRAM_pointer_write_11_LC_1_12_3.C_ON=1'b1;
    defparam sRAM_pointer_write_11_LC_1_12_3.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_11_LC_1_12_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_11_LC_1_12_3 (
            .in0(N__39356),
            .in1(N__35737),
            .in2(_gnd_net_),
            .in3(N__20390),
            .lcout(sRAM_pointer_writeZ0Z_11),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_10),
            .carryout(sRAM_pointer_write_cry_11),
            .clk(N__52348),
            .ce(N__20365),
            .sr(N__51788));
    defparam sRAM_pointer_write_12_LC_1_12_4.C_ON=1'b1;
    defparam sRAM_pointer_write_12_LC_1_12_4.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_12_LC_1_12_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_12_LC_1_12_4 (
            .in0(N__39404),
            .in1(N__35689),
            .in2(_gnd_net_),
            .in3(N__20387),
            .lcout(sRAM_pointer_writeZ0Z_12),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_11),
            .carryout(sRAM_pointer_write_cry_12),
            .clk(N__52348),
            .ce(N__20365),
            .sr(N__51788));
    defparam sRAM_pointer_write_13_LC_1_12_5.C_ON=1'b1;
    defparam sRAM_pointer_write_13_LC_1_12_5.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_13_LC_1_12_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_13_LC_1_12_5 (
            .in0(N__39357),
            .in1(N__35605),
            .in2(_gnd_net_),
            .in3(N__20384),
            .lcout(sRAM_pointer_writeZ0Z_13),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_12),
            .carryout(sRAM_pointer_write_cry_13),
            .clk(N__52348),
            .ce(N__20365),
            .sr(N__51788));
    defparam sRAM_pointer_write_14_LC_1_12_6.C_ON=1'b1;
    defparam sRAM_pointer_write_14_LC_1_12_6.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_14_LC_1_12_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_14_LC_1_12_6 (
            .in0(N__39405),
            .in1(N__35560),
            .in2(_gnd_net_),
            .in3(N__20381),
            .lcout(sRAM_pointer_writeZ0Z_14),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_13),
            .carryout(sRAM_pointer_write_cry_14),
            .clk(N__52348),
            .ce(N__20365),
            .sr(N__51788));
    defparam sRAM_pointer_write_15_LC_1_12_7.C_ON=1'b1;
    defparam sRAM_pointer_write_15_LC_1_12_7.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_15_LC_1_12_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_15_LC_1_12_7 (
            .in0(N__39358),
            .in1(N__35464),
            .in2(_gnd_net_),
            .in3(N__20378),
            .lcout(sRAM_pointer_writeZ0Z_15),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_14),
            .carryout(sRAM_pointer_write_cry_15),
            .clk(N__52348),
            .ce(N__20365),
            .sr(N__51788));
    defparam sRAM_pointer_write_16_LC_1_13_0.C_ON=1'b1;
    defparam sRAM_pointer_write_16_LC_1_13_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_16_LC_1_13_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_16_LC_1_13_0 (
            .in0(N__39397),
            .in1(N__35395),
            .in2(_gnd_net_),
            .in3(N__20375),
            .lcout(sRAM_pointer_writeZ0Z_16),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(sRAM_pointer_write_cry_16),
            .clk(N__52349),
            .ce(N__20366),
            .sr(N__51776));
    defparam sRAM_pointer_write_17_LC_1_13_1.C_ON=1'b1;
    defparam sRAM_pointer_write_17_LC_1_13_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_17_LC_1_13_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_17_LC_1_13_1 (
            .in0(N__39396),
            .in1(N__36388),
            .in2(_gnd_net_),
            .in3(N__20372),
            .lcout(sRAM_pointer_writeZ0Z_17),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_16),
            .carryout(sRAM_pointer_write_cry_17),
            .clk(N__52349),
            .ce(N__20366),
            .sr(N__51776));
    defparam sRAM_pointer_write_18_LC_1_13_2.C_ON=1'b0;
    defparam sRAM_pointer_write_18_LC_1_13_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_18_LC_1_13_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_18_LC_1_13_2 (
            .in0(N__39398),
            .in1(N__36322),
            .in2(_gnd_net_),
            .in3(N__20369),
            .lcout(sRAM_pointer_writeZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52349),
            .ce(N__20366),
            .sr(N__51776));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_RNIPPNJ2_LC_2_6_1 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_RNIPPNJ2_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_RNIPPNJ2_LC_2_6_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_start_i_RNIPPNJ2_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__20577),
            .in2(_gnd_net_),
            .in3(N__20505),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIIUTC1_7_LC_2_6_6 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIIUTC1_7_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIIUTC1_7_LC_2_6_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIIUTC1_7_LC_2_6_6  (
            .in0(N__20904),
            .in1(N__21006),
            .in2(N__20935),
            .in3(N__20961),
            .lcout(),
            .ltout(\spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIL2KE2_1_LC_2_6_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIL2KE2_1_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIL2KE2_1_LC_2_6_7 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIL2KE2_1_LC_2_6_7  (
            .in0(N__21027),
            .in1(N__20982),
            .in2(N__20435),
            .in3(N__20593),
            .lcout(\spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4D3E3_1_LC_2_8_1 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4D3E3_1_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4D3E3_1_LC_2_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4D3E3_1_LC_2_8_1  (
            .in0(N__20672),
            .in1(N__20777),
            .in2(N__20650),
            .in3(N__21139),
            .lcout(\spi_master_inst.sclk_gen_u0.N_1531 ),
            .ltout(\spi_master_inst.sclk_gen_u0.N_1531_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0RFT3_1_LC_2_8_2 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0RFT3_1_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0RFT3_1_LC_2_8_2 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0RFT3_1_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__20769),
            .in2(N__20432),
            .in3(N__20424),
            .lcout(\spi_master_inst.sclk_gen_u0.N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_1_LC_2_8_5 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_1_LC_2_8_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_1_LC_2_8_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_1_LC_2_8_5  (
            .in0(N__20751),
            .in1(N__24378),
            .in2(N__20429),
            .in3(N__24551),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48488),
            .ce(),
            .sr(N__51818));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI1JPL3_1_LC_2_8_6 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI1JPL3_1_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI1JPL3_1_LC_2_8_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI1JPL3_1_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(N__20425),
            .in2(_gnd_net_),
            .in3(N__20750),
            .lcout(\spi_master_inst.sclk_gen_u0.N_1540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_LC_2_9_4 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_LC_2_9_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_LC_2_9_4 .LUT_INIT=16'b0010000011101111;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_start_i_LC_2_9_4  (
            .in0(N__20732),
            .in1(N__24550),
            .in2(N__24387),
            .in3(N__20849),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_start_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48489),
            .ce(),
            .sr(N__51810));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_3_LC_2_9_6 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_3_LC_2_9_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_3_LC_2_9_6 .LUT_INIT=16'b1010110010100000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_3_LC_2_9_6  (
            .in0(N__24460),
            .in1(N__20753),
            .in2(N__24513),
            .in3(N__20771),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48489),
            .ce(),
            .sr(N__51810));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_LC_2_9_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_LC_2_9_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_LC_2_9_7 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_start_i_LC_2_9_7  (
            .in0(N__20571),
            .in1(N__20842),
            .in2(N__24512),
            .in3(N__20861),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48489),
            .ce(),
            .sr(N__51810));
    defparam button_mode_ibuf_RNIN5K7_LC_2_10_5.C_ON=1'b0;
    defparam button_mode_ibuf_RNIN5K7_LC_2_10_5.SEQ_MODE=4'b0000;
    defparam button_mode_ibuf_RNIN5K7_LC_2_10_5.LUT_INIT=16'b0101010100000000;
    LogicCell40 button_mode_ibuf_RNIN5K7_LC_2_10_5 (
            .in0(N__20414),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49445),
            .lcout(button_mode_ibuf_RNIN5KZ0Z7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_12_7_LC_2_11_0.C_ON=1'b0;
    defparam sDAC_mem_12_7_LC_2_11_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_7_LC_2_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_7_LC_2_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50027),
            .lcout(sDAC_mem_12Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52341),
            .ce(N__36959),
            .sr(N__51789));
    defparam \spi_master_inst.o_slave_csn_0_LC_3_1_1 .C_ON=1'b0;
    defparam \spi_master_inst.o_slave_csn_0_LC_3_1_1 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.o_slave_csn_0_LC_3_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.o_slave_csn_0_LC_3_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21077),
            .lcout(DAC_cs_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48464),
            .ce(),
            .sr(N__51827));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_0_LC_3_6_0 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_0_LC_3_6_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_0_LC_3_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_0_LC_3_6_0  (
            .in0(_gnd_net_),
            .in1(N__20492),
            .in2(_gnd_net_),
            .in3(N__20456),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_i_s_0 ),
            .ltout(),
            .carryin(bfn_3_6_0_),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_1_LC_3_6_1 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_1_LC_3_6_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_1_LC_3_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_1_LC_3_6_1  (
            .in0(_gnd_net_),
            .in1(N__20594),
            .in2(_gnd_net_),
            .in3(N__20453),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_i_s_1 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_2_LC_3_6_2 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_2_LC_3_6_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_2_LC_3_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_2_LC_3_6_2  (
            .in0(N__20536),
            .in1(N__21028),
            .in2(_gnd_net_),
            .in3(N__20450),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2 ),
            .clk(N__48478),
            .ce(),
            .sr(N__51822));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_3_LC_3_6_3 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_3_LC_3_6_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_3_LC_3_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_3_LC_3_6_3  (
            .in0(N__20539),
            .in1(N__20983),
            .in2(_gnd_net_),
            .in3(N__20447),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3 ),
            .clk(N__48478),
            .ce(),
            .sr(N__51822));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_4_LC_3_6_4 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_4_LC_3_6_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_4_LC_3_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_4_LC_3_6_4  (
            .in0(N__20537),
            .in1(N__20965),
            .in2(_gnd_net_),
            .in3(N__20444),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4 ),
            .clk(N__48478),
            .ce(),
            .sr(N__51822));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_5_LC_3_6_5 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_5_LC_3_6_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_5_LC_3_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_5_LC_3_6_5  (
            .in0(N__20540),
            .in1(N__21010),
            .in2(_gnd_net_),
            .in3(N__20441),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5 ),
            .clk(N__48478),
            .ce(),
            .sr(N__51822));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_6_LC_3_6_6 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_6_LC_3_6_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_6_LC_3_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_6_LC_3_6_6  (
            .in0(N__20538),
            .in1(N__20905),
            .in2(_gnd_net_),
            .in3(N__20438),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6 ),
            .clk(N__48478),
            .ce(),
            .sr(N__51822));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_7_LC_3_6_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_7_LC_3_6_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_7_LC_3_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_7_LC_3_6_7  (
            .in0(N__20541),
            .in1(N__20931),
            .in2(_gnd_net_),
            .in3(N__20603),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48478),
            .ce(),
            .sr(N__51822));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_1_LC_3_7_2 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_1_LC_3_7_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_1_LC_3_7_2 .LUT_INIT=16'b1100111110101010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_1_LC_3_7_2  (
            .in0(N__20600),
            .in1(N__20507),
            .in2(N__20582),
            .in3(N__20545),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48482),
            .ce(),
            .sr(N__51819));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_0_LC_3_7_4 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_0_LC_3_7_4 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_0_LC_3_7_4 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_0_LC_3_7_4  (
            .in0(N__20578),
            .in1(N__20552),
            .in2(N__20546),
            .in3(N__20506),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48482),
            .ce(),
            .sr(N__51819));
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_LC_3_7_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_LC_3_7_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_LC_3_7_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.falling_count_start_i_LC_3_7_7  (
            .in0(N__27943),
            .in1(N__24332),
            .in2(_gnd_net_),
            .in3(N__20843),
            .lcout(\spi_master_inst.sclk_gen_u0.falling_count_start_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48482),
            .ce(),
            .sr(N__51819));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_0_LC_3_8_0 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_0_LC_3_8_0 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_0_LC_3_8_0 .LUT_INIT=16'b1011101111101110;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_0_LC_3_8_0  (
            .in0(N__20706),
            .in1(N__20687),
            .in2(_gnd_net_),
            .in3(N__20486),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0 ),
            .ltout(),
            .carryin(bfn_3_8_0_),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_0 ),
            .clk(N__48485),
            .ce(),
            .sr(N__51811));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_1_LC_3_8_1 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_1_LC_3_8_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_1_LC_3_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_1_LC_3_8_1  (
            .in0(N__20718),
            .in1(N__20671),
            .in2(_gnd_net_),
            .in3(N__20483),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_0 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_1 ),
            .clk(N__48485),
            .ce(),
            .sr(N__51811));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_2_LC_3_8_2 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_2_LC_3_8_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_2_LC_3_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_2_LC_3_8_2  (
            .in0(N__20707),
            .in1(N__20627),
            .in2(_gnd_net_),
            .in3(N__20480),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_1 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_2 ),
            .clk(N__48485),
            .ce(),
            .sr(N__51811));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_3_LC_3_8_3 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_3_LC_3_8_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_3_LC_3_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_3_LC_3_8_3  (
            .in0(N__20719),
            .in1(N__20649),
            .in2(_gnd_net_),
            .in3(N__20477),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_2 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_3 ),
            .clk(N__48485),
            .ce(),
            .sr(N__51811));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_4_LC_3_8_4 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_4_LC_3_8_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_4_LC_3_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_4_LC_3_8_4  (
            .in0(N__20708),
            .in1(N__21157),
            .in2(_gnd_net_),
            .in3(N__20474),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_3 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_4 ),
            .clk(N__48485),
            .ce(),
            .sr(N__51811));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_5_LC_3_8_5 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_5_LC_3_8_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_5_LC_3_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_5_LC_3_8_5  (
            .in0(N__20720),
            .in1(N__21190),
            .in2(_gnd_net_),
            .in3(N__20786),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_4 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_5 ),
            .clk(N__48485),
            .ce(),
            .sr(N__51811));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_6_LC_3_8_6 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_6_LC_3_8_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_6_LC_3_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_6_LC_3_8_6  (
            .in0(N__20709),
            .in1(N__21206),
            .in2(_gnd_net_),
            .in3(N__20783),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_5 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_6 ),
            .clk(N__48485),
            .ce(),
            .sr(N__51811));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_7_LC_3_8_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_7_LC_3_8_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_7_LC_3_8_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_7_LC_3_8_7  (
            .in0(N__21172),
            .in1(N__20710),
            .in2(_gnd_net_),
            .in3(N__20780),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48485),
            .ce(),
            .sr(N__51811));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4MGR_0_LC_3_9_0 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4MGR_0_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4MGR_0_LC_3_9_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4MGR_0_LC_3_9_0  (
            .in0(_gnd_net_),
            .in1(N__20625),
            .in2(_gnd_net_),
            .in3(N__20685),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI3LPL3_3_LC_3_9_2 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI3LPL3_3_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI3LPL3_3_LC_3_9_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI3LPL3_3_LC_3_9_2  (
            .in0(_gnd_net_),
            .in1(N__20770),
            .in2(_gnd_net_),
            .in3(N__20752),
            .lcout(\spi_master_inst.sclk_gen_u0.N_150_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNI6TQC_LC_3_9_4 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNI6TQC_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNI6TQC_LC_3_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNI6TQC_LC_3_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20731),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_start_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIAE1N1_0_LC_3_9_5 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIAE1N1_0_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIAE1N1_0_LC_3_9_5 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_RNIAE1N1_0_LC_3_9_5  (
            .in0(N__20686),
            .in1(N__20670),
            .in2(N__20651),
            .in3(N__20626),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4 ),
            .ltout(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0IPL3_0_LC_3_9_6 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0IPL3_0_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0IPL3_0_LC_3_9_6 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0IPL3_0_LC_3_9_6  (
            .in0(_gnd_net_),
            .in1(N__21107),
            .in2(N__20609),
            .in3(N__21143),
            .lcout(\spi_master_inst.sclk_gen_u0.N_48 ),
            .ltout(\spi_master_inst.sclk_gen_u0.N_48_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNO_0_LC_3_9_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNO_0_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNO_0_LC_3_9_7 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNO_0_LC_3_9_7  (
            .in0(N__24495),
            .in1(N__24459),
            .in2(N__20606),
            .in3(N__20860),
            .lcout(\spi_master_inst.sclk_gen_u0.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_2_LC_3_10_2 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_2_LC_3_10_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_2_LC_3_10_2 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_2_LC_3_10_2  (
            .in0(N__24385),
            .in1(N__24543),
            .in2(_gnd_net_),
            .in3(N__20838),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48490),
            .ce(),
            .sr(N__51790));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_4_LC_3_10_5 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_4_LC_3_10_5 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_4_LC_3_10_5 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_4_LC_3_10_5  (
            .in0(N__24499),
            .in1(N__24461),
            .in2(_gnd_net_),
            .in3(N__20822),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48490),
            .ce(),
            .sr(N__51790));
    defparam sAddress_7_LC_3_11_0.C_ON=1'b0;
    defparam sAddress_7_LC_3_11_0.SEQ_MODE=4'b1010;
    defparam sAddress_7_LC_3_11_0.LUT_INIT=16'b0101010100000000;
    LogicCell40 sAddress_7_LC_3_11_0 (
            .in0(N__26198),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49929),
            .lcout(sAddressZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52332),
            .ce(N__23423),
            .sr(N__51777));
    defparam sAddress_6_LC_3_11_3.C_ON=1'b0;
    defparam sAddress_6_LC_3_11_3.SEQ_MODE=4'b1010;
    defparam sAddress_6_LC_3_11_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 sAddress_6_LC_3_11_3 (
            .in0(_gnd_net_),
            .in1(N__50327),
            .in2(_gnd_net_),
            .in3(N__26197),
            .lcout(sAddressZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52332),
            .ce(N__23423),
            .sr(N__51777));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI73G42_2_LC_5_3_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI73G42_2_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI73G42_2_LC_5_3_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI73G42_2_LC_5_3_0  (
            .in0(N__21421),
            .in1(N__21236),
            .in2(_gnd_net_),
            .in3(N__20792),
            .lcout(),
            .ltout(\spi_master_inst.spi_data_path_u1.N_1414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI60IB4_1_LC_5_3_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI60IB4_1_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI60IB4_1_LC_5_3_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI60IB4_1_LC_5_3_1  (
            .in0(N__21512),
            .in1(_gnd_net_),
            .in2(N__20816),
            .in3(N__21242),
            .lcout(),
            .ltout(\spi_master_inst.spi_data_path_u1.N_1415_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI70MD9_0_LC_5_3_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI70MD9_0_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI70MD9_0_LC_5_3_2 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI70MD9_0_LC_5_3_2  (
            .in0(N__21578),
            .in1(N__21038),
            .in2(N__20813),
            .in3(N__21076),
            .lcout(DAC_mosi_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01_1_LC_5_3_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01_1_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01_1_LC_5_3_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01_1_LC_5_3_7  (
            .in0(N__25748),
            .in1(N__21797),
            .in2(_gnd_net_),
            .in3(N__24668),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01_0_LC_5_4_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01_0_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01_0_LC_5_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01_0_LC_5_4_3  (
            .in0(N__47567),
            .in1(N__21767),
            .in2(_gnd_net_),
            .in3(N__24667),
            .lcout(),
            .ltout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI3VF42_2_LC_5_4_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI3VF42_2_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI3VF42_2_LC_5_4_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI3VF42_2_LC_5_4_4  (
            .in0(_gnd_net_),
            .in1(N__23228),
            .in2(N__21044),
            .in3(N__21416),
            .lcout(),
            .ltout(\spi_master_inst.spi_data_path_u1.N_1421_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIUNHB4_1_LC_5_4_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIUNHB4_1_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIUNHB4_1_LC_5_4_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIUNHB4_1_LC_5_4_5  (
            .in0(N__21224),
            .in1(_gnd_net_),
            .in2(N__21041),
            .in3(N__21511),
            .lcout(\spi_master_inst.spi_data_path_u1.N_1422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_RNIH6AC_LC_5_6_3 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_RNIH6AC_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_RNIH6AC_LC_5_6_3 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.o_sclk_RNIH6AC_LC_5_6_3  (
            .in0(N__27989),
            .in1(N__24386),
            .in2(_gnd_net_),
            .in3(N__20875),
            .lcout(\spi_master_inst.o_sclk_RNIH6AC ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_RNO_0_LC_5_6_4 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_RNO_0_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_RNO_0_LC_5_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \spi_master_inst.sclk_gen_u0.div_clk_i_RNO_0_LC_5_6_4  (
            .in0(N__21032),
            .in1(N__21011),
            .in2(N__20990),
            .in3(N__20966),
            .lcout(\spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_LC_5_7_1 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_LC_5_7_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_LC_5_7_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.div_clk_i_LC_5_7_1  (
            .in0(N__20945),
            .in1(N__20939),
            .in2(_gnd_net_),
            .in3(N__20912),
            .lcout(\spi_master_inst.sclk_gen_u0.div_clk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48474),
            .ce(),
            .sr(N__51802));
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_LC_5_7_2 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_LC_5_7_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_LC_5_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.o_sclk_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(N__27993),
            .in2(_gnd_net_),
            .in3(N__24389),
            .lcout(DAC_sclk_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48474),
            .ce(),
            .sr(N__51802));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_2_LC_5_7_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_2_LC_5_7_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_2_LC_5_7_4 .LUT_INIT=16'b0001101000101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_2_LC_5_7_4  (
            .in0(N__21401),
            .in1(N__21331),
            .in2(N__21296),
            .in3(N__21365),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48474),
            .ce(),
            .sr(N__51802));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIL1LO1_2_LC_5_7_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIL1LO1_2_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIL1LO1_2_LC_5_7_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIL1LO1_2_LC_5_7_5  (
            .in0(N__21476),
            .in1(N__21400),
            .in2(_gnd_net_),
            .in3(N__24651),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6 ),
            .ltout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_i_LC_5_7_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_i_LC_5_7_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_i_LC_5_7_6 .LUT_INIT=16'b1110101011100010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_i_LC_5_7_6  (
            .in0(N__23170),
            .in1(N__21284),
            .in2(N__20864),
            .in3(N__21066),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48474),
            .ce(),
            .sr(N__51802));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_3_LC_5_7_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_3_LC_5_7_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_3_LC_5_7_7 .LUT_INIT=16'b0100011001001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_3_LC_5_7_7  (
            .in0(N__21283),
            .in1(N__24652),
            .in2(N__21332),
            .in3(N__21356),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48474),
            .ce(),
            .sr(N__51802));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIQU1N1_7_LC_5_8_1 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIQU1N1_7_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIQU1N1_7_LC_5_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_RNIQU1N1_7_LC_5_8_1  (
            .in0(N__21205),
            .in1(N__21191),
            .in2(N__21176),
            .in3(N__21158),
            .lcout(\spi_master_inst.sclk_gen_u0.N_1737 ),
            .ltout(\spi_master_inst.sclk_gen_u0.N_1737_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_0_LC_5_8_2 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_0_LC_5_8_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_0_LC_5_8_2 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_0_LC_5_8_2  (
            .in0(N__21089),
            .in1(N__21122),
            .in2(N__21110),
            .in3(N__21103),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48479),
            .ce(),
            .sr(N__51791));
    defparam \spi_master_inst.sclk_gen_u0.o_ss_start_LC_5_8_5 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.o_ss_start_LC_5_8_5 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.sclk_gen_u0.o_ss_start_LC_5_8_5 .LUT_INIT=16'b1111111100111010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.o_ss_start_LC_5_8_5  (
            .in0(N__21065),
            .in1(N__24454),
            .in2(N__24521),
            .in3(N__21088),
            .lcout(\spi_master_inst.ss_start_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48479),
            .ce(),
            .sr(N__51791));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52_2_LC_5_8_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52_2_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52_2_LC_5_8_6 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52_2_LC_5_8_6  (
            .in0(N__24649),
            .in1(N__21064),
            .in2(N__21415),
            .in3(N__21475),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam spi_mosi_ready64_prev_e_0_LC_5_9_2.C_ON=1'b0;
    defparam spi_mosi_ready64_prev_e_0_LC_5_9_2.SEQ_MODE=4'b1000;
    defparam spi_mosi_ready64_prev_e_0_LC_5_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 spi_mosi_ready64_prev_e_0_LC_5_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22001),
            .lcout(spi_mosi_ready64_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52340),
            .ce(N__49426),
            .sr(_gnd_net_));
    defparam spi_mosi_ready64_prev2_e_0_LC_5_10_4.C_ON=1'b0;
    defparam spi_mosi_ready64_prev2_e_0_LC_5_10_4.SEQ_MODE=4'b1000;
    defparam spi_mosi_ready64_prev2_e_0_LC_5_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 spi_mosi_ready64_prev2_e_0_LC_5_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21446),
            .lcout(spi_mosi_ready64_prevZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52331),
            .ce(N__49441),
            .sr(_gnd_net_));
    defparam spi_mosi_ready64_prev3_e_0_LC_5_10_6.C_ON=1'b0;
    defparam spi_mosi_ready64_prev3_e_0_LC_5_10_6.SEQ_MODE=4'b1000;
    defparam spi_mosi_ready64_prev3_e_0_LC_5_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 spi_mosi_ready64_prev3_e_0_LC_5_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21458),
            .lcout(spi_mosi_ready64_prevZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52331),
            .ce(N__49441),
            .sr(_gnd_net_));
    defparam sSingleCont_LC_5_12_7.C_ON=1'b0;
    defparam sSingleCont_LC_5_12_7.SEQ_MODE=4'b1010;
    defparam sSingleCont_LC_5_12_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 sSingleCont_LC_5_12_7 (
            .in0(_gnd_net_),
            .in1(N__26399),
            .in2(_gnd_net_),
            .in3(N__22526),
            .lcout(LED_MODE_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48491),
            .ce(),
            .sr(N__51736));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIMGLT1_2_LC_6_3_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIMGLT1_2_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIMGLT1_2_LC_6_3_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIMGLT1_2_LC_6_3_1  (
            .in0(N__21803),
            .in1(N__24614),
            .in2(_gnd_net_),
            .in3(N__21422),
            .lcout(\spi_master_inst.spi_data_path_u1.N_1411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4Q_14_LC_6_3_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4Q_14_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4Q_14_LC_6_3_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4Q_14_LC_6_3_5  (
            .in0(N__21218),
            .in1(N__21773),
            .in2(_gnd_net_),
            .in3(N__24693),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4Q_13_LC_6_4_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4Q_13_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4Q_13_LC_6_4_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4Q_13_LC_6_4_3  (
            .in0(N__24682),
            .in1(N__21785),
            .in2(_gnd_net_),
            .in3(N__21779),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIICLT1_2_LC_6_4_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIICLT1_2_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIICLT1_2_LC_6_4_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIICLT1_2_LC_6_4_5  (
            .in0(N__21417),
            .in1(N__21230),
            .in2(_gnd_net_),
            .in3(N__23219),
            .lcout(\spi_master_inst.spi_data_path_u1.N_1418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_6_LC_6_5_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_6_LC_6_5_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_6_LC_6_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_6_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21758),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48465),
            .ce(),
            .sr(N__51803));
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_LC_6_5_3 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_LC_6_5_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_LC_6_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_clk_i_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28000),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_clk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48465),
            .ce(),
            .sr(N__51803));
    defparam sDAC_mem_29_5_LC_6_6_6.C_ON=1'b0;
    defparam sDAC_mem_29_5_LC_6_6_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_5_LC_6_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_29_5_LC_6_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44952),
            .lcout(sDAC_mem_29Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52347),
            .ce(N__23153),
            .sr(N__51792));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_c_LC_6_7_0 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_c_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_c_LC_6_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_c_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__21253),
            .in2(N__21577),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_LUT4_0_LC_6_7_1 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_LUT4_0_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_LUT4_0_LC_6_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_LUT4_0_LC_6_7_1  (
            .in0(_gnd_net_),
            .in1(N__21504),
            .in2(_gnd_net_),
            .in3(N__21209),
            .lcout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0 ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_LUT4_0_LC_6_7_2 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_LUT4_0_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_LUT4_0_LC_6_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_LUT4_0_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__21402),
            .in2(_gnd_net_),
            .in3(N__21359),
            .lcout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1 ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_LUT4_0_LC_6_7_3 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_LUT4_0_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_LUT4_0_LC_6_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_LUT4_0_LC_6_7_3  (
            .in0(_gnd_net_),
            .in1(N__24650),
            .in2(_gnd_net_),
            .in3(N__21350),
            .lcout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2 ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_4_LC_6_7_4 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_4_LC_6_7_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_4_LC_6_7_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_4_LC_6_7_4  (
            .in0(N__21282),
            .in1(N__21526),
            .in2(_gnd_net_),
            .in3(N__21347),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3 ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4 ),
            .clk(N__48467),
            .ce(),
            .sr(N__51778));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_0_LC_6_7_5 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_0_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_0_LC_6_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_0_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__52738),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4 ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_1_LC_6_7_6 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_1_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_1_LC_6_7_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_1_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__52782),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_2_LC_6_7_7 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_2_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_2_LC_6_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_2_LC_6_7_7  (
            .in0(_gnd_net_),
            .in1(N__52742),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_5_LC_6_8_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_5_LC_6_8_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_5_LC_6_8_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_5_LC_6_8_0  (
            .in0(_gnd_net_),
            .in1(N__21544),
            .in2(_gnd_net_),
            .in3(N__21344),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48471),
            .ce(N__21297),
            .sr(N__51763));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_1_LC_6_9_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_1_LC_6_9_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_1_LC_6_9_0 .LUT_INIT=16'b0001111101000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_1_LC_6_9_0  (
            .in0(N__21327),
            .in1(N__21341),
            .in2(N__21305),
            .in3(N__21503),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48475),
            .ce(),
            .sr(N__51751));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_0_LC_6_9_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_0_LC_6_9_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_0_LC_6_9_6 .LUT_INIT=16'b0001110001001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_0_LC_6_9_6  (
            .in0(N__21326),
            .in1(N__21570),
            .in2(N__21304),
            .in3(N__21254),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48475),
            .ce(),
            .sr(N__51751));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_RNI06S51_5_LC_6_10_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_RNI06S51_5_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_RNI06S51_5_LC_6_10_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_RNI06S51_5_LC_6_10_0  (
            .in0(N__21563),
            .in1(N__21545),
            .in2(N__21530),
            .in3(N__21494),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam spi_mosi_ready64_prev3_e_0_RNICM2C1_LC_6_10_3.C_ON=1'b0;
    defparam spi_mosi_ready64_prev3_e_0_RNICM2C1_LC_6_10_3.SEQ_MODE=4'b0000;
    defparam spi_mosi_ready64_prev3_e_0_RNICM2C1_LC_6_10_3.LUT_INIT=16'b0000100000000000;
    LogicCell40 spi_mosi_ready64_prev3_e_0_RNICM2C1_LC_6_10_3 (
            .in0(N__21457),
            .in1(N__21445),
            .in2(N__21434),
            .in3(N__21991),
            .lcout(spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1),
            .ltout(spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sPointer_RNI85NC1_0_LC_6_10_4.C_ON=1'b0;
    defparam sPointer_RNI85NC1_0_LC_6_10_4.SEQ_MODE=4'b0000;
    defparam sPointer_RNI85NC1_0_LC_6_10_4.LUT_INIT=16'b1111000000000000;
    LogicCell40 sPointer_RNI85NC1_0_LC_6_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21425),
            .in3(N__26098),
            .lcout(un1_spointer11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam spi_mosi_ready_prev3_RNILKER_LC_6_10_5.C_ON=1'b0;
    defparam spi_mosi_ready_prev3_RNILKER_LC_6_10_5.SEQ_MODE=4'b0000;
    defparam spi_mosi_ready_prev3_RNILKER_LC_6_10_5.LUT_INIT=16'b0000100000000000;
    LogicCell40 spi_mosi_ready_prev3_RNILKER_LC_6_10_5 (
            .in0(N__21958),
            .in1(N__21970),
            .in2(N__21947),
            .in3(N__21992),
            .lcout(spi_mosi_ready_prev3_RNILKERZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNICMDR1_5_LC_6_10_6 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNICMDR1_5_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNICMDR1_5_LC_6_10_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_RNICMDR1_5_LC_6_10_6  (
            .in0(N__22040),
            .in1(N__21844),
            .in2(N__21863),
            .in3(N__22012),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_i6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_0_LC_6_11_0.C_ON=1'b0;
    defparam sEETrigCounter_0_LC_6_11_0.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_0_LC_6_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_0_LC_6_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46324),
            .lcout(un8_trig_prev_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52302),
            .ce(N__22682),
            .sr(N__51724));
    defparam sEETrigCounter_1_LC_6_11_1.C_ON=1'b0;
    defparam sEETrigCounter_1_LC_6_11_1.SEQ_MODE=4'b1011;
    defparam sEETrigCounter_1_LC_6_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_1_LC_6_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50984),
            .lcout(sEETrigCounterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52302),
            .ce(N__22682),
            .sr(N__51724));
    defparam sEETrigCounter_2_LC_6_11_2.C_ON=1'b0;
    defparam sEETrigCounter_2_LC_6_11_2.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_2_LC_6_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_2_LC_6_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47413),
            .lcout(sEETrigCounterZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52302),
            .ce(N__22682),
            .sr(N__51724));
    defparam sEETrigCounter_3_LC_6_11_3.C_ON=1'b0;
    defparam sEETrigCounter_3_LC_6_11_3.SEQ_MODE=4'b1011;
    defparam sEETrigCounter_3_LC_6_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_3_LC_6_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46840),
            .lcout(sEETrigCounterZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52302),
            .ce(N__22682),
            .sr(N__51724));
    defparam sEETrigCounter_4_LC_6_11_4.C_ON=1'b0;
    defparam sEETrigCounter_4_LC_6_11_4.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_4_LC_6_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_4_LC_6_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45554),
            .lcout(sEETrigCounterZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52302),
            .ce(N__22682),
            .sr(N__51724));
    defparam sEETrigCounter_5_LC_6_11_5.C_ON=1'b0;
    defparam sEETrigCounter_5_LC_6_11_5.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_5_LC_6_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_5_LC_6_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45000),
            .lcout(sEETrigCounterZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52302),
            .ce(N__22682),
            .sr(N__51724));
    defparam sEETrigCounter_6_LC_6_11_6.C_ON=1'b0;
    defparam sEETrigCounter_6_LC_6_11_6.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_6_LC_6_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_6_LC_6_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50328),
            .lcout(sEETrigCounterZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52302),
            .ce(N__22682),
            .sr(N__51724));
    defparam sEETrigCounter_7_LC_6_11_7.C_ON=1'b0;
    defparam sEETrigCounter_7_LC_6_11_7.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_7_LC_6_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_7_LC_6_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50023),
            .lcout(sEETrigCounterZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52302),
            .ce(N__22682),
            .sr(N__51724));
    defparam un8_trig_prev_0_cry_0_c_LC_6_12_0.C_ON=1'b1;
    defparam un8_trig_prev_0_cry_0_c_LC_6_12_0.SEQ_MODE=4'b0000;
    defparam un8_trig_prev_0_cry_0_c_LC_6_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un8_trig_prev_0_cry_0_c_LC_6_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22145),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_12_0_),
            .carryout(un8_trig_prev_0_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_trig_prev_0_cry_0_c_RNILB0M_LC_6_12_1.C_ON=1'b1;
    defparam un8_trig_prev_0_cry_0_c_RNILB0M_LC_6_12_1.SEQ_MODE=4'b0000;
    defparam un8_trig_prev_0_cry_0_c_RNILB0M_LC_6_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un8_trig_prev_0_cry_0_c_RNILB0M_LC_6_12_1 (
            .in0(_gnd_net_),
            .in1(N__52763),
            .in2(N__21626),
            .in3(N__21617),
            .lcout(un10_trig_prev_1),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_0),
            .carryout(un8_trig_prev_0_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_trig_prev_0_cry_1_c_RNINE1M_LC_6_12_2.C_ON=1'b1;
    defparam un8_trig_prev_0_cry_1_c_RNINE1M_LC_6_12_2.SEQ_MODE=4'b0000;
    defparam un8_trig_prev_0_cry_1_c_RNINE1M_LC_6_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un8_trig_prev_0_cry_1_c_RNINE1M_LC_6_12_2 (
            .in0(_gnd_net_),
            .in1(N__52779),
            .in2(N__21614),
            .in3(N__21605),
            .lcout(un10_trig_prev_2),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_1),
            .carryout(un8_trig_prev_0_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_trig_prev_0_cry_2_c_RNIPH2M_LC_6_12_3.C_ON=1'b1;
    defparam un8_trig_prev_0_cry_2_c_RNIPH2M_LC_6_12_3.SEQ_MODE=4'b0000;
    defparam un8_trig_prev_0_cry_2_c_RNIPH2M_LC_6_12_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un8_trig_prev_0_cry_2_c_RNIPH2M_LC_6_12_3 (
            .in0(_gnd_net_),
            .in1(N__52764),
            .in2(N__21602),
            .in3(N__21593),
            .lcout(un10_trig_prev_3),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_2),
            .carryout(un8_trig_prev_0_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_trig_prev_0_cry_3_c_RNIRK3M_LC_6_12_4.C_ON=1'b1;
    defparam un8_trig_prev_0_cry_3_c_RNIRK3M_LC_6_12_4.SEQ_MODE=4'b0000;
    defparam un8_trig_prev_0_cry_3_c_RNIRK3M_LC_6_12_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 un8_trig_prev_0_cry_3_c_RNIRK3M_LC_6_12_4 (
            .in0(_gnd_net_),
            .in1(N__52780),
            .in2(N__21590),
            .in3(N__21581),
            .lcout(un10_trig_prev_4),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_3),
            .carryout(un8_trig_prev_0_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_trig_prev_0_cry_4_c_RNITN4M_LC_6_12_5.C_ON=1'b1;
    defparam un8_trig_prev_0_cry_4_c_RNITN4M_LC_6_12_5.SEQ_MODE=4'b0000;
    defparam un8_trig_prev_0_cry_4_c_RNITN4M_LC_6_12_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 un8_trig_prev_0_cry_4_c_RNITN4M_LC_6_12_5 (
            .in0(_gnd_net_),
            .in1(N__52765),
            .in2(N__21680),
            .in3(N__21671),
            .lcout(un10_trig_prev_5),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_4),
            .carryout(un8_trig_prev_0_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_trig_prev_0_cry_5_c_RNIVQ5M_LC_6_12_6.C_ON=1'b1;
    defparam un8_trig_prev_0_cry_5_c_RNIVQ5M_LC_6_12_6.SEQ_MODE=4'b0000;
    defparam un8_trig_prev_0_cry_5_c_RNIVQ5M_LC_6_12_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un8_trig_prev_0_cry_5_c_RNIVQ5M_LC_6_12_6 (
            .in0(_gnd_net_),
            .in1(N__52781),
            .in2(N__21668),
            .in3(N__21659),
            .lcout(un10_trig_prev_6),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_5),
            .carryout(un8_trig_prev_0_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_trig_prev_0_cry_6_c_RNI1U6M_LC_6_12_7.C_ON=1'b1;
    defparam un8_trig_prev_0_cry_6_c_RNI1U6M_LC_6_12_7.SEQ_MODE=4'b0000;
    defparam un8_trig_prev_0_cry_6_c_RNI1U6M_LC_6_12_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 un8_trig_prev_0_cry_6_c_RNI1U6M_LC_6_12_7 (
            .in0(_gnd_net_),
            .in1(N__52766),
            .in2(N__21656),
            .in3(N__21647),
            .lcout(un10_trig_prev_7),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_6),
            .carryout(un8_trig_prev_0_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_trig_prev_0_cry_7_c_RNI318M_LC_6_13_0.C_ON=1'b1;
    defparam un8_trig_prev_0_cry_7_c_RNI318M_LC_6_13_0.SEQ_MODE=4'b0000;
    defparam un8_trig_prev_0_cry_7_c_RNI318M_LC_6_13_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un8_trig_prev_0_cry_7_c_RNI318M_LC_6_13_0 (
            .in0(_gnd_net_),
            .in1(N__52789),
            .in2(N__21689),
            .in3(N__21644),
            .lcout(un10_trig_prev_8),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(un8_trig_prev_0_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_trig_prev_0_cry_8_c_RNI549M_LC_6_13_1.C_ON=1'b1;
    defparam un8_trig_prev_0_cry_8_c_RNI549M_LC_6_13_1.SEQ_MODE=4'b0000;
    defparam un8_trig_prev_0_cry_8_c_RNI549M_LC_6_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un8_trig_prev_0_cry_8_c_RNI549M_LC_6_13_1 (
            .in0(_gnd_net_),
            .in1(N__52769),
            .in2(N__21812),
            .in3(N__21641),
            .lcout(un10_trig_prev_9),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_8),
            .carryout(un8_trig_prev_0_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_trig_prev_0_cry_9_c_RNIEEGI_LC_6_13_2.C_ON=1'b1;
    defparam un8_trig_prev_0_cry_9_c_RNIEEGI_LC_6_13_2.SEQ_MODE=4'b0000;
    defparam un8_trig_prev_0_cry_9_c_RNIEEGI_LC_6_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un8_trig_prev_0_cry_9_c_RNIEEGI_LC_6_13_2 (
            .in0(_gnd_net_),
            .in1(N__52790),
            .in2(N__21740),
            .in3(N__21638),
            .lcout(un10_trig_prev_10),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_9),
            .carryout(un8_trig_prev_0_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNINORL_11_LC_6_13_3.C_ON=1'b1;
    defparam sEETrigCounter_RNINORL_11_LC_6_13_3.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNINORL_11_LC_6_13_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 sEETrigCounter_RNINORL_11_LC_6_13_3 (
            .in0(_gnd_net_),
            .in1(N__52767),
            .in2(N__21731),
            .in3(N__21635),
            .lcout(un10_trig_prev_11),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_10),
            .carryout(un8_trig_prev_0_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIPRSL_12_LC_6_13_4.C_ON=1'b1;
    defparam sEETrigCounter_RNIPRSL_12_LC_6_13_4.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIPRSL_12_LC_6_13_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 sEETrigCounter_RNIPRSL_12_LC_6_13_4 (
            .in0(_gnd_net_),
            .in1(N__52787),
            .in2(N__21722),
            .in3(N__21632),
            .lcout(un10_trig_prev_12),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_11),
            .carryout(un8_trig_prev_0_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIRUTL_13_LC_6_13_5.C_ON=1'b1;
    defparam sEETrigCounter_RNIRUTL_13_LC_6_13_5.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIRUTL_13_LC_6_13_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 sEETrigCounter_RNIRUTL_13_LC_6_13_5 (
            .in0(_gnd_net_),
            .in1(N__52768),
            .in2(N__21713),
            .in3(N__21629),
            .lcout(un10_trig_prev_13),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_12),
            .carryout(un8_trig_prev_0_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIT1VL_14_LC_6_13_6.C_ON=1'b1;
    defparam sEETrigCounter_RNIT1VL_14_LC_6_13_6.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIT1VL_14_LC_6_13_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 sEETrigCounter_RNIT1VL_14_LC_6_13_6 (
            .in0(_gnd_net_),
            .in1(N__52788),
            .in2(N__21704),
            .in3(N__21746),
            .lcout(un10_trig_prev_14),
            .ltout(),
            .carryin(un8_trig_prev_0_cry_13),
            .carryout(un8_trig_prev_0_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIV40M_15_LC_6_13_7.C_ON=1'b0;
    defparam sEETrigCounter_RNIV40M_15_LC_6_13_7.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIV40M_15_LC_6_13_7.LUT_INIT=16'b1100110000110011;
    LogicCell40 sEETrigCounter_RNIV40M_15_LC_6_13_7 (
            .in0(_gnd_net_),
            .in1(N__21695),
            .in2(_gnd_net_),
            .in3(N__21743),
            .lcout(un10_trig_prev_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_10_LC_6_14_0.C_ON=1'b0;
    defparam sEETrigCounter_10_LC_6_14_0.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_10_LC_6_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_10_LC_6_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47480),
            .lcout(sEETrigCounterZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52333),
            .ce(N__21932),
            .sr(N__51695));
    defparam sEETrigCounter_11_LC_6_14_1.C_ON=1'b0;
    defparam sEETrigCounter_11_LC_6_14_1.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_11_LC_6_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_11_LC_6_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46919),
            .lcout(sEETrigCounterZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52333),
            .ce(N__21932),
            .sr(N__51695));
    defparam sEETrigCounter_12_LC_6_14_2.C_ON=1'b0;
    defparam sEETrigCounter_12_LC_6_14_2.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_12_LC_6_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_12_LC_6_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45601),
            .lcout(sEETrigCounterZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52333),
            .ce(N__21932),
            .sr(N__51695));
    defparam sEETrigCounter_13_LC_6_14_3.C_ON=1'b0;
    defparam sEETrigCounter_13_LC_6_14_3.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_13_LC_6_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_13_LC_6_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45117),
            .lcout(sEETrigCounterZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52333),
            .ce(N__21932),
            .sr(N__51695));
    defparam sEETrigCounter_14_LC_6_14_4.C_ON=1'b0;
    defparam sEETrigCounter_14_LC_6_14_4.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_14_LC_6_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_14_LC_6_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50378),
            .lcout(sEETrigCounterZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52333),
            .ce(N__21932),
            .sr(N__51695));
    defparam sEETrigCounter_15_LC_6_14_5.C_ON=1'b0;
    defparam sEETrigCounter_15_LC_6_14_5.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_15_LC_6_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_15_LC_6_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50049),
            .lcout(sEETrigCounterZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52333),
            .ce(N__21932),
            .sr(N__51695));
    defparam sEETrigCounter_8_LC_6_14_6.C_ON=1'b0;
    defparam sEETrigCounter_8_LC_6_14_6.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_8_LC_6_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_8_LC_6_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46281),
            .lcout(sEETrigCounterZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52333),
            .ce(N__21932),
            .sr(N__51695));
    defparam sEETrigCounter_9_LC_6_14_7.C_ON=1'b0;
    defparam sEETrigCounter_9_LC_6_14_7.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_9_LC_6_14_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 sEETrigCounter_9_LC_6_14_7 (
            .in0(_gnd_net_),
            .in1(N__51068),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEETrigCounterZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52333),
            .ce(N__21932),
            .sr(N__51695));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4Q_11_LC_7_3_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4Q_11_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4Q_11_LC_7_3_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4Q_11_LC_7_3_7  (
            .in0(N__25790),
            .in1(N__22316),
            .in2(_gnd_net_),
            .in3(N__24700),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_1_LC_7_4_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_1_LC_7_4_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_1_LC_7_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_1_LC_7_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23984),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48459),
            .ce(),
            .sr(N__51804));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_5_LC_7_4_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_5_LC_7_4_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_5_LC_7_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_5_LC_7_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21752),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48459),
            .ce(),
            .sr(N__51804));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_13_LC_7_4_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_13_LC_7_4_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_13_LC_7_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_13_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24041),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48459),
            .ce(),
            .sr(N__51804));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_14_LC_7_4_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_14_LC_7_4_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_14_LC_7_4_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_14_LC_7_4_6  (
            .in0(_gnd_net_),
            .in1(N__24032),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48459),
            .ce(),
            .sr(N__51804));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_0_LC_7_4_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_0_LC_7_4_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_0_LC_7_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_0_LC_7_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23993),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48459),
            .ce(),
            .sr(N__51804));
    defparam \spi_master_inst.spi_data_path_u1.data_in_6_LC_7_5_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_6_LC_7_5_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_6_LC_7_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_6_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27170),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48461),
            .ce(N__43902),
            .sr(N__51793));
    defparam \spi_master_inst.spi_data_path_u1.data_in_5_LC_7_5_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_5_LC_7_5_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_5_LC_7_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_5_LC_7_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37127),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48461),
            .ce(N__43902),
            .sr(N__51793));
    defparam sDAC_mem_35_0_LC_7_6_0.C_ON=1'b0;
    defparam sDAC_mem_35_0_LC_7_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_0_LC_7_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_0_LC_7_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46130),
            .lcout(sDAC_mem_35Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52342),
            .ce(N__22544),
            .sr(N__51779));
    defparam sDAC_mem_35_1_LC_7_6_1.C_ON=1'b0;
    defparam sDAC_mem_35_1_LC_7_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_1_LC_7_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_1_LC_7_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50717),
            .lcout(sDAC_mem_35Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52342),
            .ce(N__22544),
            .sr(N__51779));
    defparam sDAC_mem_35_2_LC_7_6_2.C_ON=1'b0;
    defparam sDAC_mem_35_2_LC_7_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_2_LC_7_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_2_LC_7_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47120),
            .lcout(sDAC_mem_35Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52342),
            .ce(N__22544),
            .sr(N__51779));
    defparam sDAC_mem_35_3_LC_7_6_3.C_ON=1'b0;
    defparam sDAC_mem_35_3_LC_7_6_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_3_LC_7_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_3_LC_7_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46520),
            .lcout(sDAC_mem_35Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52342),
            .ce(N__22544),
            .sr(N__51779));
    defparam sDAC_mem_35_4_LC_7_6_4.C_ON=1'b0;
    defparam sDAC_mem_35_4_LC_7_6_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_4_LC_7_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_4_LC_7_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45225),
            .lcout(sDAC_mem_35Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52342),
            .ce(N__22544),
            .sr(N__51779));
    defparam sDAC_mem_35_5_LC_7_6_5.C_ON=1'b0;
    defparam sDAC_mem_35_5_LC_7_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_5_LC_7_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_5_LC_7_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44732),
            .lcout(sDAC_mem_35Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52342),
            .ce(N__22544),
            .sr(N__51779));
    defparam sDAC_mem_35_6_LC_7_6_6.C_ON=1'b0;
    defparam sDAC_mem_35_6_LC_7_6_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_6_LC_7_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_6_LC_7_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50169),
            .lcout(sDAC_mem_35Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52342),
            .ce(N__22544),
            .sr(N__51779));
    defparam sDAC_mem_35_7_LC_7_6_7.C_ON=1'b0;
    defparam sDAC_mem_35_7_LC_7_6_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_7_LC_7_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_7_LC_7_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49671),
            .lcout(sDAC_mem_35Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52342),
            .ce(N__22544),
            .sr(N__51779));
    defparam sDAC_mem_22_0_LC_7_7_0.C_ON=1'b0;
    defparam sDAC_mem_22_0_LC_7_7_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_0_LC_7_7_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_22_0_LC_7_7_0 (
            .in0(N__46042),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_22Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52334),
            .ce(N__33883),
            .sr(N__51764));
    defparam sDAC_mem_22_1_LC_7_7_1.C_ON=1'b0;
    defparam sDAC_mem_22_1_LC_7_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_1_LC_7_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_1_LC_7_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50903),
            .lcout(sDAC_mem_22Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52334),
            .ce(N__33883),
            .sr(N__51764));
    defparam sDAC_mem_22_2_LC_7_7_2.C_ON=1'b0;
    defparam sDAC_mem_22_2_LC_7_7_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_2_LC_7_7_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_22_2_LC_7_7_2 (
            .in0(N__47202),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_22Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52334),
            .ce(N__33883),
            .sr(N__51764));
    defparam sDAC_mem_22_3_LC_7_7_3.C_ON=1'b0;
    defparam sDAC_mem_22_3_LC_7_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_3_LC_7_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_3_LC_7_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46604),
            .lcout(sDAC_mem_22Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52334),
            .ce(N__33883),
            .sr(N__51764));
    defparam sDAC_mem_22_7_LC_7_7_4.C_ON=1'b0;
    defparam sDAC_mem_22_7_LC_7_7_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_7_LC_7_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_7_LC_7_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49726),
            .lcout(sDAC_mem_22Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52334),
            .ce(N__33883),
            .sr(N__51764));
    defparam sAddress_RNIQ63A_6_LC_7_8_0.C_ON=1'b0;
    defparam sAddress_RNIQ63A_6_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNIQ63A_6_LC_7_8_0.LUT_INIT=16'b1111111101111111;
    LogicCell40 sAddress_RNIQ63A_6_LC_7_8_0 (
            .in0(N__21880),
            .in1(N__40861),
            .in2(N__21917),
            .in3(N__22609),
            .lcout(N_316),
            .ltout(N_316_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIUTJC_3_LC_7_8_1.C_ON=1'b0;
    defparam sAddress_RNIUTJC_3_LC_7_8_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNIUTJC_3_LC_7_8_1.LUT_INIT=16'b1111010111110101;
    LogicCell40 sAddress_RNIUTJC_3_LC_7_8_1 (
            .in0(N__40269),
            .in1(_gnd_net_),
            .in2(N__21830),
            .in3(_gnd_net_),
            .lcout(N_317),
            .ltout(N_317_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI8U0V1_1_LC_7_8_2.C_ON=1'b0;
    defparam sAddress_RNI8U0V1_1_LC_7_8_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI8U0V1_1_LC_7_8_2.LUT_INIT=16'b0000000100000000;
    LogicCell40 sAddress_RNI8U0V1_1_LC_7_8_2 (
            .in0(N__40632),
            .in1(N__40533),
            .in2(N__21827),
            .in3(N__33754),
            .lcout(sAddress_RNI8U0V1Z0Z_1),
            .ltout(sAddress_RNI8U0V1Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIETI62_1_LC_7_8_3.C_ON=1'b0;
    defparam sAddress_RNIETI62_1_LC_7_8_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNIETI62_1_LC_7_8_3.LUT_INIT=16'b0101000001010000;
    LogicCell40 sAddress_RNIETI62_1_LC_7_8_3 (
            .in0(N__23836),
            .in1(_gnd_net_),
            .in2(N__21824),
            .in3(_gnd_net_),
            .lcout(sAddress_RNIETI62Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_0_LC_7_8_4.C_ON=1'b0;
    defparam sAddress_RNI9IH12_0_LC_7_8_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_0_LC_7_8_4.LUT_INIT=16'b0101010100000000;
    LogicCell40 sAddress_RNI9IH12_0_LC_7_8_4 (
            .in0(N__40180),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21821),
            .lcout(sAddress_RNI9IH12Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPointerReset_RNO_0_LC_7_8_5.C_ON=1'b0;
    defparam sEEPointerReset_RNO_0_LC_7_8_5.SEQ_MODE=4'b0000;
    defparam sEEPointerReset_RNO_0_LC_7_8_5.LUT_INIT=16'b0000000010000000;
    LogicCell40 sEEPointerReset_RNO_0_LC_7_8_5 (
            .in0(N__33755),
            .in1(N__23345),
            .in2(N__49352),
            .in3(N__27092),
            .lcout(),
            .ltout(N_454_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPointerReset_LC_7_8_6.C_ON=1'b0;
    defparam sEEPointerReset_LC_7_8_6.SEQ_MODE=4'b1000;
    defparam sEEPointerReset_LC_7_8_6.LUT_INIT=16'b0000001011111110;
    LogicCell40 sEEPointerReset_LC_7_8_6 (
            .in0(N__39225),
            .in1(N__26006),
            .in2(N__21815),
            .in3(N__25952),
            .lcout(sEEPointerResetZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52324),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIBH15_4_LC_7_9_0.C_ON=1'b0;
    defparam sAddress_RNIBH15_4_LC_7_9_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNIBH15_4_LC_7_9_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 sAddress_RNIBH15_4_LC_7_9_0 (
            .in0(_gnd_net_),
            .in1(N__40871),
            .in2(_gnd_net_),
            .in3(N__22610),
            .lcout(),
            .ltout(N_346_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIUTJC_6_LC_7_9_1.C_ON=1'b0;
    defparam sAddress_RNIUTJC_6_LC_7_9_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNIUTJC_6_LC_7_9_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 sAddress_RNIUTJC_6_LC_7_9_1 (
            .in0(N__40410),
            .in1(N__21920),
            .in2(N__21938),
            .in3(N__21890),
            .lcout(),
            .ltout(un1_spointer11_8_0_0_a2_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI7G5E2_6_LC_7_9_2.C_ON=1'b0;
    defparam sAddress_RNI7G5E2_6_LC_7_9_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI7G5E2_6_LC_7_9_2.LUT_INIT=16'b0100000000000000;
    LogicCell40 sAddress_RNI7G5E2_6_LC_7_9_2 (
            .in0(N__23554),
            .in1(N__27093),
            .in2(N__21935),
            .in3(N__33747),
            .lcout(sAddress_RNI7G5E2Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_4_LC_7_9_3.C_ON=1'b0;
    defparam sAddress_4_LC_7_9_3.SEQ_MODE=4'b1010;
    defparam sAddress_4_LC_7_9_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 sAddress_4_LC_7_9_3 (
            .in0(_gnd_net_),
            .in1(N__45387),
            .in2(_gnd_net_),
            .in3(N__26166),
            .lcout(sAddressZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52312),
            .ce(N__23417),
            .sr(N__51738));
    defparam sAddress_5_LC_7_9_4.C_ON=1'b0;
    defparam sAddress_5_LC_7_9_4.SEQ_MODE=4'b1010;
    defparam sAddress_5_LC_7_9_4.LUT_INIT=16'b0101010100000000;
    LogicCell40 sAddress_5_LC_7_9_4 (
            .in0(N__26167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45037),
            .lcout(sAddressZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52312),
            .ce(N__23417),
            .sr(N__51738));
    defparam sAddress_RNIQ63A_0_6_LC_7_9_5.C_ON=1'b0;
    defparam sAddress_RNIQ63A_0_6_LC_7_9_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNIQ63A_0_6_LC_7_9_5.LUT_INIT=16'b0000100000000000;
    LogicCell40 sAddress_RNIQ63A_0_6_LC_7_9_5 (
            .in0(N__22611),
            .in1(N__21919),
            .in2(N__40900),
            .in3(N__21889),
            .lcout(sEEPonPoff_1_sqmuxa_0_a3_0_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIFL15_6_LC_7_9_7.C_ON=1'b0;
    defparam sAddress_RNIFL15_6_LC_7_9_7.SEQ_MODE=4'b0000;
    defparam sAddress_RNIFL15_6_LC_7_9_7.LUT_INIT=16'b0000000000110011;
    LogicCell40 sAddress_RNIFL15_6_LC_7_9_7 (
            .in0(_gnd_net_),
            .in1(N__21918),
            .in2(_gnd_net_),
            .in3(N__21888),
            .lcout(sDAC_mem_17_1_sqmuxa_0_a2_0_a2_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_0_LC_7_10_0 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_0_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_0_LC_7_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_0_LC_7_10_0  (
            .in0(N__24254),
            .in1(N__21859),
            .in2(N__24221),
            .in3(N__24220),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0 ),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51725));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_1_LC_7_10_1 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_1_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_1_LC_7_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_1_LC_7_10_1  (
            .in0(N__24256),
            .in1(N__21845),
            .in2(_gnd_net_),
            .in3(N__21833),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1 ),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51725));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_2_LC_7_10_2 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_2_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_2_LC_7_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_2_LC_7_10_2  (
            .in0(N__24255),
            .in1(N__22039),
            .in2(_gnd_net_),
            .in3(N__22025),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2 ),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51725));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_3_LC_7_10_3 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_3_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_3_LC_7_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_3_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(N__24286),
            .in2(_gnd_net_),
            .in3(N__22022),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3 ),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51725));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_4_LC_7_10_4 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_4_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_4_LC_7_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_4_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__24304),
            .in2(_gnd_net_),
            .in3(N__22019),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4 ),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51725));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_5_LC_7_10_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_5_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_5_LC_7_10_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_5_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(N__22013),
            .in2(_gnd_net_),
            .in3(N__22016),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51725));
    defparam \spi_slave_inst.rx_ready_i_LC_7_11_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_ready_i_LC_7_11_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_ready_i_LC_7_11_0 .LUT_INIT=16'b1110111111101100;
    LogicCell40 \spi_slave_inst.rx_ready_i_LC_7_11_0  (
            .in0(N__51223),
            .in1(N__22634),
            .in2(N__49353),
            .in3(N__21993),
            .lcout(spi_mosi_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52292),
            .ce(),
            .sr(N__51714));
    defparam spi_mosi_ready_prev_LC_7_11_1.C_ON=1'b0;
    defparam spi_mosi_ready_prev_LC_7_11_1.SEQ_MODE=4'b1010;
    defparam spi_mosi_ready_prev_LC_7_11_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 spi_mosi_ready_prev_LC_7_11_1 (
            .in0(N__21994),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_mosi_ready_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52292),
            .ce(),
            .sr(N__51714));
    defparam spi_mosi_ready_prev2_LC_7_11_2.C_ON=1'b0;
    defparam spi_mosi_ready_prev2_LC_7_11_2.SEQ_MODE=4'b1010;
    defparam spi_mosi_ready_prev2_LC_7_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 spi_mosi_ready_prev2_LC_7_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21971),
            .lcout(spi_mosi_ready_prevZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52292),
            .ce(),
            .sr(N__51714));
    defparam spi_mosi_ready_prev3_LC_7_11_3.C_ON=1'b0;
    defparam spi_mosi_ready_prev3_LC_7_11_3.SEQ_MODE=4'b1010;
    defparam spi_mosi_ready_prev3_LC_7_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 spi_mosi_ready_prev3_LC_7_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21959),
            .lcout(spi_mosi_ready_prevZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52292),
            .ce(),
            .sr(N__51714));
    defparam trig_prev_LC_7_11_4.C_ON=1'b0;
    defparam trig_prev_LC_7_11_4.SEQ_MODE=4'b1010;
    defparam trig_prev_LC_7_11_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 trig_prev_LC_7_11_4 (
            .in0(N__22798),
            .in1(N__22828),
            .in2(_gnd_net_),
            .in3(N__22758),
            .lcout(trig_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52292),
            .ce(),
            .sr(N__51714));
    defparam sEETrigCounter_RNIR6CE_0_LC_7_11_5.C_ON=1'b0;
    defparam sEETrigCounter_RNIR6CE_0_LC_7_11_5.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIR6CE_0_LC_7_11_5.LUT_INIT=16'b0011001100110011;
    LogicCell40 sEETrigCounter_RNIR6CE_0_LC_7_11_5 (
            .in0(_gnd_net_),
            .in1(N__22144),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un10_trig_prev_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_done_reg3_i_LC_7_11_7 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_reg3_i_LC_7_11_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_done_reg3_i_LC_7_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_done_reg3_i_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22670),
            .lcout(\spi_slave_inst.rx_done_reg3_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52292),
            .ce(),
            .sr(N__51714));
    defparam un10_trig_prev_cry_0_c_inv_LC_7_12_0.C_ON=1'b1;
    defparam un10_trig_prev_cry_0_c_inv_LC_7_12_0.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_0_c_inv_LC_7_12_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_0_c_inv_LC_7_12_0 (
            .in0(_gnd_net_),
            .in1(N__22121),
            .in2(N__22130),
            .in3(N__26562),
            .lcout(sTrigCounter_i_0),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(un10_trig_prev_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_1_c_inv_LC_7_12_1.C_ON=1'b1;
    defparam un10_trig_prev_cry_1_c_inv_LC_7_12_1.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_1_c_inv_LC_7_12_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_1_c_inv_LC_7_12_1 (
            .in0(_gnd_net_),
            .in1(N__22106),
            .in2(N__22115),
            .in3(N__26949),
            .lcout(sTrigCounter_i_1),
            .ltout(),
            .carryin(un10_trig_prev_cry_0),
            .carryout(un10_trig_prev_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_2_c_inv_LC_7_12_2.C_ON=1'b1;
    defparam un10_trig_prev_cry_2_c_inv_LC_7_12_2.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_2_c_inv_LC_7_12_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_2_c_inv_LC_7_12_2 (
            .in0(_gnd_net_),
            .in1(N__22091),
            .in2(N__22100),
            .in3(N__22858),
            .lcout(sTrigCounter_i_2),
            .ltout(),
            .carryin(un10_trig_prev_cry_1),
            .carryout(un10_trig_prev_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_3_c_inv_LC_7_12_3.C_ON=1'b1;
    defparam un10_trig_prev_cry_3_c_inv_LC_7_12_3.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_3_c_inv_LC_7_12_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_3_c_inv_LC_7_12_3 (
            .in0(_gnd_net_),
            .in1(N__22076),
            .in2(N__22085),
            .in3(N__22843),
            .lcout(sTrigCounter_i_3),
            .ltout(),
            .carryin(un10_trig_prev_cry_2),
            .carryout(un10_trig_prev_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_4_c_inv_LC_7_12_4.C_ON=1'b1;
    defparam un10_trig_prev_cry_4_c_inv_LC_7_12_4.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_4_c_inv_LC_7_12_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_4_c_inv_LC_7_12_4 (
            .in0(_gnd_net_),
            .in1(N__22061),
            .in2(N__22070),
            .in3(N__23071),
            .lcout(sTrigCounter_i_4),
            .ltout(),
            .carryin(un10_trig_prev_cry_3),
            .carryout(un10_trig_prev_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_5_c_inv_LC_7_12_5.C_ON=1'b1;
    defparam un10_trig_prev_cry_5_c_inv_LC_7_12_5.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_5_c_inv_LC_7_12_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 un10_trig_prev_cry_5_c_inv_LC_7_12_5 (
            .in0(N__23056),
            .in1(N__22046),
            .in2(N__22055),
            .in3(_gnd_net_),
            .lcout(sTrigCounter_i_5),
            .ltout(),
            .carryin(un10_trig_prev_cry_4),
            .carryout(un10_trig_prev_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_6_c_inv_LC_7_12_6.C_ON=1'b1;
    defparam un10_trig_prev_cry_6_c_inv_LC_7_12_6.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_6_c_inv_LC_7_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_6_c_inv_LC_7_12_6 (
            .in0(_gnd_net_),
            .in1(N__22256),
            .in2(N__22265),
            .in3(N__23041),
            .lcout(sTrigCounter_i_6),
            .ltout(),
            .carryin(un10_trig_prev_cry_5),
            .carryout(un10_trig_prev_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_7_c_inv_LC_7_12_7.C_ON=1'b1;
    defparam un10_trig_prev_cry_7_c_inv_LC_7_12_7.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_7_c_inv_LC_7_12_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_7_c_inv_LC_7_12_7 (
            .in0(_gnd_net_),
            .in1(N__22241),
            .in2(N__22250),
            .in3(N__23026),
            .lcout(sTrigCounter_i_7),
            .ltout(),
            .carryin(un10_trig_prev_cry_6),
            .carryout(un10_trig_prev_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_8_c_inv_LC_7_13_0.C_ON=1'b1;
    defparam un10_trig_prev_cry_8_c_inv_LC_7_13_0.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_8_c_inv_LC_7_13_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_8_c_inv_LC_7_13_0 (
            .in0(_gnd_net_),
            .in1(N__22226),
            .in2(N__22235),
            .in3(N__23011),
            .lcout(sTrigCounter_i_8),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(un10_trig_prev_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_9_c_inv_LC_7_13_1.C_ON=1'b1;
    defparam un10_trig_prev_cry_9_c_inv_LC_7_13_1.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_9_c_inv_LC_7_13_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_9_c_inv_LC_7_13_1 (
            .in0(_gnd_net_),
            .in1(N__22211),
            .in2(N__22220),
            .in3(N__22996),
            .lcout(sTrigCounter_i_9),
            .ltout(),
            .carryin(un10_trig_prev_cry_8),
            .carryout(un10_trig_prev_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_10_c_inv_LC_7_13_2.C_ON=1'b1;
    defparam un10_trig_prev_cry_10_c_inv_LC_7_13_2.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_10_c_inv_LC_7_13_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 un10_trig_prev_cry_10_c_inv_LC_7_13_2 (
            .in0(N__22981),
            .in1(N__22196),
            .in2(N__22205),
            .in3(_gnd_net_),
            .lcout(sTrigCounter_i_10),
            .ltout(),
            .carryin(un10_trig_prev_cry_9),
            .carryout(un10_trig_prev_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_11_c_inv_LC_7_13_3.C_ON=1'b1;
    defparam un10_trig_prev_cry_11_c_inv_LC_7_13_3.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_11_c_inv_LC_7_13_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_11_c_inv_LC_7_13_3 (
            .in0(_gnd_net_),
            .in1(N__22181),
            .in2(N__22190),
            .in3(N__22966),
            .lcout(sTrigCounter_i_11),
            .ltout(),
            .carryin(un10_trig_prev_cry_10),
            .carryout(un10_trig_prev_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_12_c_inv_LC_7_13_4.C_ON=1'b1;
    defparam un10_trig_prev_cry_12_c_inv_LC_7_13_4.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_12_c_inv_LC_7_13_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 un10_trig_prev_cry_12_c_inv_LC_7_13_4 (
            .in0(N__22951),
            .in1(N__22166),
            .in2(N__22175),
            .in3(_gnd_net_),
            .lcout(sTrigCounter_i_12),
            .ltout(),
            .carryin(un10_trig_prev_cry_11),
            .carryout(un10_trig_prev_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_13_c_inv_LC_7_13_5.C_ON=1'b1;
    defparam un10_trig_prev_cry_13_c_inv_LC_7_13_5.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_13_c_inv_LC_7_13_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_13_c_inv_LC_7_13_5 (
            .in0(_gnd_net_),
            .in1(N__22151),
            .in2(N__22160),
            .in3(N__23128),
            .lcout(sTrigCounter_i_13),
            .ltout(),
            .carryin(un10_trig_prev_cry_12),
            .carryout(un10_trig_prev_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_14_c_inv_LC_7_13_6.C_ON=1'b1;
    defparam un10_trig_prev_cry_14_c_inv_LC_7_13_6.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_14_c_inv_LC_7_13_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_14_c_inv_LC_7_13_6 (
            .in0(_gnd_net_),
            .in1(N__22301),
            .in2(N__22310),
            .in3(N__23113),
            .lcout(sTrigCounter_i_14),
            .ltout(),
            .carryin(un10_trig_prev_cry_13),
            .carryout(un10_trig_prev_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_15_c_inv_LC_7_13_7.C_ON=1'b1;
    defparam un10_trig_prev_cry_15_c_inv_LC_7_13_7.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_15_c_inv_LC_7_13_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_15_c_inv_LC_7_13_7 (
            .in0(_gnd_net_),
            .in1(N__22286),
            .in2(N__22295),
            .in3(N__23095),
            .lcout(sTrigCounter_i_15),
            .ltout(),
            .carryin(un10_trig_prev_cry_14),
            .carryout(un10_trig_prev_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_15_THRU_LUT4_0_LC_7_14_0.C_ON=1'b0;
    defparam un10_trig_prev_cry_15_THRU_LUT4_0_LC_7_14_0.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_15_THRU_LUT4_0_LC_7_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un10_trig_prev_cry_15_THRU_LUT4_0_LC_7_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22280),
            .lcout(un10_trig_prev_cry_15_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_rpi_ibuf_RNI4GQD1_LC_7_14_4.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNI4GQD1_LC_7_14_4.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNI4GQD1_LC_7_14_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 reset_rpi_ibuf_RNI4GQD1_LC_7_14_4 (
            .in0(_gnd_net_),
            .in1(N__49354),
            .in2(_gnd_net_),
            .in3(N__22277),
            .lcout(N_82_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_prev_RNIIHS91_LC_7_14_5.C_ON=1'b0;
    defparam trig_prev_RNIIHS91_LC_7_14_5.SEQ_MODE=4'b0000;
    defparam trig_prev_RNIIHS91_LC_7_14_5.LUT_INIT=16'b1011101110110000;
    LogicCell40 trig_prev_RNIIHS91_LC_7_14_5 (
            .in0(N__23656),
            .in1(N__23720),
            .in2(N__22381),
            .in3(N__22726),
            .lcout(N_173),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_ft_ibuf_RNI4OFN_LC_7_14_6.C_ON=1'b0;
    defparam trig_ft_ibuf_RNI4OFN_LC_7_14_6.SEQ_MODE=4'b0000;
    defparam trig_ft_ibuf_RNI4OFN_LC_7_14_6.LUT_INIT=16'b0000000000010001;
    LogicCell40 trig_ft_ibuf_RNI4OFN_LC_7_14_6 (
            .in0(N__22785),
            .in1(N__22829),
            .in2(_gnd_net_),
            .in3(N__22766),
            .lcout(un3_trig_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_done_neg_sclk_i_LC_7_15_2 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_neg_sclk_i_LC_7_15_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_done_neg_sclk_i_LC_7_15_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \spi_slave_inst.rx_done_neg_sclk_i_LC_7_15_2  (
            .in0(N__51227),
            .in1(N__22576),
            .in2(_gnd_net_),
            .in3(N__24257),
            .lcout(\spi_slave_inst.rx_done_neg_sclk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVspi_slave_inst.rx_done_neg_sclk_iC_net ),
            .ce(),
            .sr(N__51681));
    defparam sEEADC_freq_RNICSIA1_4_LC_7_16_0.C_ON=1'b0;
    defparam sEEADC_freq_RNICSIA1_4_LC_7_16_0.SEQ_MODE=4'b0000;
    defparam sEEADC_freq_RNICSIA1_4_LC_7_16_0.LUT_INIT=16'b1000001001000001;
    LogicCell40 sEEADC_freq_RNICSIA1_4_LC_7_16_0 (
            .in0(N__22271),
            .in1(N__43052),
            .in2(N__22364),
            .in3(N__43079),
            .lcout(un11_sacqtime_NE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEADC_freq_4_LC_7_16_1.C_ON=1'b0;
    defparam sEEADC_freq_4_LC_7_16_1.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_4_LC_7_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEADC_freq_4_LC_7_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45576),
            .lcout(sEEADC_freqZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52343),
            .ce(N__49561),
            .sr(_gnd_net_));
    defparam sTrigInternal_RNO_2_LC_7_16_3.C_ON=1'b0;
    defparam sTrigInternal_RNO_2_LC_7_16_3.SEQ_MODE=4'b0000;
    defparam sTrigInternal_RNO_2_LC_7_16_3.LUT_INIT=16'b0100010001001111;
    LogicCell40 sTrigInternal_RNO_2_LC_7_16_3 (
            .in0(N__23655),
            .in1(N__23719),
            .in2(N__22385),
            .in3(N__22727),
            .lcout(un1_scounter_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEADC_freq_5_LC_7_16_6.C_ON=1'b0;
    defparam sEEADC_freq_5_LC_7_16_6.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_5_LC_7_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEADC_freq_5_LC_7_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45009),
            .lcout(sEEADC_freqZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52343),
            .ce(N__49561),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_1_LC_8_2_1 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_1_LC_8_2_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_1_LC_8_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_1_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22480),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48259),
            .ce(N__48231),
            .sr(N__51812));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_0_LC_8_2_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_0_LC_8_2_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_0_LC_8_2_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_0_LC_8_2_5  (
            .in0(N__22355),
            .in1(N__48011),
            .in2(_gnd_net_),
            .in3(N__22337),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48259),
            .ce(N__48231),
            .sr(N__51812));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_11_LC_8_3_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_11_LC_8_3_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_11_LC_8_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_11_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24053),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48455),
            .ce(),
            .sr(N__51805));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_6_LC_8_4_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_6_LC_8_4_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_6_LC_8_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_6_LC_8_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22414),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48260),
            .ce(N__48236),
            .sr(N__51794));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_2_LC_8_4_2 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_2_LC_8_4_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_2_LC_8_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_2_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22465),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48260),
            .ce(N__48236),
            .sr(N__51794));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_3_LC_8_4_3 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_3_LC_8_4_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_3_LC_8_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_3_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22450),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48260),
            .ce(N__48236),
            .sr(N__51794));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_4_LC_8_4_4 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_4_LC_8_4_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_4_LC_8_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_4_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22438),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48260),
            .ce(N__48236),
            .sr(N__51794));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_5_LC_8_4_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_5_LC_8_4_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_5_LC_8_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_5_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22426),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48260),
            .ce(N__48236),
            .sr(N__51794));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_7_LC_8_4_7 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_7_LC_8_4_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_7_LC_8_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_7_LC_8_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22402),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48260),
            .ce(N__48236),
            .sr(N__51794));
    defparam \spi_slave_inst.rxdata_reg_i_0_LC_8_5_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_0_LC_8_5_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_0_LC_8_5_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_0_LC_8_5_0  (
            .in0(N__22484),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_data_mosi_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52344),
            .ce(N__22565),
            .sr(N__51780));
    defparam \spi_slave_inst.rxdata_reg_i_1_LC_8_5_1 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_1_LC_8_5_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_1_LC_8_5_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_1_LC_8_5_1  (
            .in0(N__22469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_data_mosi_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52344),
            .ce(N__22565),
            .sr(N__51780));
    defparam \spi_slave_inst.rxdata_reg_i_2_LC_8_5_2 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_2_LC_8_5_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_2_LC_8_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_2_LC_8_5_2  (
            .in0(N__22451),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_data_mosi_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52344),
            .ce(N__22565),
            .sr(N__51780));
    defparam \spi_slave_inst.rxdata_reg_i_3_LC_8_5_3 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_3_LC_8_5_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_3_LC_8_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_3_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22439),
            .lcout(spi_data_mosi_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52344),
            .ce(N__22565),
            .sr(N__51780));
    defparam \spi_slave_inst.rxdata_reg_i_4_LC_8_5_4 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_4_LC_8_5_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_4_LC_8_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_4_LC_8_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22427),
            .lcout(spi_data_mosi_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52344),
            .ce(N__22565),
            .sr(N__51780));
    defparam \spi_slave_inst.rxdata_reg_i_5_LC_8_5_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_5_LC_8_5_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_5_LC_8_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_5_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22415),
            .lcout(spi_data_mosi_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52344),
            .ce(N__22565),
            .sr(N__51780));
    defparam \spi_slave_inst.rxdata_reg_i_6_LC_8_5_6 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_6_LC_8_5_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_6_LC_8_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_6_LC_8_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22403),
            .lcout(spi_data_mosi_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52344),
            .ce(N__22565),
            .sr(N__51780));
    defparam \spi_slave_inst.rxdata_reg_i_7_LC_8_5_7 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_7_LC_8_5_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_7_LC_8_5_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_7_LC_8_5_7  (
            .in0(N__22391),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_data_mosi_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52344),
            .ce(N__22565),
            .sr(N__51780));
    defparam sDAC_mem_11_0_LC_8_6_0.C_ON=1'b0;
    defparam sDAC_mem_11_0_LC_8_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_0_LC_8_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_0_LC_8_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45978),
            .lcout(sDAC_mem_11Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52335),
            .ce(N__22493),
            .sr(N__51765));
    defparam sDAC_mem_11_1_LC_8_6_1.C_ON=1'b0;
    defparam sDAC_mem_11_1_LC_8_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_1_LC_8_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_1_LC_8_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50716),
            .lcout(sDAC_mem_11Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52335),
            .ce(N__22493),
            .sr(N__51765));
    defparam sDAC_mem_11_2_LC_8_6_2.C_ON=1'b0;
    defparam sDAC_mem_11_2_LC_8_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_2_LC_8_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_2_LC_8_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47119),
            .lcout(sDAC_mem_11Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52335),
            .ce(N__22493),
            .sr(N__51765));
    defparam sDAC_mem_11_3_LC_8_6_3.C_ON=1'b0;
    defparam sDAC_mem_11_3_LC_8_6_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_3_LC_8_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_3_LC_8_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46519),
            .lcout(sDAC_mem_11Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52335),
            .ce(N__22493),
            .sr(N__51765));
    defparam sDAC_mem_11_4_LC_8_6_4.C_ON=1'b0;
    defparam sDAC_mem_11_4_LC_8_6_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_4_LC_8_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_4_LC_8_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45388),
            .lcout(sDAC_mem_11Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52335),
            .ce(N__22493),
            .sr(N__51765));
    defparam sDAC_mem_11_5_LC_8_6_5.C_ON=1'b0;
    defparam sDAC_mem_11_5_LC_8_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_5_LC_8_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_5_LC_8_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44731),
            .lcout(sDAC_mem_11Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52335),
            .ce(N__22493),
            .sr(N__51765));
    defparam sDAC_mem_11_6_LC_8_6_6.C_ON=1'b0;
    defparam sDAC_mem_11_6_LC_8_6_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_6_LC_8_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_6_LC_8_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50168),
            .lcout(sDAC_mem_11Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52335),
            .ce(N__22493),
            .sr(N__51765));
    defparam sDAC_mem_11_7_LC_8_6_7.C_ON=1'b0;
    defparam sDAC_mem_11_7_LC_8_6_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_7_LC_8_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_7_LC_8_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49655),
            .lcout(sDAC_mem_11Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52335),
            .ce(N__22493),
            .sr(N__51765));
    defparam sAddress_RNI9IH12_15_5_LC_8_7_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_15_5_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_15_5_LC_8_7_0.LUT_INIT=16'b0000010000000000;
    LogicCell40 sAddress_RNI9IH12_15_5_LC_8_7_0 (
            .in0(N__34857),
            .in1(N__40306),
            .in2(N__40998),
            .in3(N__40753),
            .lcout(sDAC_mem_11_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_19_5_LC_8_7_1.C_ON=1'b0;
    defparam sAddress_RNI9IH12_19_5_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_19_5_LC_8_7_1.LUT_INIT=16'b0000000000000010;
    LogicCell40 sAddress_RNI9IH12_19_5_LC_8_7_1 (
            .in0(N__40751),
            .in1(N__40294),
            .in2(N__40976),
            .in3(N__34858),
            .lcout(sDAC_mem_3_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_3_LC_8_7_2.C_ON=1'b0;
    defparam sAddress_3_LC_8_7_2.SEQ_MODE=4'b1010;
    defparam sAddress_3_LC_8_7_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 sAddress_3_LC_8_7_2 (
            .in0(_gnd_net_),
            .in1(N__46603),
            .in2(_gnd_net_),
            .in3(N__26163),
            .lcout(sAddressZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52325),
            .ce(N__23413),
            .sr(N__51752));
    defparam sEETrigInternal_RNO_2_LC_8_7_3.C_ON=1'b0;
    defparam sEETrigInternal_RNO_2_LC_8_7_3.SEQ_MODE=4'b0000;
    defparam sEETrigInternal_RNO_2_LC_8_7_3.LUT_INIT=16'b1111111111011101;
    LogicCell40 sEETrigInternal_RNO_2_LC_8_7_3 (
            .in0(N__40307),
            .in1(N__34853),
            .in2(_gnd_net_),
            .in3(N__23445),
            .lcout(),
            .ltout(N_344_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigInternal_RNO_1_LC_8_7_4.C_ON=1'b0;
    defparam sEETrigInternal_RNO_1_LC_8_7_4.SEQ_MODE=4'b0000;
    defparam sEETrigInternal_RNO_1_LC_8_7_4.LUT_INIT=16'b1000100010001101;
    LogicCell40 sEETrigInternal_RNO_1_LC_8_7_4 (
            .in0(N__26087),
            .in1(N__23705),
            .in2(N__22547),
            .in3(N__25945),
            .lcout(sEETrigInternal_3_iv_0_0_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_6_5_LC_8_7_5.C_ON=1'b0;
    defparam sAddress_RNI9IH12_6_5_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_6_5_LC_8_7_5.LUT_INIT=16'b0000000000100000;
    LogicCell40 sAddress_RNI9IH12_6_5_LC_8_7_5 (
            .in0(N__40752),
            .in1(N__40295),
            .in2(N__40977),
            .in3(N__34859),
            .lcout(sDAC_mem_35_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigInternal_RNO_0_LC_8_7_6.C_ON=1'b0;
    defparam sEETrigInternal_RNO_0_LC_8_7_6.SEQ_MODE=4'b0000;
    defparam sEETrigInternal_RNO_0_LC_8_7_6.LUT_INIT=16'b1100100000000000;
    LogicCell40 sEETrigInternal_RNO_0_LC_8_7_6 (
            .in0(N__27091),
            .in1(N__23704),
            .in2(N__34866),
            .in3(N__26162),
            .lcout(N_1631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEESingleCont_RNO_0_LC_8_7_7.C_ON=1'b0;
    defparam sEESingleCont_RNO_0_LC_8_7_7.SEQ_MODE=4'b0000;
    defparam sEESingleCont_RNO_0_LC_8_7_7.LUT_INIT=16'b0000000000100000;
    LogicCell40 sEESingleCont_RNO_0_LC_8_7_7 (
            .in0(N__26041),
            .in1(N__26088),
            .in2(N__26184),
            .in3(N__27090),
            .lcout(sEESingleCont_RNOZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEESingleCont_LC_8_8_0.C_ON=1'b0;
    defparam sEESingleCont_LC_8_8_0.SEQ_MODE=4'b1010;
    defparam sEESingleCont_LC_8_8_0.LUT_INIT=16'b1110010011001100;
    LogicCell40 sEESingleCont_LC_8_8_0 (
            .in0(N__23490),
            .in1(N__22522),
            .in2(N__46211),
            .in3(N__22532),
            .lcout(sEESingleContZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52313),
            .ce(),
            .sr(N__51739));
    defparam sEETrigInternal_LC_8_8_1.C_ON=1'b0;
    defparam sEETrigInternal_LC_8_8_1.SEQ_MODE=4'b1010;
    defparam sEETrigInternal_LC_8_8_1.LUT_INIT=16'b1111101111001000;
    LogicCell40 sEETrigInternal_LC_8_8_1 (
            .in0(N__22508),
            .in1(N__26043),
            .in2(N__22502),
            .in3(N__23706),
            .lcout(sEETrigInternalZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52313),
            .ce(),
            .sr(N__51739));
    defparam sEETrigInternal_prev_LC_8_8_2.C_ON=1'b0;
    defparam sEETrigInternal_prev_LC_8_8_2.SEQ_MODE=4'b1010;
    defparam sEETrigInternal_prev_LC_8_8_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEETrigInternal_prev_LC_8_8_2 (
            .in0(N__23707),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEETrigInternal_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52313),
            .ce(),
            .sr(N__51739));
    defparam sPointer_1_LC_8_8_3.C_ON=1'b0;
    defparam sPointer_1_LC_8_8_3.SEQ_MODE=4'b1010;
    defparam sPointer_1_LC_8_8_3.LUT_INIT=16'b0011100000111000;
    LogicCell40 sPointer_1_LC_8_8_3 (
            .in0(N__26089),
            .in1(N__26042),
            .in2(N__26193),
            .in3(_gnd_net_),
            .lcout(sPointerZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52313),
            .ce(),
            .sr(N__51739));
    defparam sPointer_0_LC_8_8_4.C_ON=1'b0;
    defparam sPointer_0_LC_8_8_4.SEQ_MODE=4'b1010;
    defparam sPointer_0_LC_8_8_4.LUT_INIT=16'b0101010100100000;
    LogicCell40 sPointer_0_LC_8_8_4 (
            .in0(N__26044),
            .in1(N__26174),
            .in2(N__25046),
            .in3(N__26090),
            .lcout(sPointerZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52313),
            .ce(),
            .sr(N__51739));
    defparam \spi_slave_inst.rx_done_reg1_i_LC_8_8_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_reg1_i_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_done_reg1_i_LC_8_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi_slave_inst.rx_done_reg1_i_LC_8_8_5  (
            .in0(N__51216),
            .in1(N__48284),
            .in2(_gnd_net_),
            .in3(N__22586),
            .lcout(\spi_slave_inst.rx_done_reg1_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52313),
            .ce(),
            .sr(N__51739));
    defparam \spi_slave_inst.rx_done_reg1_i_RNID541_LC_8_8_6 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_reg1_i_RNID541_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_done_reg1_i_RNID541_LC_8_8_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \spi_slave_inst.rx_done_reg1_i_RNID541_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__22555),
            .in2(_gnd_net_),
            .in3(N__22663),
            .lcout(\spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_done_reg2_i_LC_8_8_7 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_reg2_i_LC_8_8_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_done_reg2_i_LC_8_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.rx_done_reg2_i_LC_8_8_7  (
            .in0(N__22556),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_inst.rx_done_reg2_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52313),
            .ce(),
            .sr(N__51739));
    defparam sAddress_RNI9IH12_5_LC_8_9_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_5_LC_8_9_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_5_LC_8_9_0.LUT_INIT=16'b1010000000000000;
    LogicCell40 sAddress_RNI9IH12_5_LC_8_9_0 (
            .in0(N__40895),
            .in1(_gnd_net_),
            .in2(N__26977),
            .in3(N__40744),
            .lcout(sDAC_mem_37_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_18_5_LC_8_9_1.C_ON=1'b0;
    defparam sAddress_RNI9IH12_18_5_LC_8_9_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_18_5_LC_8_9_1.LUT_INIT=16'b0000000000000010;
    LogicCell40 sAddress_RNI9IH12_18_5_LC_8_9_1 (
            .in0(N__40742),
            .in1(N__40407),
            .in2(N__23565),
            .in3(N__40894),
            .lcout(sDAC_mem_7_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_0_3_LC_8_9_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_0_3_LC_8_9_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_0_3_LC_8_9_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 sAddress_RNI9IH12_0_3_LC_8_9_2 (
            .in0(N__23340),
            .in1(N__40406),
            .in2(_gnd_net_),
            .in3(N__39970),
            .lcout(sDAC_mem_32_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_7_5_LC_8_9_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_7_5_LC_8_9_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_7_5_LC_8_9_3.LUT_INIT=16'b0000001000000000;
    LogicCell40 sAddress_RNI9IH12_7_5_LC_8_9_3 (
            .in0(N__40743),
            .in1(N__40409),
            .in2(N__23566),
            .in3(N__40896),
            .lcout(sDAC_mem_39_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI6VH7_1_1_LC_8_9_4.C_ON=1'b0;
    defparam sAddress_RNI6VH7_1_1_LC_8_9_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI6VH7_1_1_LC_8_9_4.LUT_INIT=16'b1111011111110111;
    LogicCell40 sAddress_RNI6VH7_1_1_LC_8_9_4 (
            .in0(N__40620),
            .in1(N__40500),
            .in2(N__40195),
            .in3(_gnd_net_),
            .lcout(N_319),
            .ltout(N_319_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_9_3_LC_8_9_5.C_ON=1'b0;
    defparam sAddress_RNI9IH12_9_3_LC_8_9_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_9_3_LC_8_9_5.LUT_INIT=16'b0000000000001010;
    LogicCell40 sAddress_RNI9IH12_9_3_LC_8_9_5 (
            .in0(N__39971),
            .in1(_gnd_net_),
            .in2(N__22685),
            .in3(N__40408),
            .lcout(sDAC_mem_23_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_2_1_LC_8_9_6.C_ON=1'b0;
    defparam sAddress_RNI9IH12_2_1_LC_8_9_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_2_1_LC_8_9_6.LUT_INIT=16'b0001000100000000;
    LogicCell40 sAddress_RNI9IH12_2_1_LC_8_9_6 (
            .in0(N__23561),
            .in1(N__27094),
            .in2(_gnd_net_),
            .in3(N__33744),
            .lcout(sAddress_RNI9IH12_2Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_ready_i_RNO_0_LC_8_9_7 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_ready_i_RNO_0_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_ready_i_RNO_0_LC_8_9_7 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \spi_slave_inst.rx_ready_i_RNO_0_LC_8_9_7  (
            .in0(N__22662),
            .in1(_gnd_net_),
            .in2(N__22646),
            .in3(_gnd_net_),
            .lcout(\spi_slave_inst.rx_ready_i_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_10_5_LC_8_10_1.C_ON=1'b0;
    defparam sAddress_RNI9IH12_10_5_LC_8_10_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_10_5_LC_8_10_1.LUT_INIT=16'b0100000000000000;
    LogicCell40 sAddress_RNI9IH12_10_5_LC_8_10_1 (
            .in0(N__40864),
            .in1(N__40404),
            .in2(N__27061),
            .in3(N__40747),
            .lcout(sDAC_mem_13_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_3_LC_8_10_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_3_LC_8_10_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_3_LC_8_10_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 sAddress_RNI9IH12_3_LC_8_10_2 (
            .in0(N__40405),
            .in1(N__27057),
            .in2(_gnd_net_),
            .in3(N__39969),
            .lcout(sDAC_mem_29_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sPointer_RNI5LBD1_0_LC_8_10_3.C_ON=1'b0;
    defparam sPointer_RNI5LBD1_0_LC_8_10_3.SEQ_MODE=4'b0000;
    defparam sPointer_RNI5LBD1_0_LC_8_10_3.LUT_INIT=16'b0010001000000000;
    LogicCell40 sPointer_RNI5LBD1_0_LC_8_10_3 (
            .in0(N__26178),
            .in1(N__26091),
            .in2(_gnd_net_),
            .in3(N__26027),
            .lcout(sPointer_RNI5LBD1Z0Z_0),
            .ltout(sPointer_RNI5LBD1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIVREN1_4_LC_8_10_4.C_ON=1'b0;
    defparam sAddress_RNIVREN1_4_LC_8_10_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNIVREN1_4_LC_8_10_4.LUT_INIT=16'b0100000000000000;
    LogicCell40 sAddress_RNIVREN1_4_LC_8_10_4 (
            .in0(N__22613),
            .in1(N__22622),
            .in2(N__22625),
            .in3(N__40862),
            .lcout(sAddress_RNIVREN1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIP2UK1_4_LC_8_10_5.C_ON=1'b0;
    defparam sAddress_RNIP2UK1_4_LC_8_10_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNIP2UK1_4_LC_8_10_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 sAddress_RNIP2UK1_4_LC_8_10_5 (
            .in0(N__22621),
            .in1(N__22612),
            .in2(_gnd_net_),
            .in3(N__33732),
            .lcout(sAddress_RNIP2UK1Z0Z_4),
            .ltout(sAddress_RNIP2UK1Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_11_5_LC_8_10_6.C_ON=1'b0;
    defparam sAddress_RNI9IH12_11_5_LC_8_10_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_11_5_LC_8_10_6.LUT_INIT=16'b0000000010000000;
    LogicCell40 sAddress_RNI9IH12_11_5_LC_8_10_6 (
            .in0(N__40403),
            .in1(N__23344),
            .in2(N__22589),
            .in3(N__40863),
            .lcout(sDAC_mem_16_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_1_1_LC_8_10_7.C_ON=1'b0;
    defparam sAddress_RNI9IH12_1_1_LC_8_10_7.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_1_1_LC_8_10_7.LUT_INIT=16'b0010001000000000;
    LogicCell40 sAddress_RNI9IH12_1_1_LC_8_10_7 (
            .in0(N__40073),
            .in1(N__23464),
            .in2(_gnd_net_),
            .in3(N__33733),
            .lcout(sEEPon_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_prev_RNIM2UO_LC_8_11_0.C_ON=1'b0;
    defparam trig_prev_RNIM2UO_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam trig_prev_RNIM2UO_LC_8_11_0.LUT_INIT=16'b1111111100000001;
    LogicCell40 trig_prev_RNIM2UO_LC_8_11_0 (
            .in0(N__22827),
            .in1(N__22799),
            .in2(N__22762),
            .in3(N__22716),
            .lcout(g3_0),
            .ltout(g3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigInternal_prev_RNIIHS91_LC_8_11_1.C_ON=1'b0;
    defparam sEETrigInternal_prev_RNIIHS91_LC_8_11_1.SEQ_MODE=4'b0000;
    defparam sEETrigInternal_prev_RNIIHS91_LC_8_11_1.LUT_INIT=16'b1010000011110000;
    LogicCell40 sEETrigInternal_prev_RNIIHS91_LC_8_11_1 (
            .in0(N__23645),
            .in1(_gnd_net_),
            .in2(N__22703),
            .in3(N__23711),
            .lcout(g1_i_a4_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI70I7_1_LC_8_11_3.C_ON=1'b0;
    defparam sAddress_RNI70I7_1_LC_8_11_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI70I7_1_LC_8_11_3.LUT_INIT=16'b0010001000000000;
    LogicCell40 sAddress_RNI70I7_1_LC_8_11_3 (
            .in0(N__40175),
            .in1(N__40402),
            .in2(_gnd_net_),
            .in3(N__40509),
            .lcout(sAddress_RNI70I7Z0Z_1),
            .ltout(sAddress_RNI70I7Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_5_2_LC_8_11_4.C_ON=1'b0;
    defparam sAddress_RNI9IH12_5_2_LC_8_11_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_5_2_LC_8_11_4.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNI9IH12_5_2_LC_8_11_4 (
            .in0(N__40950),
            .in1(N__40647),
            .in2(N__22700),
            .in3(N__40740),
            .lcout(sDAC_mem_4_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI25GS1_1_LC_8_11_5.C_ON=1'b0;
    defparam sAddress_RNI25GS1_1_LC_8_11_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNI25GS1_1_LC_8_11_5.LUT_INIT=16'b0001001000000000;
    LogicCell40 sAddress_RNI25GS1_1_LC_8_11_5 (
            .in0(N__40176),
            .in1(N__23461),
            .in2(N__40531),
            .in3(N__33739),
            .lcout(un1_spointer11_5_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_rpi_ibuf_RNI3E6DF_LC_8_12_0.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNI3E6DF_LC_8_12_0.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNI3E6DF_LC_8_12_0.LUT_INIT=16'b1100111111001101;
    LogicCell40 reset_rpi_ibuf_RNI3E6DF_LC_8_12_0 (
            .in0(N__22697),
            .in1(N__22691),
            .in2(N__23762),
            .in3(N__22925),
            .lcout(un1_reset_rpi_inv_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_15_c_RNIGF876_LC_8_12_1.C_ON=1'b0;
    defparam un10_trig_prev_cry_15_c_RNIGF876_LC_8_12_1.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_15_c_RNIGF876_LC_8_12_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 un10_trig_prev_cry_15_c_RNIGF876_LC_8_12_1 (
            .in0(N__23798),
            .in1(N__23507),
            .in2(N__23849),
            .in3(N__22938),
            .lcout(N_8_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigInternal_RNO_1_LC_8_12_2.C_ON=1'b0;
    defparam sTrigInternal_RNO_1_LC_8_12_2.SEQ_MODE=4'b0000;
    defparam sTrigInternal_RNO_1_LC_8_12_2.LUT_INIT=16'b1111100011110000;
    LogicCell40 sTrigInternal_RNO_1_LC_8_12_2 (
            .in0(N__22940),
            .in1(N__23608),
            .in2(N__31048),
            .in3(N__22893),
            .lcout(N_96),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_15_c_RNI3GF11_LC_8_12_3.C_ON=1'b0;
    defparam un10_trig_prev_cry_15_c_RNI3GF11_LC_8_12_3.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_15_c_RNI3GF11_LC_8_12_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 un10_trig_prev_cry_15_c_RNI3GF11_LC_8_12_3 (
            .in0(N__23607),
            .in1(N__25159),
            .in2(N__22895),
            .in3(N__22939),
            .lcout(N_178),
            .ltout(N_178_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigInternal_RNO_0_LC_8_12_4.C_ON=1'b0;
    defparam sTrigInternal_RNO_0_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam sTrigInternal_RNO_0_LC_8_12_4.LUT_INIT=16'b1111101111111010;
    LogicCell40 sTrigInternal_RNO_0_LC_8_12_4 (
            .in0(N__22919),
            .in1(N__29554),
            .in2(N__22907),
            .in3(N__22904),
            .lcout(),
            .ltout(N_77_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigInternal_LC_8_12_5.C_ON=1'b0;
    defparam sTrigInternal_LC_8_12_5.SEQ_MODE=4'b1010;
    defparam sTrigInternal_LC_8_12_5.LUT_INIT=16'b1111110001011100;
    LogicCell40 sTrigInternal_LC_8_12_5 (
            .in0(N__31033),
            .in1(N__25206),
            .in2(N__22898),
            .in3(N__29556),
            .lcout(sTrigInternalZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52293),
            .ce(),
            .sr(N__51696));
    defparam sPeriod_prev_LC_8_12_6.C_ON=1'b0;
    defparam sPeriod_prev_LC_8_12_6.SEQ_MODE=4'b1010;
    defparam sPeriod_prev_LC_8_12_6.LUT_INIT=16'b0101010101000100;
    LogicCell40 sPeriod_prev_LC_8_12_6 (
            .in0(N__25160),
            .in1(N__29555),
            .in2(_gnd_net_),
            .in3(N__31034),
            .lcout(sPeriod_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52293),
            .ce(),
            .sr(N__51696));
    defparam sPeriod_prev_RNI43A11_LC_8_12_7.C_ON=1'b0;
    defparam sPeriod_prev_RNI43A11_LC_8_12_7.SEQ_MODE=4'b0000;
    defparam sPeriod_prev_RNI43A11_LC_8_12_7.LUT_INIT=16'b0000000000010000;
    LogicCell40 sPeriod_prev_RNI43A11_LC_8_12_7 (
            .in0(N__31569),
            .in1(N__30674),
            .in2(N__22894),
            .in3(N__30888),
            .lcout(g0_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_0_LC_8_13_0.C_ON=1'b1;
    defparam sTrigCounter_0_LC_8_13_0.SEQ_MODE=4'b1000;
    defparam sTrigCounter_0_LC_8_13_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_0_LC_8_13_0 (
            .in0(_gnd_net_),
            .in1(N__26563),
            .in2(N__22877),
            .in3(N__22876),
            .lcout(sTrigCounterZ0Z_0),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(un1_sTrigCounter_cry_0),
            .clk(N__52303),
            .ce(),
            .sr(N__23084));
    defparam sTrigCounter_1_LC_8_13_1.C_ON=1'b1;
    defparam sTrigCounter_1_LC_8_13_1.SEQ_MODE=4'b1000;
    defparam sTrigCounter_1_LC_8_13_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_1_LC_8_13_1 (
            .in0(_gnd_net_),
            .in1(N__26950),
            .in2(_gnd_net_),
            .in3(N__22862),
            .lcout(sTrigCounterZ0Z_1),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_0),
            .carryout(un1_sTrigCounter_cry_1),
            .clk(N__52303),
            .ce(),
            .sr(N__23084));
    defparam sTrigCounter_2_LC_8_13_2.C_ON=1'b1;
    defparam sTrigCounter_2_LC_8_13_2.SEQ_MODE=4'b1000;
    defparam sTrigCounter_2_LC_8_13_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_2_LC_8_13_2 (
            .in0(_gnd_net_),
            .in1(N__22859),
            .in2(_gnd_net_),
            .in3(N__22847),
            .lcout(sTrigCounterZ0Z_2),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_1),
            .carryout(un1_sTrigCounter_cry_2),
            .clk(N__52303),
            .ce(),
            .sr(N__23084));
    defparam sTrigCounter_3_LC_8_13_3.C_ON=1'b1;
    defparam sTrigCounter_3_LC_8_13_3.SEQ_MODE=4'b1000;
    defparam sTrigCounter_3_LC_8_13_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_3_LC_8_13_3 (
            .in0(_gnd_net_),
            .in1(N__22844),
            .in2(_gnd_net_),
            .in3(N__22832),
            .lcout(sTrigCounterZ0Z_3),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_2),
            .carryout(un1_sTrigCounter_cry_3),
            .clk(N__52303),
            .ce(),
            .sr(N__23084));
    defparam sTrigCounter_4_LC_8_13_4.C_ON=1'b1;
    defparam sTrigCounter_4_LC_8_13_4.SEQ_MODE=4'b1000;
    defparam sTrigCounter_4_LC_8_13_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_4_LC_8_13_4 (
            .in0(_gnd_net_),
            .in1(N__23072),
            .in2(_gnd_net_),
            .in3(N__23060),
            .lcout(sTrigCounterZ0Z_4),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_3),
            .carryout(un1_sTrigCounter_cry_4),
            .clk(N__52303),
            .ce(),
            .sr(N__23084));
    defparam sTrigCounter_5_LC_8_13_5.C_ON=1'b1;
    defparam sTrigCounter_5_LC_8_13_5.SEQ_MODE=4'b1000;
    defparam sTrigCounter_5_LC_8_13_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_5_LC_8_13_5 (
            .in0(_gnd_net_),
            .in1(N__23057),
            .in2(_gnd_net_),
            .in3(N__23045),
            .lcout(sTrigCounterZ0Z_5),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_4),
            .carryout(un1_sTrigCounter_cry_5),
            .clk(N__52303),
            .ce(),
            .sr(N__23084));
    defparam sTrigCounter_6_LC_8_13_6.C_ON=1'b1;
    defparam sTrigCounter_6_LC_8_13_6.SEQ_MODE=4'b1000;
    defparam sTrigCounter_6_LC_8_13_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_6_LC_8_13_6 (
            .in0(_gnd_net_),
            .in1(N__23042),
            .in2(_gnd_net_),
            .in3(N__23030),
            .lcout(sTrigCounterZ0Z_6),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_5),
            .carryout(un1_sTrigCounter_cry_6),
            .clk(N__52303),
            .ce(),
            .sr(N__23084));
    defparam sTrigCounter_7_LC_8_13_7.C_ON=1'b1;
    defparam sTrigCounter_7_LC_8_13_7.SEQ_MODE=4'b1000;
    defparam sTrigCounter_7_LC_8_13_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_7_LC_8_13_7 (
            .in0(_gnd_net_),
            .in1(N__23027),
            .in2(_gnd_net_),
            .in3(N__23015),
            .lcout(sTrigCounterZ0Z_7),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_6),
            .carryout(un1_sTrigCounter_cry_7),
            .clk(N__52303),
            .ce(),
            .sr(N__23084));
    defparam sTrigCounter_8_LC_8_14_0.C_ON=1'b1;
    defparam sTrigCounter_8_LC_8_14_0.SEQ_MODE=4'b1000;
    defparam sTrigCounter_8_LC_8_14_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_8_LC_8_14_0 (
            .in0(_gnd_net_),
            .in1(N__23012),
            .in2(_gnd_net_),
            .in3(N__23000),
            .lcout(sTrigCounterZ0Z_8),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(un1_sTrigCounter_cry_8),
            .clk(N__52314),
            .ce(),
            .sr(N__23083));
    defparam sTrigCounter_9_LC_8_14_1.C_ON=1'b1;
    defparam sTrigCounter_9_LC_8_14_1.SEQ_MODE=4'b1000;
    defparam sTrigCounter_9_LC_8_14_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_9_LC_8_14_1 (
            .in0(_gnd_net_),
            .in1(N__22997),
            .in2(_gnd_net_),
            .in3(N__22985),
            .lcout(sTrigCounterZ0Z_9),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_8),
            .carryout(un1_sTrigCounter_cry_9),
            .clk(N__52314),
            .ce(),
            .sr(N__23083));
    defparam sTrigCounter_10_LC_8_14_2.C_ON=1'b1;
    defparam sTrigCounter_10_LC_8_14_2.SEQ_MODE=4'b1000;
    defparam sTrigCounter_10_LC_8_14_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_10_LC_8_14_2 (
            .in0(_gnd_net_),
            .in1(N__22982),
            .in2(_gnd_net_),
            .in3(N__22970),
            .lcout(sTrigCounterZ0Z_10),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_9),
            .carryout(un1_sTrigCounter_cry_10),
            .clk(N__52314),
            .ce(),
            .sr(N__23083));
    defparam sTrigCounter_11_LC_8_14_3.C_ON=1'b1;
    defparam sTrigCounter_11_LC_8_14_3.SEQ_MODE=4'b1000;
    defparam sTrigCounter_11_LC_8_14_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_11_LC_8_14_3 (
            .in0(_gnd_net_),
            .in1(N__22967),
            .in2(_gnd_net_),
            .in3(N__22955),
            .lcout(sTrigCounterZ0Z_11),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_10),
            .carryout(un1_sTrigCounter_cry_11),
            .clk(N__52314),
            .ce(),
            .sr(N__23083));
    defparam sTrigCounter_12_LC_8_14_4.C_ON=1'b1;
    defparam sTrigCounter_12_LC_8_14_4.SEQ_MODE=4'b1000;
    defparam sTrigCounter_12_LC_8_14_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_12_LC_8_14_4 (
            .in0(_gnd_net_),
            .in1(N__22952),
            .in2(_gnd_net_),
            .in3(N__23132),
            .lcout(sTrigCounterZ0Z_12),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_11),
            .carryout(un1_sTrigCounter_cry_12),
            .clk(N__52314),
            .ce(),
            .sr(N__23083));
    defparam sTrigCounter_13_LC_8_14_5.C_ON=1'b1;
    defparam sTrigCounter_13_LC_8_14_5.SEQ_MODE=4'b1000;
    defparam sTrigCounter_13_LC_8_14_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_13_LC_8_14_5 (
            .in0(_gnd_net_),
            .in1(N__23129),
            .in2(_gnd_net_),
            .in3(N__23117),
            .lcout(sTrigCounterZ0Z_13),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_12),
            .carryout(un1_sTrigCounter_cry_13),
            .clk(N__52314),
            .ce(),
            .sr(N__23083));
    defparam sTrigCounter_14_LC_8_14_6.C_ON=1'b1;
    defparam sTrigCounter_14_LC_8_14_6.SEQ_MODE=4'b1000;
    defparam sTrigCounter_14_LC_8_14_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 sTrigCounter_14_LC_8_14_6 (
            .in0(_gnd_net_),
            .in1(N__23114),
            .in2(_gnd_net_),
            .in3(N__23102),
            .lcout(sTrigCounterZ0Z_14),
            .ltout(),
            .carryin(un1_sTrigCounter_cry_13),
            .carryout(un1_sTrigCounter_cry_14),
            .clk(N__52314),
            .ce(),
            .sr(N__23083));
    defparam sTrigCounter_15_LC_8_14_7.C_ON=1'b0;
    defparam sTrigCounter_15_LC_8_14_7.SEQ_MODE=4'b1000;
    defparam sTrigCounter_15_LC_8_14_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 sTrigCounter_15_LC_8_14_7 (
            .in0(_gnd_net_),
            .in1(N__23096),
            .in2(_gnd_net_),
            .in3(N__23099),
            .lcout(sTrigCounterZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52314),
            .ce(),
            .sr(N__23083));
    defparam sDAC_mem_29_0_LC_8_15_0.C_ON=1'b0;
    defparam sDAC_mem_29_0_LC_8_15_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_0_LC_8_15_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_29_0_LC_8_15_0 (
            .in0(N__46149),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_29Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52326),
            .ce(N__23149),
            .sr(N__51674));
    defparam sDAC_mem_29_1_LC_8_15_1.C_ON=1'b0;
    defparam sDAC_mem_29_1_LC_8_15_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_1_LC_8_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_29_1_LC_8_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50883),
            .lcout(sDAC_mem_29Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52326),
            .ce(N__23149),
            .sr(N__51674));
    defparam sDAC_mem_29_2_LC_8_15_2.C_ON=1'b0;
    defparam sDAC_mem_29_2_LC_8_15_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_2_LC_8_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_29_2_LC_8_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47379),
            .lcout(sDAC_mem_29Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52326),
            .ce(N__23149),
            .sr(N__51674));
    defparam sDAC_mem_29_3_LC_8_15_3.C_ON=1'b0;
    defparam sDAC_mem_29_3_LC_8_15_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_3_LC_8_15_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_29_3_LC_8_15_3 (
            .in0(N__46650),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_29Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52326),
            .ce(N__23149),
            .sr(N__51674));
    defparam sDAC_mem_29_4_LC_8_15_4.C_ON=1'b0;
    defparam sDAC_mem_29_4_LC_8_15_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_4_LC_8_15_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_29_4_LC_8_15_4 (
            .in0(N__45574),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_29Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52326),
            .ce(N__23149),
            .sr(N__51674));
    defparam sDAC_mem_29_6_LC_8_15_6.C_ON=1'b0;
    defparam sDAC_mem_29_6_LC_8_15_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_6_LC_8_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_29_6_LC_8_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50329),
            .lcout(sDAC_mem_29Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52326),
            .ce(N__23149),
            .sr(N__51674));
    defparam sDAC_mem_29_7_LC_8_15_7.C_ON=1'b0;
    defparam sDAC_mem_29_7_LC_8_15_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_7_LC_8_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_29_7_LC_8_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50060),
            .lcout(sDAC_mem_29Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52326),
            .ce(N__23149),
            .sr(N__51674));
    defparam sDAC_mem_16_0_LC_8_16_0.C_ON=1'b0;
    defparam sDAC_mem_16_0_LC_8_16_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_0_LC_8_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_0_LC_8_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46279),
            .lcout(sDAC_mem_16Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52336),
            .ce(N__33504),
            .sr(N__51665));
    defparam sDAC_mem_16_1_LC_8_16_1.C_ON=1'b0;
    defparam sDAC_mem_16_1_LC_8_16_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_1_LC_8_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_1_LC_8_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50881),
            .lcout(sDAC_mem_16Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52336),
            .ce(N__33504),
            .sr(N__51665));
    defparam sDAC_mem_16_2_LC_8_16_2.C_ON=1'b0;
    defparam sDAC_mem_16_2_LC_8_16_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_2_LC_8_16_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_16_2_LC_8_16_2 (
            .in0(_gnd_net_),
            .in1(N__47380),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_16Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52336),
            .ce(N__33504),
            .sr(N__51665));
    defparam sEEPon_0_LC_8_17_0.C_ON=1'b0;
    defparam sEEPon_0_LC_8_17_0.SEQ_MODE=4'b1010;
    defparam sEEPon_0_LC_8_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_0_LC_8_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46280),
            .lcout(sEEPonZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52345),
            .ce(N__23207),
            .sr(N__51660));
    defparam sEEPon_1_LC_8_17_1.C_ON=1'b0;
    defparam sEEPon_1_LC_8_17_1.SEQ_MODE=4'b1010;
    defparam sEEPon_1_LC_8_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_1_LC_8_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50882),
            .lcout(sEEPonZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52345),
            .ce(N__23207),
            .sr(N__51660));
    defparam sEEPon_2_LC_8_17_2.C_ON=1'b0;
    defparam sEEPon_2_LC_8_17_2.SEQ_MODE=4'b1011;
    defparam sEEPon_2_LC_8_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_2_LC_8_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47457),
            .lcout(sEEPonZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52345),
            .ce(N__23207),
            .sr(N__51660));
    defparam sEEPon_3_LC_8_17_3.C_ON=1'b0;
    defparam sEEPon_3_LC_8_17_3.SEQ_MODE=4'b1010;
    defparam sEEPon_3_LC_8_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_3_LC_8_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46909),
            .lcout(sEEPonZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52345),
            .ce(N__23207),
            .sr(N__51660));
    defparam sEEPon_4_LC_8_17_4.C_ON=1'b0;
    defparam sEEPon_4_LC_8_17_4.SEQ_MODE=4'b1011;
    defparam sEEPon_4_LC_8_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_4_LC_8_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45575),
            .lcout(sEEPonZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52345),
            .ce(N__23207),
            .sr(N__51660));
    defparam sEEPon_5_LC_8_17_5.C_ON=1'b0;
    defparam sEEPon_5_LC_8_17_5.SEQ_MODE=4'b1010;
    defparam sEEPon_5_LC_8_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_5_LC_8_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45085),
            .lcout(sEEPonZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52345),
            .ce(N__23207),
            .sr(N__51660));
    defparam sEEPon_6_LC_8_17_6.C_ON=1'b0;
    defparam sEEPon_6_LC_8_17_6.SEQ_MODE=4'b1010;
    defparam sEEPon_6_LC_8_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_6_LC_8_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50330),
            .lcout(sEEPonZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52345),
            .ce(N__23207),
            .sr(N__51660));
    defparam sEEPon_7_LC_8_17_7.C_ON=1'b0;
    defparam sEEPon_7_LC_8_17_7.SEQ_MODE=4'b1010;
    defparam sEEPon_7_LC_8_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_7_LC_8_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49990),
            .lcout(sEEPonZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52345),
            .ce(N__23207),
            .sr(N__51660));
    defparam \spi_master_inst.spi_data_path_u1.tx_ready_i_LC_9_3_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_ready_i_LC_9_3_1 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.spi_data_path_u1.tx_ready_i_LC_9_3_1 .LUT_INIT=16'b0000000011110100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_ready_i_LC_9_3_1  (
            .in0(N__23195),
            .in1(N__23188),
            .in2(N__43888),
            .in3(N__47554),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_ready_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48451),
            .ce(),
            .sr(N__51795));
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg3_i_LC_9_3_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg3_i_LC_9_3_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg3_i_LC_9_3_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_done_reg3_i_LC_9_3_2  (
            .in0(N__23189),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48451),
            .ce(),
            .sr(N__51795));
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg2_i_LC_9_3_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg2_i_LC_9_3_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg2_i_LC_9_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_done_reg2_i_LC_9_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23159),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48451),
            .ce(),
            .sr(N__51795));
    defparam \spi_master_inst.sclk_gen_u0.spi_start_i_LC_9_3_4 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spi_start_i_LC_9_3_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.spi_start_i_LC_9_3_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spi_start_i_LC_9_3_4  (
            .in0(N__47555),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_master_inst.sclk_gen_u0.spi_start_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48451),
            .ce(),
            .sr(N__51795));
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg1_i_LC_9_3_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg1_i_LC_9_3_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg1_i_LC_9_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_done_reg1_i_LC_9_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23180),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48451),
            .ce(),
            .sr(N__51795));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_4_LC_9_3_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_4_LC_9_3_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_4_LC_9_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_4_LC_9_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31778),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48451),
            .ce(),
            .sr(N__51795));
    defparam reset_rpi_ibuf_RNIRGF52_LC_9_4_0.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNIRGF52_LC_9_4_0.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNIRGF52_LC_9_4_0.LUT_INIT=16'b0010000000000000;
    LogicCell40 reset_rpi_ibuf_RNIRGF52_LC_9_4_0 (
            .in0(N__23300),
            .in1(N__27106),
            .in2(N__49355),
            .in3(N__33768),
            .lcout(sEEADC_freq_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4Q_12_LC_9_4_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4Q_12_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4Q_12_LC_9_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4Q_12_LC_9_4_3  (
            .in0(N__25766),
            .in1(N__23234),
            .in2(_gnd_net_),
            .in3(N__24692),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4Q_10_LC_9_4_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4Q_10_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4Q_10_LC_9_4_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4Q_10_LC_9_4_5  (
            .in0(N__43847),
            .in1(N__23999),
            .in2(_gnd_net_),
            .in3(N__24691),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_10_0_LC_9_5_0.C_ON=1'b0;
    defparam sDAC_mem_10_0_LC_9_5_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_0_LC_9_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_0_LC_9_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45977),
            .lcout(sDAC_mem_10Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52337),
            .ce(N__23264),
            .sr(N__51766));
    defparam sDAC_mem_10_1_LC_9_5_1.C_ON=1'b0;
    defparam sDAC_mem_10_1_LC_9_5_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_1_LC_9_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_1_LC_9_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50715),
            .lcout(sDAC_mem_10Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52337),
            .ce(N__23264),
            .sr(N__51766));
    defparam sDAC_mem_10_2_LC_9_5_2.C_ON=1'b0;
    defparam sDAC_mem_10_2_LC_9_5_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_2_LC_9_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_2_LC_9_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47118),
            .lcout(sDAC_mem_10Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52337),
            .ce(N__23264),
            .sr(N__51766));
    defparam sDAC_mem_10_3_LC_9_5_3.C_ON=1'b0;
    defparam sDAC_mem_10_3_LC_9_5_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_3_LC_9_5_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_10_3_LC_9_5_3 (
            .in0(N__46518),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_10Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52337),
            .ce(N__23264),
            .sr(N__51766));
    defparam sDAC_mem_10_4_LC_9_5_4.C_ON=1'b0;
    defparam sDAC_mem_10_4_LC_9_5_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_4_LC_9_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_4_LC_9_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45224),
            .lcout(sDAC_mem_10Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52337),
            .ce(N__23264),
            .sr(N__51766));
    defparam sDAC_mem_10_5_LC_9_5_5.C_ON=1'b0;
    defparam sDAC_mem_10_5_LC_9_5_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_5_LC_9_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_5_LC_9_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44730),
            .lcout(sDAC_mem_10Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52337),
            .ce(N__23264),
            .sr(N__51766));
    defparam sDAC_mem_10_6_LC_9_5_6.C_ON=1'b0;
    defparam sDAC_mem_10_6_LC_9_5_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_6_LC_9_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_6_LC_9_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50224),
            .lcout(sDAC_mem_10Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52337),
            .ce(N__23264),
            .sr(N__51766));
    defparam sDAC_mem_10_7_LC_9_5_7.C_ON=1'b0;
    defparam sDAC_mem_10_7_LC_9_5_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_7_LC_9_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_7_LC_9_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49654),
            .lcout(sDAC_mem_10Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52337),
            .ce(N__23264),
            .sr(N__51766));
    defparam sDAC_mem_38_0_LC_9_6_0.C_ON=1'b0;
    defparam sDAC_mem_38_0_LC_9_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_0_LC_9_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_0_LC_9_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45979),
            .lcout(sDAC_mem_38Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52327),
            .ce(N__23246),
            .sr(N__51753));
    defparam sDAC_mem_38_1_LC_9_6_1.C_ON=1'b0;
    defparam sDAC_mem_38_1_LC_9_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_1_LC_9_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_1_LC_9_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50718),
            .lcout(sDAC_mem_38Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52327),
            .ce(N__23246),
            .sr(N__51753));
    defparam sDAC_mem_38_2_LC_9_6_2.C_ON=1'b0;
    defparam sDAC_mem_38_2_LC_9_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_2_LC_9_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_2_LC_9_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47121),
            .lcout(sDAC_mem_38Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52327),
            .ce(N__23246),
            .sr(N__51753));
    defparam sDAC_mem_38_3_LC_9_6_3.C_ON=1'b0;
    defparam sDAC_mem_38_3_LC_9_6_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_3_LC_9_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_3_LC_9_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46521),
            .lcout(sDAC_mem_38Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52327),
            .ce(N__23246),
            .sr(N__51753));
    defparam sDAC_mem_38_4_LC_9_6_4.C_ON=1'b0;
    defparam sDAC_mem_38_4_LC_9_6_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_4_LC_9_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_4_LC_9_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45226),
            .lcout(sDAC_mem_38Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52327),
            .ce(N__23246),
            .sr(N__51753));
    defparam sDAC_mem_38_5_LC_9_6_5.C_ON=1'b0;
    defparam sDAC_mem_38_5_LC_9_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_5_LC_9_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_5_LC_9_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44733),
            .lcout(sDAC_mem_38Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52327),
            .ce(N__23246),
            .sr(N__51753));
    defparam sDAC_mem_38_6_LC_9_6_6.C_ON=1'b0;
    defparam sDAC_mem_38_6_LC_9_6_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_6_LC_9_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_6_LC_9_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50170),
            .lcout(sDAC_mem_38Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52327),
            .ce(N__23246),
            .sr(N__51753));
    defparam sDAC_mem_38_7_LC_9_6_7.C_ON=1'b0;
    defparam sDAC_mem_38_7_LC_9_6_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_7_LC_9_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_7_LC_9_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49672),
            .lcout(sDAC_mem_38Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52327),
            .ce(N__23246),
            .sr(N__51753));
    defparam sAddress_RNI9IH12_12_5_LC_9_7_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_12_5_LC_9_7_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_12_5_LC_9_7_0.LUT_INIT=16'b0010000000000000;
    LogicCell40 sAddress_RNI9IH12_12_5_LC_9_7_0 (
            .in0(N__40298),
            .in1(N__40961),
            .in2(N__23298),
            .in3(N__40785),
            .lcout(sDAC_mem_14_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_5_5_LC_9_7_1.C_ON=1'b0;
    defparam sAddress_RNI9IH12_5_5_LC_9_7_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_5_5_LC_9_7_1.LUT_INIT=16'b0000000010000000;
    LogicCell40 sAddress_RNI9IH12_5_5_LC_9_7_1 (
            .in0(N__40786),
            .in1(N__23293),
            .in2(N__40995),
            .in3(N__40300),
            .lcout(sDAC_mem_38_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_17_5_LC_9_7_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_17_5_LC_9_7_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_17_5_LC_9_7_2.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNI9IH12_17_5_LC_9_7_2 (
            .in0(N__40296),
            .in1(N__40960),
            .in2(N__23299),
            .in3(N__40784),
            .lcout(sDAC_mem_6_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_3_3_LC_9_7_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_3_3_LC_9_7_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_3_3_LC_9_7_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 sAddress_RNI9IH12_3_3_LC_9_7_3 (
            .in0(N__23294),
            .in1(N__40299),
            .in2(_gnd_net_),
            .in3(N__39997),
            .lcout(sDAC_mem_30_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI6VH7_3_1_LC_9_7_4.C_ON=1'b0;
    defparam sAddress_RNI6VH7_3_1_LC_9_7_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI6VH7_3_1_LC_9_7_4.LUT_INIT=16'b0000110000000000;
    LogicCell40 sAddress_RNI6VH7_3_1_LC_9_7_4 (
            .in0(_gnd_net_),
            .in1(N__40120),
            .in2(N__40532),
            .in3(N__40603),
            .lcout(sAddress_RNI6VH7_3Z0Z_1),
            .ltout(sAddress_RNI6VH7_3Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_7_3_LC_9_7_5.C_ON=1'b0;
    defparam sAddress_RNI9IH12_7_3_LC_9_7_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_7_3_LC_9_7_5.LUT_INIT=16'b0011000000000000;
    LogicCell40 sAddress_RNI9IH12_7_3_LC_9_7_5 (
            .in0(_gnd_net_),
            .in1(N__40297),
            .in2(N__23267),
            .in3(N__39998),
            .lcout(sDAC_mem_22_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_0_LC_9_7_6.C_ON=1'b0;
    defparam sAddress_0_LC_9_7_6.SEQ_MODE=4'b1010;
    defparam sAddress_0_LC_9_7_6.LUT_INIT=16'b0000000011001100;
    LogicCell40 sAddress_0_LC_9_7_6 (
            .in0(_gnd_net_),
            .in1(N__46015),
            .in2(_gnd_net_),
            .in3(N__26165),
            .lcout(sAddressZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52315),
            .ce(N__23418),
            .sr(N__51740));
    defparam sAddress_RNI6VH7_0_1_LC_9_7_7.C_ON=1'b0;
    defparam sAddress_RNI6VH7_0_1_LC_9_7_7.SEQ_MODE=4'b0000;
    defparam sAddress_RNI6VH7_0_1_LC_9_7_7.LUT_INIT=16'b1111101111111011;
    LogicCell40 sAddress_RNI6VH7_0_1_LC_9_7_7 (
            .in0(N__40604),
            .in1(N__40516),
            .in2(N__40157),
            .in3(_gnd_net_),
            .lcout(N_333),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_16_5_LC_9_8_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_16_5_LC_9_8_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_16_5_LC_9_8_0.LUT_INIT=16'b0000001000000000;
    LogicCell40 sAddress_RNI9IH12_16_5_LC_9_8_0 (
            .in0(N__40302),
            .in1(N__40968),
            .in2(N__23834),
            .in3(N__40794),
            .lcout(sDAC_mem_10_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI6VH7_1_LC_9_8_1.C_ON=1'b0;
    defparam sAddress_RNI6VH7_1_LC_9_8_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI6VH7_1_LC_9_8_1.LUT_INIT=16'b1110111011111111;
    LogicCell40 sAddress_RNI6VH7_1_LC_9_8_1 (
            .in0(N__40615),
            .in1(N__40520),
            .in2(_gnd_net_),
            .in3(N__40139),
            .lcout(N_326),
            .ltout(N_326_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_10_3_LC_9_8_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_10_3_LC_9_8_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_10_3_LC_9_8_2.LUT_INIT=16'b0000001100000000;
    LogicCell40 sAddress_RNI9IH12_10_3_LC_9_8_2 (
            .in0(_gnd_net_),
            .in1(N__40301),
            .in2(N__23249),
            .in3(N__40002),
            .lcout(sDAC_mem_18_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_2_5_LC_9_8_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_2_5_LC_9_8_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_2_5_LC_9_8_3.LUT_INIT=16'b0010000000000000;
    LogicCell40 sAddress_RNI9IH12_2_5_LC_9_8_3 (
            .in0(N__40796),
            .in1(N__23824),
            .in2(N__40997),
            .in3(N__40305),
            .lcout(sDAC_mem_42_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_8_5_LC_9_8_4.C_ON=1'b0;
    defparam sAddress_RNI9IH12_8_5_LC_9_8_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_8_5_LC_9_8_4.LUT_INIT=16'b0000010000000000;
    LogicCell40 sAddress_RNI9IH12_8_5_LC_9_8_4 (
            .in0(N__40304),
            .in1(N__40969),
            .in2(N__23835),
            .in3(N__40795),
            .lcout(sDAC_mem_34_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_20_5_LC_9_8_5.C_ON=1'b0;
    defparam sAddress_RNI9IH12_20_5_LC_9_8_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_20_5_LC_9_8_5.LUT_INIT=16'b0000000000000010;
    LogicCell40 sAddress_RNI9IH12_20_5_LC_9_8_5 (
            .in0(N__40793),
            .in1(N__23823),
            .in2(N__40996),
            .in3(N__40303),
            .lcout(sDAC_mem_2_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_2_LC_9_8_7.C_ON=1'b0;
    defparam sAddress_2_LC_9_8_7.SEQ_MODE=4'b1010;
    defparam sAddress_2_LC_9_8_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 sAddress_2_LC_9_8_7 (
            .in0(_gnd_net_),
            .in1(N__47174),
            .in2(_gnd_net_),
            .in3(N__26164),
            .lcout(sAddressZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52304),
            .ce(N__23422),
            .sr(N__51726));
    defparam sAddress_RNI6VH7_5_1_LC_9_9_0.C_ON=1'b0;
    defparam sAddress_RNI6VH7_5_1_LC_9_9_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI6VH7_5_1_LC_9_9_0.LUT_INIT=16'b0100010000000000;
    LogicCell40 sAddress_RNI6VH7_5_1_LC_9_9_0 (
            .in0(N__40616),
            .in1(N__40507),
            .in2(_gnd_net_),
            .in3(N__40158),
            .lcout(sAddress_RNI6VH7_5Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_ready_i_RNIBLID_LC_9_9_1 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_ready_i_RNIBLID_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_ready_i_RNIBLID_LC_9_9_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \spi_slave_inst.tx_ready_i_RNIBLID_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__49365),
            .in2(_gnd_net_),
            .in3(N__44570),
            .lcout(\spi_slave_inst.un4_i_wr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_14_5_LC_9_9_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_14_5_LC_9_9_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_14_5_LC_9_9_2.LUT_INIT=16'b0000000000001000;
    LogicCell40 sAddress_RNI9IH12_14_5_LC_9_9_2 (
            .in0(N__40746),
            .in1(N__40385),
            .in2(N__40994),
            .in3(N__23550),
            .lcout(sDAC_mem_15_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LED_ACQ_obuf_RNO_LC_9_9_3.C_ON=1'b0;
    defparam LED_ACQ_obuf_RNO_LC_9_9_3.SEQ_MODE=4'b0000;
    defparam LED_ACQ_obuf_RNO_LC_9_9_3.LUT_INIT=16'b1100110000000100;
    LogicCell40 LED_ACQ_obuf_RNO_LC_9_9_3 (
            .in0(N__25158),
            .in1(N__49364),
            .in2(N__25187),
            .in3(N__25213),
            .lcout(LED_ACQ_obuf_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_1_2_LC_9_9_4.C_ON=1'b0;
    defparam sAddress_RNI9IH12_1_2_LC_9_9_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_1_2_LC_9_9_4.LUT_INIT=16'b0010000000000000;
    LogicCell40 sAddress_RNI9IH12_1_2_LC_9_9_4 (
            .in0(N__40618),
            .in1(N__23463),
            .in2(N__27023),
            .in3(N__33743),
            .lcout(sAddress_RNI9IH12_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_2_LC_9_9_5.C_ON=1'b0;
    defparam sAddress_RNI9IH12_2_LC_9_9_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_2_LC_9_9_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 sAddress_RNI9IH12_2_LC_9_9_5 (
            .in0(N__27015),
            .in1(N__40619),
            .in2(_gnd_net_),
            .in3(N__39973),
            .lcout(sDAC_mem_24_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIAM2A_0_1_LC_9_9_6.C_ON=1'b0;
    defparam sAddress_RNIAM2A_0_1_LC_9_9_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNIAM2A_0_1_LC_9_9_6.LUT_INIT=16'b0000000000000010;
    LogicCell40 sAddress_RNIAM2A_0_1_LC_9_9_6 (
            .in0(N__40617),
            .in1(N__40508),
            .in2(N__40377),
            .in3(N__40159),
            .lcout(sAddress_RNIAM2A_0Z0Z_1),
            .ltout(sAddress_RNIAM2A_0Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_3_5_LC_9_9_7.C_ON=1'b0;
    defparam sAddress_RNI9IH12_3_5_LC_9_9_7.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_3_5_LC_9_9_7.LUT_INIT=16'b0011000000000000;
    LogicCell40 sAddress_RNI9IH12_3_5_LC_9_9_7 (
            .in0(_gnd_net_),
            .in1(N__40956),
            .in2(N__23501),
            .in3(N__40745),
            .lcout(sDAC_mem_5_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIAM2A_1_LC_9_10_0.C_ON=1'b0;
    defparam sAddress_RNIAM2A_1_LC_9_10_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNIAM2A_1_LC_9_10_0.LUT_INIT=16'b0000000100100000;
    LogicCell40 sAddress_RNIAM2A_1_LC_9_10_0 (
            .in0(N__40161),
            .in1(N__40334),
            .in2(N__40521),
            .in3(N__40646),
            .lcout(N_445),
            .ltout(N_445_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_0_LC_9_10_1.C_ON=1'b0;
    defparam sAddress_RNIA6242_0_LC_9_10_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_0_LC_9_10_1.LUT_INIT=16'b0010000000000000;
    LogicCell40 sAddress_RNIA6242_0_LC_9_10_1 (
            .in0(N__40162),
            .in1(N__23462),
            .in2(N__23498),
            .in3(N__33745),
            .lcout(sAddress_RNIA6242Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_13_5_LC_9_10_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_13_5_LC_9_10_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_13_5_LC_9_10_2.LUT_INIT=16'b0010000000000000;
    LogicCell40 sAddress_RNI9IH12_13_5_LC_9_10_2 (
            .in0(N__40336),
            .in1(N__40949),
            .in2(N__23495),
            .in3(N__40741),
            .lcout(sDAC_mem_12_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_2_3_LC_9_10_4.C_ON=1'b0;
    defparam sAddress_RNI9IH12_2_3_LC_9_10_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_2_3_LC_9_10_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 sAddress_RNI9IH12_2_3_LC_9_10_4 (
            .in0(N__23494),
            .in1(N__40335),
            .in2(_gnd_net_),
            .in3(N__39972),
            .lcout(sDAC_mem_28_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_4_0_LC_9_10_5.C_ON=1'b0;
    defparam sAddress_RNIA6242_4_0_LC_9_10_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_4_0_LC_9_10_5.LUT_INIT=16'b0000010000000000;
    LogicCell40 sAddress_RNIA6242_4_0_LC_9_10_5 (
            .in0(N__40163),
            .in1(N__23474),
            .in2(N__23468),
            .in3(N__33746),
            .lcout(sAddress_RNIA6242_4Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_1_LC_9_10_6.C_ON=1'b0;
    defparam sAddress_1_LC_9_10_6.SEQ_MODE=4'b1010;
    defparam sAddress_1_LC_9_10_6.LUT_INIT=16'b0000000011001100;
    LogicCell40 sAddress_1_LC_9_10_6 (
            .in0(_gnd_net_),
            .in1(N__50851),
            .in2(_gnd_net_),
            .in3(N__26196),
            .lcout(sAddressZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52282),
            .ce(N__23409),
            .sr(N__51703));
    defparam sAddress_RNI6VH7_2_1_LC_9_10_7.C_ON=1'b0;
    defparam sAddress_RNI6VH7_2_1_LC_9_10_7.SEQ_MODE=4'b0000;
    defparam sAddress_RNI6VH7_2_1_LC_9_10_7.LUT_INIT=16'b1000100000000000;
    LogicCell40 sAddress_RNI6VH7_2_1_LC_9_10_7 (
            .in0(N__40645),
            .in1(N__40496),
            .in2(_gnd_net_),
            .in3(N__40160),
            .lcout(sAddress_RNI6VH7_2Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIM4BU_20_LC_9_11_0.C_ON=1'b0;
    defparam sCounter_RNIM4BU_20_LC_9_11_0.SEQ_MODE=4'b0000;
    defparam sCounter_RNIM4BU_20_LC_9_11_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNIM4BU_20_LC_9_11_0 (
            .in0(N__33362),
            .in1(N__29872),
            .in2(N__33165),
            .in3(N__29998),
            .lcout(g0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigInternal_prev_RNIH3OJ1_LC_9_11_2.C_ON=1'b0;
    defparam sEETrigInternal_prev_RNIH3OJ1_LC_9_11_2.SEQ_MODE=4'b0000;
    defparam sEETrigInternal_prev_RNIH3OJ1_LC_9_11_2.LUT_INIT=16'b1111111111000100;
    LogicCell40 sEETrigInternal_prev_RNIH3OJ1_LC_9_11_2 (
            .in0(N__23718),
            .in1(N__23666),
            .in2(N__23657),
            .in3(N__31029),
            .lcout(sEETrigInternal_prev_RNIH3OJZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sSingleCont_RNIUP5M_LC_9_11_3.C_ON=1'b0;
    defparam sSingleCont_RNIUP5M_LC_9_11_3.SEQ_MODE=4'b0000;
    defparam sSingleCont_RNIUP5M_LC_9_11_3.LUT_INIT=16'b0010001000000000;
    LogicCell40 sSingleCont_RNIUP5M_LC_9_11_3 (
            .in0(N__49253),
            .in1(N__30555),
            .in2(_gnd_net_),
            .in3(N__23606),
            .lcout(g0_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_4_3_LC_9_11_4.C_ON=1'b0;
    defparam sAddress_RNI9IH12_4_3_LC_9_11_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_4_3_LC_9_11_4.LUT_INIT=16'b0000000010001000;
    LogicCell40 sAddress_RNI9IH12_4_3_LC_9_11_4 (
            .in0(N__39991),
            .in1(N__40384),
            .in2(_gnd_net_),
            .in3(N__34867),
            .lcout(sDAC_mem_27_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIUB4L_12_LC_9_11_5.C_ON=1'b0;
    defparam sCounter_RNIUB4L_12_LC_9_11_5.SEQ_MODE=4'b0000;
    defparam sCounter_RNIUB4L_12_LC_9_11_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNIUB4L_12_LC_9_11_5 (
            .in0(N__31722),
            .in1(N__31550),
            .in2(N__31468),
            .in3(N__31643),
            .lcout(N_831_16),
            .ltout(N_831_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIP69T1_10_LC_9_11_6.C_ON=1'b0;
    defparam sCounter_RNIP69T1_10_LC_9_11_6.SEQ_MODE=4'b0000;
    defparam sCounter_RNIP69T1_10_LC_9_11_6.LUT_INIT=16'b1111111111101111;
    LogicCell40 sCounter_RNIP69T1_10_LC_9_11_6 (
            .in0(N__24182),
            .in1(N__33053),
            .in2(N__23570),
            .in3(N__30345),
            .lcout(un1_reset_rpi_inv_2_0_o2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_5_3_LC_9_12_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_5_3_LC_9_12_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_5_3_LC_9_12_0.LUT_INIT=16'b0010000000100000;
    LogicCell40 sAddress_RNI9IH12_5_3_LC_9_12_0 (
            .in0(N__40009),
            .in1(N__23567),
            .in2(N__40412),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_31_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIEQR21_10_LC_9_12_1.C_ON=1'b0;
    defparam sCounter_RNIEQR21_10_LC_9_12_1.SEQ_MODE=4'b0000;
    defparam sCounter_RNIEQR21_10_LC_9_12_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNIEQR21_10_LC_9_12_1 (
            .in0(N__30457),
            .in1(N__30563),
            .in2(N__30361),
            .in3(N__30233),
            .lcout(),
            .ltout(g0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNID5AA2_5_LC_9_12_2.C_ON=1'b0;
    defparam sCounter_RNID5AA2_5_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam sCounter_RNID5AA2_5_LC_9_12_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNID5AA2_5_LC_9_12_2 (
            .in0(N__24161),
            .in1(N__30781),
            .in2(N__23519),
            .in3(N__30898),
            .lcout(g0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIN61V1_10_LC_9_12_3.C_ON=1'b0;
    defparam sCounter_RNIN61V1_10_LC_9_12_3.SEQ_MODE=4'b0000;
    defparam sCounter_RNIN61V1_10_LC_9_12_3.LUT_INIT=16'b0000000000100000;
    LogicCell40 sCounter_RNIN61V1_10_LC_9_12_3 (
            .in0(N__24173),
            .in1(N__30346),
            .in2(N__23516),
            .in3(N__30458),
            .lcout(g0_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNI3LAJ2_1_LC_9_12_5.C_ON=1'b0;
    defparam sCounter_RNI3LAJ2_1_LC_9_12_5.SEQ_MODE=4'b0000;
    defparam sCounter_RNI3LAJ2_1_LC_9_12_5.LUT_INIT=16'b0000000000100000;
    LogicCell40 sCounter_RNI3LAJ2_1_LC_9_12_5 (
            .in0(N__24566),
            .in1(N__29873),
            .in2(N__23858),
            .in3(N__30111),
            .lcout(g0_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_6_3_LC_9_12_6.C_ON=1'b0;
    defparam sAddress_RNI9IH12_6_3_LC_9_12_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_6_3_LC_9_12_6.LUT_INIT=16'b0010000000100000;
    LogicCell40 sAddress_RNI9IH12_6_3_LC_9_12_6 (
            .in0(N__40010),
            .in1(N__23840),
            .in2(N__40411),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_26_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIDCVE1_18_LC_9_12_7.C_ON=1'b0;
    defparam sCounter_RNIDCVE1_18_LC_9_12_7.SEQ_MODE=4'b0000;
    defparam sCounter_RNIDCVE1_18_LC_9_12_7.LUT_INIT=16'b0000000000100000;
    LogicCell40 sCounter_RNIDCVE1_18_LC_9_12_7 (
            .in0(N__25850),
            .in1(N__31163),
            .in2(N__32951),
            .in3(N__30005),
            .lcout(g0_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNITBBU_23_LC_9_13_0.C_ON=1'b0;
    defparam sCounter_RNITBBU_23_LC_9_13_0.SEQ_MODE=4'b0000;
    defparam sCounter_RNITBBU_23_LC_9_13_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNITBBU_23_LC_9_13_0 (
            .in0(N__32045),
            .in1(N__30667),
            .in2(N__31930),
            .in3(N__30110),
            .lcout(g1_i_a4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIES4L_0_16_LC_9_13_1.C_ON=1'b0;
    defparam sCounter_RNIES4L_0_16_LC_9_13_1.SEQ_MODE=4'b0000;
    defparam sCounter_RNIES4L_0_16_LC_9_13_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNIES4L_0_16_LC_9_13_1 (
            .in0(N__31161),
            .in1(N__31276),
            .in2(N__33276),
            .in3(N__31366),
            .lcout(),
            .ltout(g1_i_a4_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNI2KI53_16_LC_9_13_2.C_ON=1'b0;
    defparam sCounter_RNI2KI53_16_LC_9_13_2.SEQ_MODE=4'b0000;
    defparam sCounter_RNI2KI53_16_LC_9_13_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 sCounter_RNI2KI53_16_LC_9_13_2 (
            .in0(N__24314),
            .in1(N__23792),
            .in2(N__23786),
            .in3(N__25712),
            .lcout(),
            .ltout(g1_i_a4_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_rpi_ibuf_RNIUSHQ6_LC_9_13_3.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNIUSHQ6_LC_9_13_3.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNIUSHQ6_LC_9_13_3.LUT_INIT=16'b0111010101010101;
    LogicCell40 reset_rpi_ibuf_RNIUSHQ6_LC_9_13_3 (
            .in0(N__49116),
            .in1(N__23783),
            .in2(N__23774),
            .in3(N__23771),
            .lcout(g0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIRQR25_18_LC_9_13_4.C_ON=1'b0;
    defparam sCounter_RNIRQR25_18_LC_9_13_4.SEQ_MODE=4'b0000;
    defparam sCounter_RNIRQR25_18_LC_9_13_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNIRQR25_18_LC_9_13_4 (
            .in0(N__24575),
            .in1(N__23747),
            .in2(N__23741),
            .in3(N__23726),
            .lcout(N_106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIKSV41_18_LC_9_13_7.C_ON=1'b0;
    defparam sCounter_RNIKSV41_18_LC_9_13_7.SEQ_MODE=4'b0000;
    defparam sCounter_RNIKSV41_18_LC_9_13_7.LUT_INIT=16'b1111111111111011;
    LogicCell40 sCounter_RNIKSV41_18_LC_9_13_7 (
            .in0(N__31160),
            .in1(N__24136),
            .in2(N__33275),
            .in3(N__33048),
            .lcout(g0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_26_0_LC_9_14_0.C_ON=1'b0;
    defparam sDAC_mem_26_0_LC_9_14_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_0_LC_9_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_26_0_LC_9_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46343),
            .lcout(sDAC_mem_26Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52305),
            .ce(N__28045),
            .sr(N__51675));
    defparam sDAC_mem_26_1_LC_9_14_1.C_ON=1'b0;
    defparam sDAC_mem_26_1_LC_9_14_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_1_LC_9_14_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_26_1_LC_9_14_1 (
            .in0(N__51069),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_26Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52305),
            .ce(N__28045),
            .sr(N__51675));
    defparam sDAC_mem_26_3_LC_9_14_2.C_ON=1'b0;
    defparam sDAC_mem_26_3_LC_9_14_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_3_LC_9_14_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_26_3_LC_9_14_2 (
            .in0(N__46866),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_26Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52305),
            .ce(N__28045),
            .sr(N__51675));
    defparam sDAC_mem_26_4_LC_9_14_3.C_ON=1'b0;
    defparam sDAC_mem_26_4_LC_9_14_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_4_LC_9_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_26_4_LC_9_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45577),
            .lcout(sDAC_mem_26Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52305),
            .ce(N__28045),
            .sr(N__51675));
    defparam sDAC_mem_26_6_LC_9_14_4.C_ON=1'b0;
    defparam sDAC_mem_26_6_LC_9_14_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_6_LC_9_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_26_6_LC_9_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50495),
            .lcout(sDAC_mem_26Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52305),
            .ce(N__28045),
            .sr(N__51675));
    defparam sDAC_mem_26_7_LC_9_14_5.C_ON=1'b0;
    defparam sDAC_mem_26_7_LC_9_14_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_7_LC_9_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_26_7_LC_9_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49875),
            .lcout(sDAC_mem_26Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52305),
            .ce(N__28045),
            .sr(N__51675));
    defparam sDAC_mem_30_0_LC_9_15_0.C_ON=1'b0;
    defparam sDAC_mem_30_0_LC_9_15_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_0_LC_9_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_0_LC_9_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46148),
            .lcout(sDAC_mem_30Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52316),
            .ce(N__23921),
            .sr(N__51666));
    defparam sDAC_mem_30_1_LC_9_15_1.C_ON=1'b0;
    defparam sDAC_mem_30_1_LC_9_15_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_1_LC_9_15_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_30_1_LC_9_15_1 (
            .in0(N__51039),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_30Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52316),
            .ce(N__23921),
            .sr(N__51666));
    defparam sDAC_mem_30_2_LC_9_15_2.C_ON=1'b0;
    defparam sDAC_mem_30_2_LC_9_15_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_2_LC_9_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_2_LC_9_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47363),
            .lcout(sDAC_mem_30Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52316),
            .ce(N__23921),
            .sr(N__51666));
    defparam sDAC_mem_30_3_LC_9_15_3.C_ON=1'b0;
    defparam sDAC_mem_30_3_LC_9_15_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_3_LC_9_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_3_LC_9_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46908),
            .lcout(sDAC_mem_30Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52316),
            .ce(N__23921),
            .sr(N__51666));
    defparam sDAC_mem_30_4_LC_9_15_4.C_ON=1'b0;
    defparam sDAC_mem_30_4_LC_9_15_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_4_LC_9_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_4_LC_9_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45578),
            .lcout(sDAC_mem_30Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52316),
            .ce(N__23921),
            .sr(N__51666));
    defparam sDAC_mem_30_5_LC_9_15_5.C_ON=1'b0;
    defparam sDAC_mem_30_5_LC_9_15_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_5_LC_9_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_5_LC_9_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45096),
            .lcout(sDAC_mem_30Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52316),
            .ce(N__23921),
            .sr(N__51666));
    defparam sDAC_mem_30_6_LC_9_15_6.C_ON=1'b0;
    defparam sDAC_mem_30_6_LC_9_15_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_6_LC_9_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_6_LC_9_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50528),
            .lcout(sDAC_mem_30Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52316),
            .ce(N__23921),
            .sr(N__51666));
    defparam sDAC_mem_30_7_LC_9_15_7.C_ON=1'b0;
    defparam sDAC_mem_30_7_LC_9_15_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_7_LC_9_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_7_LC_9_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49876),
            .lcout(sDAC_mem_30Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52316),
            .ce(N__23921),
            .sr(N__51666));
    defparam sCounter_RNIQB8L_23_LC_9_16_5.C_ON=1'b0;
    defparam sCounter_RNIQB8L_23_LC_9_16_5.SEQ_MODE=4'b0000;
    defparam sCounter_RNIQB8L_23_LC_9_16_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNIQB8L_23_LC_9_16_5 (
            .in0(N__32046),
            .in1(N__33161),
            .in2(N__31937),
            .in3(N__33376),
            .lcout(un21_trig_prev_21_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_0_c_inv_LC_9_17_0.C_ON=1'b1;
    defparam un7_spon_cry_0_c_inv_LC_9_17_0.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_0_c_inv_LC_9_17_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 un7_spon_cry_0_c_inv_LC_9_17_0 (
            .in0(N__23909),
            .in1(N__30241),
            .in2(N__23903),
            .in3(_gnd_net_),
            .lcout(sEEPon_i_0),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(un7_spon_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_1_c_inv_LC_9_17_1.C_ON=1'b1;
    defparam un7_spon_cry_1_c_inv_LC_9_17_1.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_1_c_inv_LC_9_17_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un7_spon_cry_1_c_inv_LC_9_17_1 (
            .in0(_gnd_net_),
            .in1(N__23888),
            .in2(N__30130),
            .in3(N__23894),
            .lcout(sEEPon_i_1),
            .ltout(),
            .carryin(un7_spon_cry_0),
            .carryout(un7_spon_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_2_c_inv_LC_9_17_2.C_ON=1'b1;
    defparam un7_spon_cry_2_c_inv_LC_9_17_2.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_2_c_inv_LC_9_17_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 un7_spon_cry_2_c_inv_LC_9_17_2 (
            .in0(N__23882),
            .in1(N__23876),
            .in2(N__30013),
            .in3(_gnd_net_),
            .lcout(sEEPon_i_2),
            .ltout(),
            .carryin(un7_spon_cry_1),
            .carryout(un7_spon_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_3_c_inv_LC_9_17_3.C_ON=1'b1;
    defparam un7_spon_cry_3_c_inv_LC_9_17_3.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_3_c_inv_LC_9_17_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 un7_spon_cry_3_c_inv_LC_9_17_3 (
            .in0(N__23870),
            .in1(N__23864),
            .in2(N__29885),
            .in3(_gnd_net_),
            .lcout(sEEPon_i_3),
            .ltout(),
            .carryin(un7_spon_cry_2),
            .carryout(un7_spon_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_4_c_inv_LC_9_17_4.C_ON=1'b1;
    defparam un7_spon_cry_4_c_inv_LC_9_17_4.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_4_c_inv_LC_9_17_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un7_spon_cry_4_c_inv_LC_9_17_4 (
            .in0(_gnd_net_),
            .in1(N__23963),
            .in2(N__31061),
            .in3(N__23969),
            .lcout(sEEPon_i_4),
            .ltout(),
            .carryin(un7_spon_cry_3),
            .carryout(un7_spon_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_5_c_inv_LC_9_17_5.C_ON=1'b1;
    defparam un7_spon_cry_5_c_inv_LC_9_17_5.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_5_c_inv_LC_9_17_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 un7_spon_cry_5_c_inv_LC_9_17_5 (
            .in0(N__23957),
            .in1(N__23951),
            .in2(N__30907),
            .in3(_gnd_net_),
            .lcout(sEEPon_i_5),
            .ltout(),
            .carryin(un7_spon_cry_4),
            .carryout(un7_spon_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_6_c_inv_LC_9_17_6.C_ON=1'b1;
    defparam un7_spon_cry_6_c_inv_LC_9_17_6.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_6_c_inv_LC_9_17_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un7_spon_cry_6_c_inv_LC_9_17_6 (
            .in0(N__23945),
            .in1(N__23939),
            .in2(N__30790),
            .in3(_gnd_net_),
            .lcout(sEEPon_i_6),
            .ltout(),
            .carryin(un7_spon_cry_5),
            .carryout(un7_spon_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_7_c_inv_LC_9_17_7.C_ON=1'b1;
    defparam un7_spon_cry_7_c_inv_LC_9_17_7.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_7_c_inv_LC_9_17_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un7_spon_cry_7_c_inv_LC_9_17_7 (
            .in0(N__23933),
            .in1(N__23927),
            .in2(N__30682),
            .in3(_gnd_net_),
            .lcout(sEEPon_i_7),
            .ltout(),
            .carryin(un7_spon_cry_6),
            .carryout(un7_spon_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_8_c_LC_9_18_0.C_ON=1'b1;
    defparam un7_spon_cry_8_c_LC_9_18_0.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_8_c_LC_9_18_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_8_c_LC_9_18_0 (
            .in0(_gnd_net_),
            .in1(N__52684),
            .in2(N__30575),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(un7_spon_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_9_c_LC_9_18_1.C_ON=1'b1;
    defparam un7_spon_cry_9_c_LC_9_18_1.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_9_c_LC_9_18_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_9_c_LC_9_18_1 (
            .in0(_gnd_net_),
            .in1(N__30466),
            .in2(N__52746),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_8),
            .carryout(un7_spon_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_10_c_LC_9_18_2.C_ON=1'b1;
    defparam un7_spon_cry_10_c_LC_9_18_2.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_10_c_LC_9_18_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_10_c_LC_9_18_2 (
            .in0(_gnd_net_),
            .in1(N__52672),
            .in2(N__30362),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_9),
            .carryout(un7_spon_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_11_c_LC_9_18_3.C_ON=1'b1;
    defparam un7_spon_cry_11_c_LC_9_18_3.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_11_c_LC_9_18_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_11_c_LC_9_18_3 (
            .in0(_gnd_net_),
            .in1(N__33058),
            .in2(N__52743),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_10),
            .carryout(un7_spon_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_12_c_LC_9_18_4.C_ON=1'b1;
    defparam un7_spon_cry_12_c_LC_9_18_4.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_12_c_LC_9_18_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_12_c_LC_9_18_4 (
            .in0(_gnd_net_),
            .in1(N__52676),
            .in2(N__31748),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_11),
            .carryout(un7_spon_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_13_c_LC_9_18_5.C_ON=1'b1;
    defparam un7_spon_cry_13_c_LC_9_18_5.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_13_c_LC_9_18_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_13_c_LC_9_18_5 (
            .in0(_gnd_net_),
            .in1(N__31660),
            .in2(N__52744),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_12),
            .carryout(un7_spon_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_14_c_LC_9_18_6.C_ON=1'b1;
    defparam un7_spon_cry_14_c_LC_9_18_6.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_14_c_LC_9_18_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_14_c_LC_9_18_6 (
            .in0(_gnd_net_),
            .in1(N__52680),
            .in2(N__31580),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_13),
            .carryout(un7_spon_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_15_c_LC_9_18_7.C_ON=1'b1;
    defparam un7_spon_cry_15_c_LC_9_18_7.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_15_c_LC_9_18_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_15_c_LC_9_18_7 (
            .in0(_gnd_net_),
            .in1(N__31480),
            .in2(N__52745),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_14),
            .carryout(un7_spon_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_16_c_LC_9_19_0.C_ON=1'b1;
    defparam un7_spon_cry_16_c_LC_9_19_0.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_16_c_LC_9_19_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_16_c_LC_9_19_0 (
            .in0(_gnd_net_),
            .in1(N__52747),
            .in2(N__31393),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(un7_spon_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_17_c_LC_9_19_1.C_ON=1'b1;
    defparam un7_spon_cry_17_c_LC_9_19_1.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_17_c_LC_9_19_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_17_c_LC_9_19_1 (
            .in0(_gnd_net_),
            .in1(N__31285),
            .in2(N__52783),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_16),
            .carryout(un7_spon_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_18_c_LC_9_19_2.C_ON=1'b1;
    defparam un7_spon_cry_18_c_LC_9_19_2.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_18_c_LC_9_19_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_18_c_LC_9_19_2 (
            .in0(_gnd_net_),
            .in1(N__52751),
            .in2(N__31178),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_17),
            .carryout(un7_spon_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_19_c_LC_9_19_3.C_ON=1'b1;
    defparam un7_spon_cry_19_c_LC_9_19_3.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_19_c_LC_9_19_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_19_c_LC_9_19_3 (
            .in0(_gnd_net_),
            .in1(N__33277),
            .in2(N__52784),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_18),
            .carryout(un7_spon_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_20_c_LC_9_19_4.C_ON=1'b1;
    defparam un7_spon_cry_20_c_LC_9_19_4.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_20_c_LC_9_19_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_20_c_LC_9_19_4 (
            .in0(_gnd_net_),
            .in1(N__52755),
            .in2(N__33389),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_19),
            .carryout(un7_spon_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_21_c_LC_9_19_5.C_ON=1'b1;
    defparam un7_spon_cry_21_c_LC_9_19_5.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_21_c_LC_9_19_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_21_c_LC_9_19_5 (
            .in0(_gnd_net_),
            .in1(N__33170),
            .in2(N__52785),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_20),
            .carryout(un7_spon_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_22_c_LC_9_19_6.C_ON=1'b1;
    defparam un7_spon_cry_22_c_LC_9_19_6.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_22_c_LC_9_19_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_22_c_LC_9_19_6 (
            .in0(_gnd_net_),
            .in1(N__52759),
            .in2(N__32047),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_21),
            .carryout(un7_spon_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_23_c_LC_9_19_7.C_ON=1'b1;
    defparam un7_spon_cry_23_c_LC_9_19_7.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_23_c_LC_9_19_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_23_c_LC_9_19_7 (
            .in0(_gnd_net_),
            .in1(N__31934),
            .in2(N__52786),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_22),
            .carryout(un7_spon_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pon_obuf_RNO_LC_9_20_0.C_ON=1'b0;
    defparam pon_obuf_RNO_LC_9_20_0.SEQ_MODE=4'b0000;
    defparam pon_obuf_RNO_LC_9_20_0.LUT_INIT=16'b0000000011101110;
    LogicCell40 pon_obuf_RNO_LC_9_20_0 (
            .in0(N__31059),
            .in1(N__29561),
            .in2(_gnd_net_),
            .in3(N__24017),
            .lcout(pon_obuf_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_10_LC_10_3_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_10_LC_10_3_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_10_LC_10_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_10_LC_10_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23975),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48448),
            .ce(),
            .sr(N__51781));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_15_LC_10_3_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_15_LC_10_3_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_15_LC_10_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_15_LC_10_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24023),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48448),
            .ce(),
            .sr(N__51781));
    defparam \spi_master_inst.spi_data_path_u1.data_in_0_LC_10_4_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_0_LC_10_4_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_0_LC_10_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_0_LC_10_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24782),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48452),
            .ce(N__43901),
            .sr(N__51767));
    defparam \spi_master_inst.spi_data_path_u1.data_in_1_LC_10_4_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_1_LC_10_4_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_1_LC_10_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_1_LC_10_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24776),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48452),
            .ce(N__43901),
            .sr(N__51767));
    defparam \spi_master_inst.spi_data_path_u1.data_in_10_LC_10_4_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_10_LC_10_4_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_10_LC_10_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_10_LC_10_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29498),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48452),
            .ce(N__43901),
            .sr(N__51767));
    defparam \spi_master_inst.spi_data_path_u1.data_in_11_LC_10_4_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_11_LC_10_4_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_11_LC_10_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_11_LC_10_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24770),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48452),
            .ce(N__43901),
            .sr(N__51767));
    defparam \spi_master_inst.spi_data_path_u1.data_in_12_LC_10_4_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_12_LC_10_4_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_12_LC_10_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_12_LC_10_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24764),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48452),
            .ce(N__43901),
            .sr(N__51767));
    defparam \spi_master_inst.spi_data_path_u1.data_in_13_LC_10_4_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_13_LC_10_4_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_13_LC_10_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_13_LC_10_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24758),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48452),
            .ce(N__43901),
            .sr(N__51767));
    defparam \spi_master_inst.spi_data_path_u1.data_in_14_LC_10_4_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_14_LC_10_4_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_14_LC_10_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_14_LC_10_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24752),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48452),
            .ce(N__43901),
            .sr(N__51767));
    defparam \spi_master_inst.spi_data_path_u1.data_in_15_LC_10_4_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_15_LC_10_4_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_15_LC_10_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_15_LC_10_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24746),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48452),
            .ce(N__43901),
            .sr(N__51767));
    defparam sDAC_mem_42_0_LC_10_5_0.C_ON=1'b0;
    defparam sDAC_mem_42_0_LC_10_5_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_0_LC_10_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_42_0_LC_10_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46050),
            .lcout(sDAC_mem_42Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52328),
            .ce(N__24062),
            .sr(N__51754));
    defparam sDAC_mem_42_1_LC_10_5_1.C_ON=1'b0;
    defparam sDAC_mem_42_1_LC_10_5_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_1_LC_10_5_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_42_1_LC_10_5_1 (
            .in0(N__50814),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_42Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52328),
            .ce(N__24062),
            .sr(N__51754));
    defparam sDAC_mem_42_2_LC_10_5_2.C_ON=1'b0;
    defparam sDAC_mem_42_2_LC_10_5_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_2_LC_10_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_42_2_LC_10_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47169),
            .lcout(sDAC_mem_42Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52328),
            .ce(N__24062),
            .sr(N__51754));
    defparam sDAC_mem_42_3_LC_10_5_3.C_ON=1'b0;
    defparam sDAC_mem_42_3_LC_10_5_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_3_LC_10_5_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_42_3_LC_10_5_3 (
            .in0(N__46598),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_42Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52328),
            .ce(N__24062),
            .sr(N__51754));
    defparam sDAC_mem_42_4_LC_10_5_4.C_ON=1'b0;
    defparam sDAC_mem_42_4_LC_10_5_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_4_LC_10_5_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_42_4_LC_10_5_4 (
            .in0(N__45296),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_42Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52328),
            .ce(N__24062),
            .sr(N__51754));
    defparam sDAC_mem_42_5_LC_10_5_5.C_ON=1'b0;
    defparam sDAC_mem_42_5_LC_10_5_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_5_LC_10_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_42_5_LC_10_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44951),
            .lcout(sDAC_mem_42Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52328),
            .ce(N__24062),
            .sr(N__51754));
    defparam sDAC_mem_42_6_LC_10_5_6.C_ON=1'b0;
    defparam sDAC_mem_42_6_LC_10_5_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_6_LC_10_5_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_42_6_LC_10_5_6 (
            .in0(N__50225),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_42Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52328),
            .ce(N__24062),
            .sr(N__51754));
    defparam sDAC_mem_42_7_LC_10_5_7.C_ON=1'b0;
    defparam sDAC_mem_42_7_LC_10_5_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_7_LC_10_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_42_7_LC_10_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49727),
            .lcout(sDAC_mem_42Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52328),
            .ce(N__24062),
            .sr(N__51754));
    defparam sDAC_mem_14_0_LC_10_6_0.C_ON=1'b0;
    defparam sDAC_mem_14_0_LC_10_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_0_LC_10_6_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_14_0_LC_10_6_0 (
            .in0(N__46210),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_14Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52317),
            .ce(N__24092),
            .sr(N__51741));
    defparam sDAC_mem_14_1_LC_10_6_1.C_ON=1'b0;
    defparam sDAC_mem_14_1_LC_10_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_1_LC_10_6_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_14_1_LC_10_6_1 (
            .in0(N__50896),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_14Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52317),
            .ce(N__24092),
            .sr(N__51741));
    defparam sDAC_mem_14_2_LC_10_6_2.C_ON=1'b0;
    defparam sDAC_mem_14_2_LC_10_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_2_LC_10_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_2_LC_10_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47275),
            .lcout(sDAC_mem_14Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52317),
            .ce(N__24092),
            .sr(N__51741));
    defparam sDAC_mem_14_3_LC_10_6_3.C_ON=1'b0;
    defparam sDAC_mem_14_3_LC_10_6_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_3_LC_10_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_3_LC_10_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46708),
            .lcout(sDAC_mem_14Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52317),
            .ce(N__24092),
            .sr(N__51741));
    defparam sDAC_mem_14_4_LC_10_6_4.C_ON=1'b0;
    defparam sDAC_mem_14_4_LC_10_6_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_4_LC_10_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_4_LC_10_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45410),
            .lcout(sDAC_mem_14Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52317),
            .ce(N__24092),
            .sr(N__51741));
    defparam sDAC_mem_14_5_LC_10_6_5.C_ON=1'b0;
    defparam sDAC_mem_14_5_LC_10_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_5_LC_10_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_5_LC_10_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44928),
            .lcout(sDAC_mem_14Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52317),
            .ce(N__24092),
            .sr(N__51741));
    defparam sDAC_mem_14_6_LC_10_6_6.C_ON=1'b0;
    defparam sDAC_mem_14_6_LC_10_6_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_6_LC_10_6_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_14_6_LC_10_6_6 (
            .in0(N__50306),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_14Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52317),
            .ce(N__24092),
            .sr(N__51741));
    defparam sDAC_mem_14_7_LC_10_6_7.C_ON=1'b0;
    defparam sDAC_mem_14_7_LC_10_6_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_7_LC_10_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_7_LC_10_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49832),
            .lcout(sDAC_mem_14Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52317),
            .ce(N__24092),
            .sr(N__51741));
    defparam sEEPeriod_10_LC_10_7_0.C_ON=1'b0;
    defparam sEEPeriod_10_LC_10_7_0.SEQ_MODE=4'b1011;
    defparam sEEPeriod_10_LC_10_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_10_LC_10_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47393),
            .lcout(sEEPeriodZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52306),
            .ce(N__24077),
            .sr(N__51727));
    defparam sEEPeriod_11_LC_10_7_1.C_ON=1'b0;
    defparam sEEPeriod_11_LC_10_7_1.SEQ_MODE=4'b1010;
    defparam sEEPeriod_11_LC_10_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_11_LC_10_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46829),
            .lcout(sEEPeriodZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52306),
            .ce(N__24077),
            .sr(N__51727));
    defparam sEEPeriod_12_LC_10_7_2.C_ON=1'b0;
    defparam sEEPeriod_12_LC_10_7_2.SEQ_MODE=4'b1010;
    defparam sEEPeriod_12_LC_10_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_12_LC_10_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45411),
            .lcout(sEEPeriodZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52306),
            .ce(N__24077),
            .sr(N__51727));
    defparam sEEPeriod_13_LC_10_7_3.C_ON=1'b0;
    defparam sEEPeriod_13_LC_10_7_3.SEQ_MODE=4'b1010;
    defparam sEEPeriod_13_LC_10_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_13_LC_10_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44923),
            .lcout(sEEPeriodZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52306),
            .ce(N__24077),
            .sr(N__51727));
    defparam sEEPeriod_14_LC_10_7_4.C_ON=1'b0;
    defparam sEEPeriod_14_LC_10_7_4.SEQ_MODE=4'b1010;
    defparam sEEPeriod_14_LC_10_7_4.LUT_INIT=16'b1100110011001100;
    LogicCell40 sEEPeriod_14_LC_10_7_4 (
            .in0(_gnd_net_),
            .in1(N__50307),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52306),
            .ce(N__24077),
            .sr(N__51727));
    defparam sEEPeriod_15_LC_10_7_5.C_ON=1'b0;
    defparam sEEPeriod_15_LC_10_7_5.SEQ_MODE=4'b1011;
    defparam sEEPeriod_15_LC_10_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_15_LC_10_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49789),
            .lcout(sEEPeriodZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52306),
            .ce(N__24077),
            .sr(N__51727));
    defparam sEEPeriod_8_LC_10_7_6.C_ON=1'b0;
    defparam sEEPeriod_8_LC_10_7_6.SEQ_MODE=4'b1010;
    defparam sEEPeriod_8_LC_10_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_8_LC_10_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46054),
            .lcout(sEEPeriodZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52306),
            .ce(N__24077),
            .sr(N__51727));
    defparam sEEPeriod_9_LC_10_7_7.C_ON=1'b0;
    defparam sEEPeriod_9_LC_10_7_7.SEQ_MODE=4'b1011;
    defparam sEEPeriod_9_LC_10_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_9_LC_10_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50898),
            .lcout(sEEPeriodZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52306),
            .ce(N__24077),
            .sr(N__51727));
    defparam sEEPeriod_16_LC_10_8_0.C_ON=1'b0;
    defparam sEEPeriod_16_LC_10_8_0.SEQ_MODE=4'b1011;
    defparam sEEPeriod_16_LC_10_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_16_LC_10_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46391),
            .lcout(sEEPeriodZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52294),
            .ce(N__24107),
            .sr(N__51715));
    defparam sEEPeriod_17_LC_10_8_1.C_ON=1'b0;
    defparam sEEPeriod_17_LC_10_8_1.SEQ_MODE=4'b1010;
    defparam sEEPeriod_17_LC_10_8_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPeriod_17_LC_10_8_1 (
            .in0(N__50897),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52294),
            .ce(N__24107),
            .sr(N__51715));
    defparam sEEPeriod_18_LC_10_8_2.C_ON=1'b0;
    defparam sEEPeriod_18_LC_10_8_2.SEQ_MODE=4'b1010;
    defparam sEEPeriod_18_LC_10_8_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPeriod_18_LC_10_8_2 (
            .in0(N__47394),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52294),
            .ce(N__24107),
            .sr(N__51715));
    defparam sEEPeriod_19_LC_10_8_3.C_ON=1'b0;
    defparam sEEPeriod_19_LC_10_8_3.SEQ_MODE=4'b1010;
    defparam sEEPeriod_19_LC_10_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_19_LC_10_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46769),
            .lcout(sEEPeriodZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52294),
            .ce(N__24107),
            .sr(N__51715));
    defparam sEEPeriod_20_LC_10_8_4.C_ON=1'b0;
    defparam sEEPeriod_20_LC_10_8_4.SEQ_MODE=4'b1010;
    defparam sEEPeriod_20_LC_10_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_20_LC_10_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45412),
            .lcout(sEEPeriodZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52294),
            .ce(N__24107),
            .sr(N__51715));
    defparam sEEPeriod_21_LC_10_8_5.C_ON=1'b0;
    defparam sEEPeriod_21_LC_10_8_5.SEQ_MODE=4'b1010;
    defparam sEEPeriod_21_LC_10_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_21_LC_10_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44929),
            .lcout(sEEPeriodZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52294),
            .ce(N__24107),
            .sr(N__51715));
    defparam sEEPeriod_22_LC_10_8_6.C_ON=1'b0;
    defparam sEEPeriod_22_LC_10_8_6.SEQ_MODE=4'b1010;
    defparam sEEPeriod_22_LC_10_8_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPeriod_22_LC_10_8_6 (
            .in0(N__50308),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52294),
            .ce(N__24107),
            .sr(N__51715));
    defparam sEEPeriod_23_LC_10_8_7.C_ON=1'b0;
    defparam sEEPeriod_23_LC_10_8_7.SEQ_MODE=4'b1010;
    defparam sEEPeriod_23_LC_10_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_23_LC_10_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49833),
            .lcout(sEEPeriodZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52294),
            .ce(N__24107),
            .sr(N__51715));
    defparam sDAC_mem_15_0_LC_10_9_0.C_ON=1'b0;
    defparam sDAC_mem_15_0_LC_10_9_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_0_LC_10_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_0_LC_10_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46375),
            .lcout(sDAC_mem_15Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52283),
            .ce(N__24113),
            .sr(N__51704));
    defparam sDAC_mem_15_1_LC_10_9_1.C_ON=1'b0;
    defparam sDAC_mem_15_1_LC_10_9_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_1_LC_10_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_1_LC_10_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50899),
            .lcout(sDAC_mem_15Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52283),
            .ce(N__24113),
            .sr(N__51704));
    defparam sDAC_mem_15_2_LC_10_9_2.C_ON=1'b0;
    defparam sDAC_mem_15_2_LC_10_9_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_2_LC_10_9_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_15_2_LC_10_9_2 (
            .in0(N__47395),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_15Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52283),
            .ce(N__24113),
            .sr(N__51704));
    defparam sDAC_mem_15_3_LC_10_9_3.C_ON=1'b0;
    defparam sDAC_mem_15_3_LC_10_9_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_3_LC_10_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_3_LC_10_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46852),
            .lcout(sDAC_mem_15Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52283),
            .ce(N__24113),
            .sr(N__51704));
    defparam sDAC_mem_15_4_LC_10_9_4.C_ON=1'b0;
    defparam sDAC_mem_15_4_LC_10_9_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_4_LC_10_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_4_LC_10_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45413),
            .lcout(sDAC_mem_15Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52283),
            .ce(N__24113),
            .sr(N__51704));
    defparam sDAC_mem_15_5_LC_10_9_5.C_ON=1'b0;
    defparam sDAC_mem_15_5_LC_10_9_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_5_LC_10_9_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_15_5_LC_10_9_5 (
            .in0(N__44924),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_15Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52283),
            .ce(N__24113),
            .sr(N__51704));
    defparam sDAC_mem_15_6_LC_10_9_6.C_ON=1'b0;
    defparam sDAC_mem_15_6_LC_10_9_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_6_LC_10_9_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_15_6_LC_10_9_6 (
            .in0(N__50309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_15Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52283),
            .ce(N__24113),
            .sr(N__51704));
    defparam sDAC_mem_15_7_LC_10_9_7.C_ON=1'b0;
    defparam sDAC_mem_15_7_LC_10_9_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_7_LC_10_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_7_LC_10_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49834),
            .lcout(sDAC_mem_15Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52283),
            .ce(N__24113),
            .sr(N__51704));
    defparam sDAC_mem_18_0_LC_10_10_0.C_ON=1'b0;
    defparam sDAC_mem_18_0_LC_10_10_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_0_LC_10_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_0_LC_10_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46209),
            .lcout(sDAC_mem_18Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52272),
            .ce(N__28540),
            .sr(N__51697));
    defparam sDAC_mem_18_1_LC_10_10_1.C_ON=1'b0;
    defparam sDAC_mem_18_1_LC_10_10_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_1_LC_10_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_1_LC_10_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50983),
            .lcout(sDAC_mem_18Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52272),
            .ce(N__28540),
            .sr(N__51697));
    defparam sDAC_mem_18_2_LC_10_10_2.C_ON=1'b0;
    defparam sDAC_mem_18_2_LC_10_10_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_2_LC_10_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_2_LC_10_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47461),
            .lcout(sDAC_mem_18Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52272),
            .ce(N__28540),
            .sr(N__51697));
    defparam sDAC_mem_18_7_LC_10_10_3.C_ON=1'b0;
    defparam sDAC_mem_18_7_LC_10_10_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_7_LC_10_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_7_LC_10_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49939),
            .lcout(sDAC_mem_18Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52272),
            .ce(N__28540),
            .sr(N__51697));
    defparam sCounter_RNI0D9U_10_LC_10_11_0.C_ON=1'b0;
    defparam sCounter_RNI0D9U_10_LC_10_11_0.SEQ_MODE=4'b0000;
    defparam sCounter_RNI0D9U_10_LC_10_11_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNI0D9U_10_LC_10_11_0 (
            .in0(N__30534),
            .in1(N__33039),
            .in2(N__30446),
            .in3(N__30314),
            .lcout(op_gt_op_gt_un13_striginternallto23_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIQB5R1_1_LC_10_11_1.C_ON=1'b0;
    defparam sCounter_RNIQB5R1_1_LC_10_11_1.SEQ_MODE=4'b0000;
    defparam sCounter_RNIQB5R1_1_LC_10_11_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNIQB5R1_1_LC_10_11_1 (
            .in0(N__30081),
            .in1(N__29841),
            .in2(N__24155),
            .in3(N__29970),
            .lcout(),
            .ltout(op_gt_op_gt_un13_striginternallto23_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIVUR25_16_LC_10_11_2.C_ON=1'b0;
    defparam sCounter_RNIVUR25_16_LC_10_11_2.SEQ_MODE=4'b0000;
    defparam sCounter_RNIVUR25_16_LC_10_11_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 sCounter_RNIVUR25_16_LC_10_11_2 (
            .in0(N__24119),
            .in1(N__24197),
            .in2(N__24185),
            .in3(N__24167),
            .lcout(op_gt_op_gt_un13_striginternal_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNI2RIT_8_LC_10_11_3.C_ON=1'b0;
    defparam sCounter_RNI2RIT_8_LC_10_11_3.SEQ_MODE=4'b0000;
    defparam sCounter_RNI2RIT_8_LC_10_11_3.LUT_INIT=16'b1111111111101110;
    LogicCell40 sCounter_RNI2RIT_8_LC_10_11_3 (
            .in0(N__30204),
            .in1(N__30422),
            .in2(_gnd_net_),
            .in3(N__30533),
            .lcout(un1_reset_rpi_inv_2_0_o2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNI9MMP_12_LC_10_11_4.C_ON=1'b0;
    defparam sCounter_RNI9MMP_12_LC_10_11_4.SEQ_MODE=4'b0000;
    defparam sCounter_RNI9MMP_12_LC_10_11_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNI9MMP_12_LC_10_11_4 (
            .in0(N__31630),
            .in1(N__31717),
            .in2(N__31467),
            .in3(N__30205),
            .lcout(g0_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIES4L_16_LC_10_11_5.C_ON=1'b0;
    defparam sCounter_RNIES4L_16_LC_10_11_5.SEQ_MODE=4'b0000;
    defparam sCounter_RNIES4L_16_LC_10_11_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNIES4L_16_LC_10_11_5 (
            .in0(N__31336),
            .in1(N__33223),
            .in2(N__31268),
            .in3(N__31123),
            .lcout(un21_trig_prev_21_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIU3NJ_1_LC_10_11_6.C_ON=1'b0;
    defparam sCounter_RNIU3NJ_1_LC_10_11_6.SEQ_MODE=4'b0000;
    defparam sCounter_RNIU3NJ_1_LC_10_11_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 sCounter_RNIU3NJ_1_LC_10_11_6 (
            .in0(_gnd_net_),
            .in1(N__30080),
            .in2(_gnd_net_),
            .in3(N__30634),
            .lcout(g0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNI3SIT_5_LC_10_12_0.C_ON=1'b0;
    defparam sCounter_RNI3SIT_5_LC_10_12_0.SEQ_MODE=4'b0000;
    defparam sCounter_RNI3SIT_5_LC_10_12_0.LUT_INIT=16'b1111111111101110;
    LogicCell40 sCounter_RNI3SIT_5_LC_10_12_0 (
            .in0(N__30675),
            .in1(N__30773),
            .in2(_gnd_net_),
            .in3(N__30880),
            .lcout(N_99),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNITA9T1_4_LC_10_12_1.C_ON=1'b0;
    defparam sCounter_RNITA9T1_4_LC_10_12_1.SEQ_MODE=4'b0000;
    defparam sCounter_RNITA9T1_4_LC_10_12_1.LUT_INIT=16'b0100000001000000;
    LogicCell40 sCounter_RNITA9T1_4_LC_10_12_1 (
            .in0(N__31000),
            .in1(N__24143),
            .in2(N__24137),
            .in3(_gnd_net_),
            .lcout(op_gt_op_gt_un13_striginternallto23_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNIJFMR_1_LC_10_12_3 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNIJFMR_1_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNIJFMR_1_LC_10_12_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNIJFMR_1_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__25489),
            .in2(_gnd_net_),
            .in3(N__25255),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNILEDN1_7_LC_10_12_4 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNILEDN1_7_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNILEDN1_7_LC_10_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNILEDN1_7_LC_10_12_4  (
            .in0(N__25399),
            .in1(N__25474),
            .in2(N__25436),
            .in3(N__25417),
            .lcout(),
            .ltout(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNISEQE3_0_LC_10_12_5 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNISEQE3_0_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNISEQE3_0_LC_10_12_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNISEQE3_0_LC_10_12_5  (
            .in0(N__25460),
            .in1(N__25270),
            .in2(N__24560),
            .in3(N__24557),
            .lcout(\spi_master_inst.sclk_gen_u0.N_158_7 ),
            .ltout(\spi_master_inst.sclk_gen_u0.N_158_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNO_0_LC_10_12_6 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNO_0_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNO_0_LC_10_12_6 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNO_0_LC_10_12_6  (
            .in0(N__24520),
            .in1(N__24455),
            .in2(N__24392),
            .in3(N__24388),
            .lcout(\spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIS7E71_2_LC_10_12_7.C_ON=1'b0;
    defparam sCounter_RNIS7E71_2_LC_10_12_7.SEQ_MODE=4'b0000;
    defparam sCounter_RNIS7E71_2_LC_10_12_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNIS7E71_2_LC_10_12_7 (
            .in0(N__30879),
            .in1(N__29851),
            .in2(N__30785),
            .in3(N__29983),
            .lcout(g2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNILK4P2_3_LC_10_13_1 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNILK4P2_3_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNILK4P2_3_LC_10_13_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_RNILK4P2_3_LC_10_13_1  (
            .in0(N__24308),
            .in1(N__24290),
            .in2(_gnd_net_),
            .in3(N__24272),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_i6 ),
            .ltout(\spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3_3_LC_10_13_2 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3_3_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3_3_LC_10_13_2 .LUT_INIT=16'b0000010000000111;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3_3_LC_10_13_2  (
            .in0(N__47892),
            .in1(N__48006),
            .in2(N__24224),
            .in3(N__47956),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNICH5T1_5_LC_10_13_3 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNICH5T1_5_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNICH5T1_5_LC_10_13_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_RNICH5T1_5_LC_10_13_3  (
            .in0(N__42773),
            .in1(N__42683),
            .in2(N__42740),
            .in3(N__38657),
            .lcout(\spi_slave_inst.un23_i_ssn_3 ),
            .ltout(\spi_slave_inst.un23_i_ssn_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI5DOR2_3_LC_10_13_4 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI5DOR2_3_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI5DOR2_3_LC_10_13_4 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_RNI5DOR2_3_LC_10_13_4  (
            .in0(N__48304),
            .in1(_gnd_net_),
            .in2(N__24200),
            .in3(N__48329),
            .lcout(\spi_slave_inst.un23_i_ssn ),
            .ltout(\spi_slave_inst.un23_i_ssn_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI4ODL3_3_LC_10_13_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI4ODL3_3_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI4ODL3_3_LC_10_13_5 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_RNI4ODL3_3_LC_10_13_5  (
            .in0(N__47957),
            .in1(N__48007),
            .in2(N__24578),
            .in3(N__47893),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNI4K6L_23_LC_10_13_6.C_ON=1'b0;
    defparam sCounter_RNI4K6L_23_LC_10_13_6.SEQ_MODE=4'b0000;
    defparam sCounter_RNI4K6L_23_LC_10_13_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNI4K6L_23_LC_10_13_6 (
            .in0(N__31376),
            .in1(N__31239),
            .in2(N__31905),
            .in3(N__31990),
            .lcout(g0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNI5I9U_16_LC_10_13_7.C_ON=1'b0;
    defparam sCounter_RNI5I9U_16_LC_10_13_7.SEQ_MODE=4'b0000;
    defparam sCounter_RNI5I9U_16_LC_10_13_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNI5I9U_16_LC_10_13_7 (
            .in0(N__30769),
            .in1(N__31377),
            .in2(N__31267),
            .in3(N__30999),
            .lcout(g0_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_31_0_LC_10_14_0.C_ON=1'b0;
    defparam sDAC_mem_31_0_LC_10_14_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_0_LC_10_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_0_LC_10_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46338),
            .lcout(sDAC_mem_31Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52295),
            .ce(N__24593),
            .sr(N__51667));
    defparam sDAC_mem_31_1_LC_10_14_1.C_ON=1'b0;
    defparam sDAC_mem_31_1_LC_10_14_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_1_LC_10_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_1_LC_10_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50878),
            .lcout(sDAC_mem_31Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52295),
            .ce(N__24593),
            .sr(N__51667));
    defparam sDAC_mem_31_2_LC_10_14_2.C_ON=1'b0;
    defparam sDAC_mem_31_2_LC_10_14_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_2_LC_10_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_2_LC_10_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47499),
            .lcout(sDAC_mem_31Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52295),
            .ce(N__24593),
            .sr(N__51667));
    defparam sDAC_mem_31_3_LC_10_14_3.C_ON=1'b0;
    defparam sDAC_mem_31_3_LC_10_14_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_3_LC_10_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_3_LC_10_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46913),
            .lcout(sDAC_mem_31Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52295),
            .ce(N__24593),
            .sr(N__51667));
    defparam sDAC_mem_31_4_LC_10_14_4.C_ON=1'b0;
    defparam sDAC_mem_31_4_LC_10_14_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_4_LC_10_14_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_31_4_LC_10_14_4 (
            .in0(N__45579),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_31Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52295),
            .ce(N__24593),
            .sr(N__51667));
    defparam sDAC_mem_31_5_LC_10_14_5.C_ON=1'b0;
    defparam sDAC_mem_31_5_LC_10_14_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_5_LC_10_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_5_LC_10_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45090),
            .lcout(sDAC_mem_31Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52295),
            .ce(N__24593),
            .sr(N__51667));
    defparam sDAC_mem_31_6_LC_10_14_6.C_ON=1'b0;
    defparam sDAC_mem_31_6_LC_10_14_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_6_LC_10_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_6_LC_10_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50529),
            .lcout(sDAC_mem_31Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52295),
            .ce(N__24593),
            .sr(N__51667));
    defparam sDAC_mem_31_7_LC_10_14_7.C_ON=1'b0;
    defparam sDAC_mem_31_7_LC_10_14_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_7_LC_10_14_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_31_7_LC_10_14_7 (
            .in0(N__50028),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_31Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52295),
            .ce(N__24593),
            .sr(N__51667));
    defparam sDAC_mem_24_0_LC_10_15_0.C_ON=1'b0;
    defparam sDAC_mem_24_0_LC_10_15_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_0_LC_10_15_0.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_24_0_LC_10_15_0 (
            .in0(_gnd_net_),
            .in1(N__46322),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_24Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52307),
            .ce(N__27745),
            .sr(N__51661));
    defparam sDAC_mem_24_2_LC_10_15_1.C_ON=1'b0;
    defparam sDAC_mem_24_2_LC_10_15_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_2_LC_10_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_2_LC_10_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47500),
            .lcout(sDAC_mem_24Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52307),
            .ce(N__27745),
            .sr(N__51661));
    defparam sDAC_mem_24_3_LC_10_15_2.C_ON=1'b0;
    defparam sDAC_mem_24_3_LC_10_15_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_3_LC_10_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_3_LC_10_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46847),
            .lcout(sDAC_mem_24Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52307),
            .ce(N__27745),
            .sr(N__51661));
    defparam sDAC_mem_24_5_LC_10_15_3.C_ON=1'b0;
    defparam sDAC_mem_24_5_LC_10_15_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_5_LC_10_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_5_LC_10_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45094),
            .lcout(sDAC_mem_24Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52307),
            .ce(N__27745),
            .sr(N__51661));
    defparam sDAC_mem_24_6_LC_10_15_4.C_ON=1'b0;
    defparam sDAC_mem_24_6_LC_10_15_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_6_LC_10_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_6_LC_10_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50391),
            .lcout(sDAC_mem_24Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52307),
            .ce(N__27745),
            .sr(N__51661));
    defparam sDAC_mem_24_7_LC_10_15_5.C_ON=1'b0;
    defparam sDAC_mem_24_7_LC_10_15_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_7_LC_10_15_5.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_24_7_LC_10_15_5 (
            .in0(_gnd_net_),
            .in1(N__50029),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_24Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52307),
            .ce(N__27745),
            .sr(N__51661));
    defparam sDAC_mem_28_0_LC_10_16_0.C_ON=1'b0;
    defparam sDAC_mem_28_0_LC_10_16_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_0_LC_10_16_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_28_0_LC_10_16_0 (
            .in0(N__46321),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_28Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52318),
            .ce(N__37789),
            .sr(N__51655));
    defparam sDAC_mem_28_1_LC_10_16_1.C_ON=1'b0;
    defparam sDAC_mem_28_1_LC_10_16_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_1_LC_10_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_1_LC_10_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51037),
            .lcout(sDAC_mem_28Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52318),
            .ce(N__37789),
            .sr(N__51655));
    defparam sDAC_mem_28_3_LC_10_16_2.C_ON=1'b0;
    defparam sDAC_mem_28_3_LC_10_16_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_3_LC_10_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_3_LC_10_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46762),
            .lcout(sDAC_mem_28Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52318),
            .ce(N__37789),
            .sr(N__51655));
    defparam sDAC_mem_28_4_LC_10_16_3.C_ON=1'b0;
    defparam sDAC_mem_28_4_LC_10_16_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_4_LC_10_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_4_LC_10_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45580),
            .lcout(sDAC_mem_28Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52318),
            .ce(N__37789),
            .sr(N__51655));
    defparam sEEDelayACQ_0_LC_10_17_0.C_ON=1'b0;
    defparam sEEDelayACQ_0_LC_10_17_0.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_0_LC_10_17_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEDelayACQ_0_LC_10_17_0 (
            .in0(N__46323),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52329),
            .ce(N__24605),
            .sr(N__51652));
    defparam sEEDelayACQ_1_LC_10_17_1.C_ON=1'b0;
    defparam sEEDelayACQ_1_LC_10_17_1.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_1_LC_10_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_1_LC_10_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51038),
            .lcout(sEEDelayACQZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52329),
            .ce(N__24605),
            .sr(N__51652));
    defparam sEEDelayACQ_2_LC_10_17_2.C_ON=1'b0;
    defparam sEEDelayACQ_2_LC_10_17_2.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_2_LC_10_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_2_LC_10_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47502),
            .lcout(sEEDelayACQZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52329),
            .ce(N__24605),
            .sr(N__51652));
    defparam sEEDelayACQ_3_LC_10_17_3.C_ON=1'b0;
    defparam sEEDelayACQ_3_LC_10_17_3.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_3_LC_10_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_3_LC_10_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46851),
            .lcout(sEEDelayACQZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52329),
            .ce(N__24605),
            .sr(N__51652));
    defparam sEEDelayACQ_4_LC_10_17_4.C_ON=1'b0;
    defparam sEEDelayACQ_4_LC_10_17_4.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_4_LC_10_17_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEDelayACQ_4_LC_10_17_4 (
            .in0(N__45581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52329),
            .ce(N__24605),
            .sr(N__51652));
    defparam sEEDelayACQ_5_LC_10_17_5.C_ON=1'b0;
    defparam sEEDelayACQ_5_LC_10_17_5.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_5_LC_10_17_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEDelayACQ_5_LC_10_17_5 (
            .in0(N__45095),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52329),
            .ce(N__24605),
            .sr(N__51652));
    defparam sEEDelayACQ_6_LC_10_17_6.C_ON=1'b0;
    defparam sEEDelayACQ_6_LC_10_17_6.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_6_LC_10_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_6_LC_10_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50392),
            .lcout(sEEDelayACQZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52329),
            .ce(N__24605),
            .sr(N__51652));
    defparam sEEDelayACQ_7_LC_10_17_7.C_ON=1'b0;
    defparam sEEDelayACQ_7_LC_10_17_7.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_7_LC_10_17_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEDelayACQ_7_LC_10_17_7 (
            .in0(N__50031),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52329),
            .ce(N__24605),
            .sr(N__51652));
    defparam sEEDelayACQ_10_LC_10_18_0.C_ON=1'b0;
    defparam sEEDelayACQ_10_LC_10_18_0.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_10_LC_10_18_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEDelayACQ_10_LC_10_18_0 (
            .in0(N__47512),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52338),
            .ce(N__24740),
            .sr(N__51649));
    defparam sEEDelayACQ_11_LC_10_18_1.C_ON=1'b0;
    defparam sEEDelayACQ_11_LC_10_18_1.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_11_LC_10_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_11_LC_10_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46924),
            .lcout(sEEDelayACQZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52338),
            .ce(N__24740),
            .sr(N__51649));
    defparam sEEDelayACQ_12_LC_10_18_2.C_ON=1'b0;
    defparam sEEDelayACQ_12_LC_10_18_2.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_12_LC_10_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_12_LC_10_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45604),
            .lcout(sEEDelayACQZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52338),
            .ce(N__24740),
            .sr(N__51649));
    defparam sEEDelayACQ_13_LC_10_18_3.C_ON=1'b0;
    defparam sEEDelayACQ_13_LC_10_18_3.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_13_LC_10_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_13_LC_10_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45116),
            .lcout(sEEDelayACQZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52338),
            .ce(N__24740),
            .sr(N__51649));
    defparam sEEDelayACQ_14_LC_10_18_4.C_ON=1'b0;
    defparam sEEDelayACQ_14_LC_10_18_4.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_14_LC_10_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_14_LC_10_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50467),
            .lcout(sEEDelayACQZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52338),
            .ce(N__24740),
            .sr(N__51649));
    defparam sEEDelayACQ_15_LC_10_18_5.C_ON=1'b0;
    defparam sEEDelayACQ_15_LC_10_18_5.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_15_LC_10_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_15_LC_10_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50051),
            .lcout(sEEDelayACQZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52338),
            .ce(N__24740),
            .sr(N__51649));
    defparam sEEDelayACQ_8_LC_10_18_6.C_ON=1'b0;
    defparam sEEDelayACQ_8_LC_10_18_6.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_8_LC_10_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_8_LC_10_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46331),
            .lcout(sEEDelayACQZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52338),
            .ce(N__24740),
            .sr(N__51649));
    defparam sEEDelayACQ_9_LC_10_18_7.C_ON=1'b0;
    defparam sEEDelayACQ_9_LC_10_18_7.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_9_LC_10_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_9_LC_10_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51030),
            .lcout(sEEDelayACQZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52338),
            .ce(N__24740),
            .sr(N__51649));
    defparam reset_rpi_ibuf_RNIIUT3_LC_10_19_1.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNIIUT3_LC_10_19_1.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNIIUT3_LC_10_19_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 reset_rpi_ibuf_RNIIUT3_LC_10_19_1 (
            .in0(N__49246),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(LED3_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4Q_15_LC_11_3_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4Q_15_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4Q_15_LC_11_3_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4Q_15_LC_11_3_7  (
            .in0(N__24710),
            .in1(N__25754),
            .in2(_gnd_net_),
            .in3(N__24704),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_0_LC_11_4_0.C_ON=1'b0;
    defparam sDAC_data_0_LC_11_4_0.SEQ_MODE=4'b1010;
    defparam sDAC_data_0_LC_11_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_0_LC_11_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48449),
            .ce(N__43958),
            .sr(N__51755));
    defparam sDAC_data_1_LC_11_4_1.C_ON=1'b0;
    defparam sDAC_data_1_LC_11_4_1.SEQ_MODE=4'b1010;
    defparam sDAC_data_1_LC_11_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_1_LC_11_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48449),
            .ce(N__43958),
            .sr(N__51755));
    defparam sDAC_data_11_LC_11_4_2.C_ON=1'b0;
    defparam sDAC_data_11_LC_11_4_2.SEQ_MODE=4'b1010;
    defparam sDAC_data_11_LC_11_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_11_LC_11_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48449),
            .ce(N__43958),
            .sr(N__51755));
    defparam sDAC_data_12_LC_11_4_3.C_ON=1'b0;
    defparam sDAC_data_12_LC_11_4_3.SEQ_MODE=4'b1010;
    defparam sDAC_data_12_LC_11_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_12_LC_11_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52649),
            .lcout(sDAC_dataZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48449),
            .ce(N__43958),
            .sr(N__51755));
    defparam sDAC_data_13_LC_11_4_4.C_ON=1'b0;
    defparam sDAC_data_13_LC_11_4_4.SEQ_MODE=4'b1010;
    defparam sDAC_data_13_LC_11_4_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_data_13_LC_11_4_4 (
            .in0(N__52650),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_dataZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48449),
            .ce(N__43958),
            .sr(N__51755));
    defparam sDAC_data_14_LC_11_4_5.C_ON=1'b0;
    defparam sDAC_data_14_LC_11_4_5.SEQ_MODE=4'b1010;
    defparam sDAC_data_14_LC_11_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_14_LC_11_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48449),
            .ce(N__43958),
            .sr(N__51755));
    defparam sDAC_data_15_LC_11_4_6.C_ON=1'b0;
    defparam sDAC_data_15_LC_11_4_6.SEQ_MODE=4'b1010;
    defparam sDAC_data_15_LC_11_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_15_LC_11_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48449),
            .ce(N__43958),
            .sr(N__51755));
    defparam sEEPeriod_0_LC_11_5_0.C_ON=1'b0;
    defparam sEEPeriod_0_LC_11_5_0.SEQ_MODE=4'b1010;
    defparam sEEPeriod_0_LC_11_5_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPeriod_0_LC_11_5_0 (
            .in0(N__46043),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52319),
            .ce(N__24836),
            .sr(N__51742));
    defparam sEEPeriod_1_LC_11_5_1.C_ON=1'b0;
    defparam sEEPeriod_1_LC_11_5_1.SEQ_MODE=4'b1010;
    defparam sEEPeriod_1_LC_11_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_1_LC_11_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50892),
            .lcout(sEEPeriodZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52319),
            .ce(N__24836),
            .sr(N__51742));
    defparam sEEPeriod_2_LC_11_5_2.C_ON=1'b0;
    defparam sEEPeriod_2_LC_11_5_2.SEQ_MODE=4'b1010;
    defparam sEEPeriod_2_LC_11_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_2_LC_11_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47170),
            .lcout(sEEPeriodZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52319),
            .ce(N__24836),
            .sr(N__51742));
    defparam sEEPeriod_3_LC_11_5_3.C_ON=1'b0;
    defparam sEEPeriod_3_LC_11_5_3.SEQ_MODE=4'b1010;
    defparam sEEPeriod_3_LC_11_5_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPeriod_3_LC_11_5_3 (
            .in0(N__46599),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52319),
            .ce(N__24836),
            .sr(N__51742));
    defparam sEEPeriod_4_LC_11_5_4.C_ON=1'b0;
    defparam sEEPeriod_4_LC_11_5_4.SEQ_MODE=4'b1010;
    defparam sEEPeriod_4_LC_11_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_4_LC_11_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45297),
            .lcout(sEEPeriodZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52319),
            .ce(N__24836),
            .sr(N__51742));
    defparam sEEPeriod_5_LC_11_5_5.C_ON=1'b0;
    defparam sEEPeriod_5_LC_11_5_5.SEQ_MODE=4'b1011;
    defparam sEEPeriod_5_LC_11_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_5_LC_11_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44763),
            .lcout(sEEPeriodZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52319),
            .ce(N__24836),
            .sr(N__51742));
    defparam sEEPeriod_6_LC_11_5_6.C_ON=1'b0;
    defparam sEEPeriod_6_LC_11_5_6.SEQ_MODE=4'b1010;
    defparam sEEPeriod_6_LC_11_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_6_LC_11_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50317),
            .lcout(sEEPeriodZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52319),
            .ce(N__24836),
            .sr(N__51742));
    defparam sEEPeriod_7_LC_11_5_7.C_ON=1'b0;
    defparam sEEPeriod_7_LC_11_5_7.SEQ_MODE=4'b1011;
    defparam sEEPeriod_7_LC_11_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_7_LC_11_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49831),
            .lcout(sEEPeriodZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52319),
            .ce(N__24836),
            .sr(N__51742));
    defparam un4_speriod_cry_0_c_inv_LC_11_6_0.C_ON=1'b1;
    defparam un4_speriod_cry_0_c_inv_LC_11_6_0.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_0_c_inv_LC_11_6_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_0_c_inv_LC_11_6_0 (
            .in0(_gnd_net_),
            .in1(N__24818),
            .in2(N__30237),
            .in3(N__24824),
            .lcout(sEEPeriod_i_0),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(un4_speriod_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_1_c_inv_LC_11_6_1.C_ON=1'b1;
    defparam un4_speriod_cry_1_c_inv_LC_11_6_1.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_1_c_inv_LC_11_6_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_1_c_inv_LC_11_6_1 (
            .in0(_gnd_net_),
            .in1(N__24806),
            .in2(N__30117),
            .in3(N__24812),
            .lcout(sEEPeriod_i_1),
            .ltout(),
            .carryin(un4_speriod_cry_0),
            .carryout(un4_speriod_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_2_c_inv_LC_11_6_2.C_ON=1'b1;
    defparam un4_speriod_cry_2_c_inv_LC_11_6_2.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_2_c_inv_LC_11_6_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_2_c_inv_LC_11_6_2 (
            .in0(_gnd_net_),
            .in1(N__24794),
            .in2(N__30006),
            .in3(N__24800),
            .lcout(sEEPeriod_i_2),
            .ltout(),
            .carryin(un4_speriod_cry_1),
            .carryout(un4_speriod_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_3_c_inv_LC_11_6_3.C_ON=1'b1;
    defparam un4_speriod_cry_3_c_inv_LC_11_6_3.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_3_c_inv_LC_11_6_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_3_c_inv_LC_11_6_3 (
            .in0(_gnd_net_),
            .in1(N__24929),
            .in2(N__29877),
            .in3(N__24788),
            .lcout(sEEPeriod_i_3),
            .ltout(),
            .carryin(un4_speriod_cry_2),
            .carryout(un4_speriod_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_4_c_inv_LC_11_6_4.C_ON=1'b1;
    defparam un4_speriod_cry_4_c_inv_LC_11_6_4.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_4_c_inv_LC_11_6_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_4_c_inv_LC_11_6_4 (
            .in0(_gnd_net_),
            .in1(N__24917),
            .in2(N__31016),
            .in3(N__24923),
            .lcout(sEEPeriod_i_4),
            .ltout(),
            .carryin(un4_speriod_cry_3),
            .carryout(un4_speriod_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_5_c_inv_LC_11_6_5.C_ON=1'b1;
    defparam un4_speriod_cry_5_c_inv_LC_11_6_5.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_5_c_inv_LC_11_6_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_speriod_cry_5_c_inv_LC_11_6_5 (
            .in0(N__24911),
            .in1(N__24905),
            .in2(N__30899),
            .in3(_gnd_net_),
            .lcout(sEEPeriod_i_5),
            .ltout(),
            .carryin(un4_speriod_cry_4),
            .carryout(un4_speriod_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_6_c_inv_LC_11_6_6.C_ON=1'b1;
    defparam un4_speriod_cry_6_c_inv_LC_11_6_6.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_6_c_inv_LC_11_6_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_6_c_inv_LC_11_6_6 (
            .in0(_gnd_net_),
            .in1(N__24893),
            .in2(N__30774),
            .in3(N__24899),
            .lcout(sEEPeriod_i_6),
            .ltout(),
            .carryin(un4_speriod_cry_5),
            .carryout(un4_speriod_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_7_c_inv_LC_11_6_7.C_ON=1'b1;
    defparam un4_speriod_cry_7_c_inv_LC_11_6_7.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_7_c_inv_LC_11_6_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_7_c_inv_LC_11_6_7 (
            .in0(_gnd_net_),
            .in1(N__30650),
            .in2(N__24881),
            .in3(N__24887),
            .lcout(sEEPeriod_i_7),
            .ltout(),
            .carryin(un4_speriod_cry_6),
            .carryout(un4_speriod_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_8_c_inv_LC_11_7_0.C_ON=1'b1;
    defparam un4_speriod_cry_8_c_inv_LC_11_7_0.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_8_c_inv_LC_11_7_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_8_c_inv_LC_11_7_0 (
            .in0(_gnd_net_),
            .in1(N__24866),
            .in2(N__30570),
            .in3(N__24872),
            .lcout(sEEPeriod_i_8),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(un4_speriod_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_9_c_inv_LC_11_7_1.C_ON=1'b1;
    defparam un4_speriod_cry_9_c_inv_LC_11_7_1.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_9_c_inv_LC_11_7_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_9_c_inv_LC_11_7_1 (
            .in0(_gnd_net_),
            .in1(N__24854),
            .in2(N__30465),
            .in3(N__24860),
            .lcout(sEEPeriod_i_9),
            .ltout(),
            .carryin(un4_speriod_cry_8),
            .carryout(un4_speriod_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_10_c_inv_LC_11_7_2.C_ON=1'b1;
    defparam un4_speriod_cry_10_c_inv_LC_11_7_2.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_10_c_inv_LC_11_7_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_10_c_inv_LC_11_7_2 (
            .in0(_gnd_net_),
            .in1(N__24842),
            .in2(N__30353),
            .in3(N__24848),
            .lcout(sEEPeriod_i_10),
            .ltout(),
            .carryin(un4_speriod_cry_9),
            .carryout(un4_speriod_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_11_c_inv_LC_11_7_3.C_ON=1'b1;
    defparam un4_speriod_cry_11_c_inv_LC_11_7_3.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_11_c_inv_LC_11_7_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_11_c_inv_LC_11_7_3 (
            .in0(_gnd_net_),
            .in1(N__25019),
            .in2(N__33057),
            .in3(N__25025),
            .lcout(sEEPeriod_i_11),
            .ltout(),
            .carryin(un4_speriod_cry_10),
            .carryout(un4_speriod_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_12_c_inv_LC_11_7_4.C_ON=1'b1;
    defparam un4_speriod_cry_12_c_inv_LC_11_7_4.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_12_c_inv_LC_11_7_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_speriod_cry_12_c_inv_LC_11_7_4 (
            .in0(N__25013),
            .in1(N__25007),
            .in2(N__31733),
            .in3(_gnd_net_),
            .lcout(sEEPeriod_i_12),
            .ltout(),
            .carryin(un4_speriod_cry_11),
            .carryout(un4_speriod_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_13_c_inv_LC_11_7_5.C_ON=1'b1;
    defparam un4_speriod_cry_13_c_inv_LC_11_7_5.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_13_c_inv_LC_11_7_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_speriod_cry_13_c_inv_LC_11_7_5 (
            .in0(N__25001),
            .in1(N__24995),
            .in2(N__31658),
            .in3(_gnd_net_),
            .lcout(sEEPeriod_i_13),
            .ltout(),
            .carryin(un4_speriod_cry_12),
            .carryout(un4_speriod_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_14_c_inv_LC_11_7_6.C_ON=1'b1;
    defparam un4_speriod_cry_14_c_inv_LC_11_7_6.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_14_c_inv_LC_11_7_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_14_c_inv_LC_11_7_6 (
            .in0(_gnd_net_),
            .in1(N__24983),
            .in2(N__31573),
            .in3(N__24989),
            .lcout(sEEPeriod_i_14),
            .ltout(),
            .carryin(un4_speriod_cry_13),
            .carryout(un4_speriod_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_15_c_inv_LC_11_7_7.C_ON=1'b1;
    defparam un4_speriod_cry_15_c_inv_LC_11_7_7.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_15_c_inv_LC_11_7_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_speriod_cry_15_c_inv_LC_11_7_7 (
            .in0(N__24977),
            .in1(N__24971),
            .in2(N__31479),
            .in3(_gnd_net_),
            .lcout(sEEPeriod_i_15),
            .ltout(),
            .carryin(un4_speriod_cry_14),
            .carryout(un4_speriod_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_16_c_inv_LC_11_8_0.C_ON=1'b1;
    defparam un4_speriod_cry_16_c_inv_LC_11_8_0.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_16_c_inv_LC_11_8_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_16_c_inv_LC_11_8_0 (
            .in0(_gnd_net_),
            .in1(N__24959),
            .in2(N__31387),
            .in3(N__24965),
            .lcout(sEEPeriod_i_16),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(un4_speriod_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_17_c_inv_LC_11_8_1.C_ON=1'b1;
    defparam un4_speriod_cry_17_c_inv_LC_11_8_1.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_17_c_inv_LC_11_8_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_17_c_inv_LC_11_8_1 (
            .in0(_gnd_net_),
            .in1(N__24947),
            .in2(N__31286),
            .in3(N__24953),
            .lcout(sEEPeriod_i_17),
            .ltout(),
            .carryin(un4_speriod_cry_16),
            .carryout(un4_speriod_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_18_c_inv_LC_11_8_2.C_ON=1'b1;
    defparam un4_speriod_cry_18_c_inv_LC_11_8_2.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_18_c_inv_LC_11_8_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_18_c_inv_LC_11_8_2 (
            .in0(_gnd_net_),
            .in1(N__24935),
            .in2(N__31177),
            .in3(N__24941),
            .lcout(sEEPeriod_i_18),
            .ltout(),
            .carryin(un4_speriod_cry_17),
            .carryout(un4_speriod_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_19_c_inv_LC_11_8_3.C_ON=1'b1;
    defparam un4_speriod_cry_19_c_inv_LC_11_8_3.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_19_c_inv_LC_11_8_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_19_c_inv_LC_11_8_3 (
            .in0(_gnd_net_),
            .in1(N__25103),
            .in2(N__33278),
            .in3(N__25109),
            .lcout(sEEPeriod_i_19),
            .ltout(),
            .carryin(un4_speriod_cry_18),
            .carryout(un4_speriod_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_20_c_inv_LC_11_8_4.C_ON=1'b1;
    defparam un4_speriod_cry_20_c_inv_LC_11_8_4.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_20_c_inv_LC_11_8_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_20_c_inv_LC_11_8_4 (
            .in0(_gnd_net_),
            .in1(N__25091),
            .in2(N__33380),
            .in3(N__25097),
            .lcout(sEEPeriod_i_20),
            .ltout(),
            .carryin(un4_speriod_cry_19),
            .carryout(un4_speriod_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_21_c_inv_LC_11_8_5.C_ON=1'b1;
    defparam un4_speriod_cry_21_c_inv_LC_11_8_5.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_21_c_inv_LC_11_8_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_speriod_cry_21_c_inv_LC_11_8_5 (
            .in0(N__25085),
            .in1(N__25079),
            .in2(N__33166),
            .in3(_gnd_net_),
            .lcout(sEEPeriod_i_21),
            .ltout(),
            .carryin(un4_speriod_cry_20),
            .carryout(un4_speriod_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_22_c_inv_LC_11_8_6.C_ON=1'b1;
    defparam un4_speriod_cry_22_c_inv_LC_11_8_6.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_22_c_inv_LC_11_8_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_22_c_inv_LC_11_8_6 (
            .in0(_gnd_net_),
            .in1(N__25067),
            .in2(N__32041),
            .in3(N__25073),
            .lcout(sEEPeriod_i_22),
            .ltout(),
            .carryin(un4_speriod_cry_21),
            .carryout(un4_speriod_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_23_c_inv_LC_11_8_7.C_ON=1'b1;
    defparam un4_speriod_cry_23_c_inv_LC_11_8_7.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_23_c_inv_LC_11_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_23_c_inv_LC_11_8_7 (
            .in0(_gnd_net_),
            .in1(N__25055),
            .in2(N__31935),
            .in3(N__25061),
            .lcout(sEEPeriod_i_23),
            .ltout(),
            .carryin(un4_speriod_cry_22),
            .carryout(un4_speriod_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_23_THRU_LUT4_0_LC_11_9_0.C_ON=1'b0;
    defparam un4_speriod_cry_23_THRU_LUT4_0_LC_11_9_0.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_23_THRU_LUT4_0_LC_11_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un4_speriod_cry_23_THRU_LUT4_0_LC_11_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25049),
            .lcout(un4_speriod_cry_23_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sPointer_RNO_0_0_LC_11_9_2.C_ON=1'b0;
    defparam sPointer_RNO_0_0_LC_11_9_2.SEQ_MODE=4'b0000;
    defparam sPointer_RNO_0_0_LC_11_9_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 sPointer_RNO_0_0_LC_11_9_2 (
            .in0(N__46770),
            .in1(N__25964),
            .in2(N__45481),
            .in3(N__25031),
            .lcout(un1_spointer11_2_0_0_a2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sPointer_RNO_1_0_LC_11_9_4.C_ON=1'b0;
    defparam sPointer_RNO_1_0_LC_11_9_4.SEQ_MODE=4'b0000;
    defparam sPointer_RNO_1_0_LC_11_9_4.LUT_INIT=16'b0000000000110011;
    LogicCell40 sPointer_RNO_1_0_LC_11_9_4 (
            .in0(_gnd_net_),
            .in1(N__50305),
            .in2(_gnd_net_),
            .in3(N__47244),
            .lcout(un1_spointer11_2_0_0_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigInternal_RNIMEFL5_LC_11_9_6.C_ON=1'b0;
    defparam sTrigInternal_RNIMEFL5_LC_11_9_6.SEQ_MODE=4'b0000;
    defparam sTrigInternal_RNIMEFL5_LC_11_9_6.LUT_INIT=16'b0101111101001111;
    LogicCell40 sTrigInternal_RNIMEFL5_LC_11_9_6 (
            .in0(N__25214),
            .in1(N__25183),
            .in2(N__49363),
            .in3(N__25152),
            .lcout(LED_ACQ_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_0_LC_11_10_0.C_ON=1'b1;
    defparam sCounter_0_LC_11_10_0.SEQ_MODE=4'b1010;
    defparam sCounter_0_LC_11_10_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_0_LC_11_10_0 (
            .in0(N__25347),
            .in1(N__30206),
            .in2(_gnd_net_),
            .in3(N__25133),
            .lcout(un7_spon_0),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(sCounter_cry_0),
            .clk(N__52262),
            .ce(),
            .sr(N__51689));
    defparam sCounter_1_LC_11_10_1.C_ON=1'b1;
    defparam sCounter_1_LC_11_10_1.SEQ_MODE=4'b1010;
    defparam sCounter_1_LC_11_10_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_1_LC_11_10_1 (
            .in0(N__25360),
            .in1(N__30089),
            .in2(_gnd_net_),
            .in3(N__25130),
            .lcout(un7_spon_1),
            .ltout(),
            .carryin(sCounter_cry_0),
            .carryout(sCounter_cry_1),
            .clk(N__52262),
            .ce(),
            .sr(N__51689));
    defparam sCounter_2_LC_11_10_2.C_ON=1'b1;
    defparam sCounter_2_LC_11_10_2.SEQ_MODE=4'b1010;
    defparam sCounter_2_LC_11_10_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_2_LC_11_10_2 (
            .in0(N__25348),
            .in1(N__29969),
            .in2(_gnd_net_),
            .in3(N__25127),
            .lcout(un7_spon_2),
            .ltout(),
            .carryin(sCounter_cry_1),
            .carryout(sCounter_cry_2),
            .clk(N__52262),
            .ce(),
            .sr(N__51689));
    defparam sCounter_3_LC_11_10_3.C_ON=1'b1;
    defparam sCounter_3_LC_11_10_3.SEQ_MODE=4'b1010;
    defparam sCounter_3_LC_11_10_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_3_LC_11_10_3 (
            .in0(N__25361),
            .in1(N__29840),
            .in2(_gnd_net_),
            .in3(N__25124),
            .lcout(un7_spon_3),
            .ltout(),
            .carryin(sCounter_cry_2),
            .carryout(sCounter_cry_3),
            .clk(N__52262),
            .ce(),
            .sr(N__51689));
    defparam sCounter_4_LC_11_10_4.C_ON=1'b1;
    defparam sCounter_4_LC_11_10_4.SEQ_MODE=4'b1010;
    defparam sCounter_4_LC_11_10_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_4_LC_11_10_4 (
            .in0(N__25349),
            .in1(N__30984),
            .in2(_gnd_net_),
            .in3(N__25121),
            .lcout(un7_spon_4),
            .ltout(),
            .carryin(sCounter_cry_3),
            .carryout(sCounter_cry_4),
            .clk(N__52262),
            .ce(),
            .sr(N__51689));
    defparam sCounter_5_LC_11_10_5.C_ON=1'b1;
    defparam sCounter_5_LC_11_10_5.SEQ_MODE=4'b1010;
    defparam sCounter_5_LC_11_10_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_5_LC_11_10_5 (
            .in0(N__25362),
            .in1(N__30863),
            .in2(_gnd_net_),
            .in3(N__25118),
            .lcout(un7_spon_5),
            .ltout(),
            .carryin(sCounter_cry_4),
            .carryout(sCounter_cry_5),
            .clk(N__52262),
            .ce(),
            .sr(N__51689));
    defparam sCounter_6_LC_11_10_6.C_ON=1'b1;
    defparam sCounter_6_LC_11_10_6.SEQ_MODE=4'b1010;
    defparam sCounter_6_LC_11_10_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_6_LC_11_10_6 (
            .in0(N__25350),
            .in1(N__30752),
            .in2(_gnd_net_),
            .in3(N__25115),
            .lcout(un7_spon_6),
            .ltout(),
            .carryin(sCounter_cry_5),
            .carryout(sCounter_cry_6),
            .clk(N__52262),
            .ce(),
            .sr(N__51689));
    defparam sCounter_7_LC_11_10_7.C_ON=1'b1;
    defparam sCounter_7_LC_11_10_7.SEQ_MODE=4'b1010;
    defparam sCounter_7_LC_11_10_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_7_LC_11_10_7 (
            .in0(N__25363),
            .in1(N__30649),
            .in2(_gnd_net_),
            .in3(N__25112),
            .lcout(un7_spon_7),
            .ltout(),
            .carryin(sCounter_cry_6),
            .carryout(sCounter_cry_7),
            .clk(N__52262),
            .ce(),
            .sr(N__51689));
    defparam sCounter_8_LC_11_11_0.C_ON=1'b1;
    defparam sCounter_8_LC_11_11_0.SEQ_MODE=4'b1010;
    defparam sCounter_8_LC_11_11_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_8_LC_11_11_0 (
            .in0(N__25354),
            .in1(N__30541),
            .in2(_gnd_net_),
            .in3(N__25241),
            .lcout(un7_spon_8),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(sCounter_cry_8),
            .clk(N__52251),
            .ce(),
            .sr(N__51682));
    defparam sCounter_9_LC_11_11_1.C_ON=1'b1;
    defparam sCounter_9_LC_11_11_1.SEQ_MODE=4'b1010;
    defparam sCounter_9_LC_11_11_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_9_LC_11_11_1 (
            .in0(N__25367),
            .in1(N__30426),
            .in2(_gnd_net_),
            .in3(N__25238),
            .lcout(un7_spon_9),
            .ltout(),
            .carryin(sCounter_cry_8),
            .carryout(sCounter_cry_9),
            .clk(N__52251),
            .ce(),
            .sr(N__51682));
    defparam sCounter_10_LC_11_11_2.C_ON=1'b1;
    defparam sCounter_10_LC_11_11_2.SEQ_MODE=4'b1010;
    defparam sCounter_10_LC_11_11_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_10_LC_11_11_2 (
            .in0(N__25351),
            .in1(N__30315),
            .in2(_gnd_net_),
            .in3(N__25235),
            .lcout(un7_spon_10),
            .ltout(),
            .carryin(sCounter_cry_9),
            .carryout(sCounter_cry_10),
            .clk(N__52251),
            .ce(),
            .sr(N__51682));
    defparam sCounter_11_LC_11_11_3.C_ON=1'b1;
    defparam sCounter_11_LC_11_11_3.SEQ_MODE=4'b1010;
    defparam sCounter_11_LC_11_11_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_11_LC_11_11_3 (
            .in0(N__25364),
            .in1(N__33017),
            .in2(_gnd_net_),
            .in3(N__25232),
            .lcout(un7_spon_11),
            .ltout(),
            .carryin(sCounter_cry_10),
            .carryout(sCounter_cry_11),
            .clk(N__52251),
            .ce(),
            .sr(N__51682));
    defparam sCounter_12_LC_11_11_4.C_ON=1'b1;
    defparam sCounter_12_LC_11_11_4.SEQ_MODE=4'b1010;
    defparam sCounter_12_LC_11_11_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_12_LC_11_11_4 (
            .in0(N__25352),
            .in1(N__31718),
            .in2(_gnd_net_),
            .in3(N__25229),
            .lcout(un7_spon_12),
            .ltout(),
            .carryin(sCounter_cry_11),
            .carryout(sCounter_cry_12),
            .clk(N__52251),
            .ce(),
            .sr(N__51682));
    defparam sCounter_13_LC_11_11_5.C_ON=1'b1;
    defparam sCounter_13_LC_11_11_5.SEQ_MODE=4'b1010;
    defparam sCounter_13_LC_11_11_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_13_LC_11_11_5 (
            .in0(N__25365),
            .in1(N__31645),
            .in2(_gnd_net_),
            .in3(N__25226),
            .lcout(un7_spon_13),
            .ltout(),
            .carryin(sCounter_cry_12),
            .carryout(sCounter_cry_13),
            .clk(N__52251),
            .ce(),
            .sr(N__51682));
    defparam sCounter_14_LC_11_11_6.C_ON=1'b1;
    defparam sCounter_14_LC_11_11_6.SEQ_MODE=4'b1010;
    defparam sCounter_14_LC_11_11_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_14_LC_11_11_6 (
            .in0(N__25353),
            .in1(N__31537),
            .in2(_gnd_net_),
            .in3(N__25223),
            .lcout(un7_spon_14),
            .ltout(),
            .carryin(sCounter_cry_13),
            .carryout(sCounter_cry_14),
            .clk(N__52251),
            .ce(),
            .sr(N__51682));
    defparam sCounter_15_LC_11_11_7.C_ON=1'b1;
    defparam sCounter_15_LC_11_11_7.SEQ_MODE=4'b1010;
    defparam sCounter_15_LC_11_11_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_15_LC_11_11_7 (
            .in0(N__25366),
            .in1(N__31450),
            .in2(_gnd_net_),
            .in3(N__25220),
            .lcout(un7_spon_15),
            .ltout(),
            .carryin(sCounter_cry_14),
            .carryout(sCounter_cry_15),
            .clk(N__52251),
            .ce(),
            .sr(N__51682));
    defparam sCounter_16_LC_11_12_0.C_ON=1'b1;
    defparam sCounter_16_LC_11_12_0.SEQ_MODE=4'b1010;
    defparam sCounter_16_LC_11_12_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_16_LC_11_12_0 (
            .in0(N__25355),
            .in1(N__31337),
            .in2(_gnd_net_),
            .in3(N__25217),
            .lcout(un7_spon_16),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(sCounter_cry_16),
            .clk(N__52263),
            .ce(),
            .sr(N__51676));
    defparam sCounter_17_LC_11_12_1.C_ON=1'b1;
    defparam sCounter_17_LC_11_12_1.SEQ_MODE=4'b1010;
    defparam sCounter_17_LC_11_12_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_17_LC_11_12_1 (
            .in0(N__25368),
            .in1(N__31261),
            .in2(_gnd_net_),
            .in3(N__25388),
            .lcout(un7_spon_17),
            .ltout(),
            .carryin(sCounter_cry_16),
            .carryout(sCounter_cry_17),
            .clk(N__52263),
            .ce(),
            .sr(N__51676));
    defparam sCounter_18_LC_11_12_2.C_ON=1'b1;
    defparam sCounter_18_LC_11_12_2.SEQ_MODE=4'b1010;
    defparam sCounter_18_LC_11_12_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_18_LC_11_12_2 (
            .in0(N__25356),
            .in1(N__31124),
            .in2(_gnd_net_),
            .in3(N__25385),
            .lcout(un7_spon_18),
            .ltout(),
            .carryin(sCounter_cry_17),
            .carryout(sCounter_cry_18),
            .clk(N__52263),
            .ce(),
            .sr(N__51676));
    defparam sCounter_19_LC_11_12_3.C_ON=1'b1;
    defparam sCounter_19_LC_11_12_3.SEQ_MODE=4'b1010;
    defparam sCounter_19_LC_11_12_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_19_LC_11_12_3 (
            .in0(N__25369),
            .in1(N__33224),
            .in2(_gnd_net_),
            .in3(N__25382),
            .lcout(un7_spon_19),
            .ltout(),
            .carryin(sCounter_cry_18),
            .carryout(sCounter_cry_19),
            .clk(N__52263),
            .ce(),
            .sr(N__51676));
    defparam sCounter_20_LC_11_12_4.C_ON=1'b1;
    defparam sCounter_20_LC_11_12_4.SEQ_MODE=4'b1010;
    defparam sCounter_20_LC_11_12_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_20_LC_11_12_4 (
            .in0(N__25357),
            .in1(N__33331),
            .in2(_gnd_net_),
            .in3(N__25379),
            .lcout(un7_spon_20),
            .ltout(),
            .carryin(sCounter_cry_19),
            .carryout(sCounter_cry_20),
            .clk(N__52263),
            .ce(),
            .sr(N__51676));
    defparam sCounter_21_LC_11_12_5.C_ON=1'b1;
    defparam sCounter_21_LC_11_12_5.SEQ_MODE=4'b1010;
    defparam sCounter_21_LC_11_12_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_21_LC_11_12_5 (
            .in0(N__25370),
            .in1(N__33115),
            .in2(_gnd_net_),
            .in3(N__25376),
            .lcout(un7_spon_21),
            .ltout(),
            .carryin(sCounter_cry_20),
            .carryout(sCounter_cry_21),
            .clk(N__52263),
            .ce(),
            .sr(N__51676));
    defparam sCounter_22_LC_11_12_6.C_ON=1'b1;
    defparam sCounter_22_LC_11_12_6.SEQ_MODE=4'b1010;
    defparam sCounter_22_LC_11_12_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_22_LC_11_12_6 (
            .in0(N__25358),
            .in1(N__31991),
            .in2(_gnd_net_),
            .in3(N__25373),
            .lcout(un7_spon_22),
            .ltout(),
            .carryin(sCounter_cry_21),
            .carryout(sCounter_cry_22),
            .clk(N__52263),
            .ce(),
            .sr(N__51676));
    defparam sCounter_23_LC_11_12_7.C_ON=1'b0;
    defparam sCounter_23_LC_11_12_7.SEQ_MODE=4'b1010;
    defparam sCounter_23_LC_11_12_7.LUT_INIT=16'b0001000100100010;
    LogicCell40 sCounter_23_LC_11_12_7 (
            .in0(N__31882),
            .in1(N__25359),
            .in2(_gnd_net_),
            .in3(N__25274),
            .lcout(un7_spon_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52263),
            .ce(),
            .sr(N__51676));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_0_LC_11_13_0 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_0_LC_11_13_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_0_LC_11_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_0_LC_11_13_0  (
            .in0(N__27927),
            .in1(N__25271),
            .in2(_gnd_net_),
            .in3(N__25259),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0 ),
            .clk(N__48472),
            .ce(N__27968),
            .sr(N__51668));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_1_LC_11_13_1 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_1_LC_11_13_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_1_LC_11_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_1_LC_11_13_1  (
            .in0(N__27922),
            .in1(N__25256),
            .in2(_gnd_net_),
            .in3(N__25244),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1 ),
            .clk(N__48472),
            .ce(N__27968),
            .sr(N__51668));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_2_LC_11_13_2 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_2_LC_11_13_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_2_LC_11_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_2_LC_11_13_2  (
            .in0(N__27928),
            .in1(N__25490),
            .in2(_gnd_net_),
            .in3(N__25478),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2 ),
            .clk(N__48472),
            .ce(N__27968),
            .sr(N__51668));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_3_LC_11_13_3 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_3_LC_11_13_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_3_LC_11_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_3_LC_11_13_3  (
            .in0(N__27923),
            .in1(N__25475),
            .in2(_gnd_net_),
            .in3(N__25463),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3 ),
            .clk(N__48472),
            .ce(N__27968),
            .sr(N__51668));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_4_LC_11_13_4 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_4_LC_11_13_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_4_LC_11_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_4_LC_11_13_4  (
            .in0(N__27929),
            .in1(N__25453),
            .in2(_gnd_net_),
            .in3(N__25439),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4 ),
            .clk(N__48472),
            .ce(N__27968),
            .sr(N__51668));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_5_LC_11_13_5 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_5_LC_11_13_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_5_LC_11_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_5_LC_11_13_5  (
            .in0(N__27924),
            .in1(N__25435),
            .in2(_gnd_net_),
            .in3(N__25421),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5 ),
            .clk(N__48472),
            .ce(N__27968),
            .sr(N__51668));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_6_LC_11_13_6 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_6_LC_11_13_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_6_LC_11_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_6_LC_11_13_6  (
            .in0(N__27925),
            .in1(N__25418),
            .in2(_gnd_net_),
            .in3(N__25406),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6 ),
            .clk(N__48472),
            .ce(N__27968),
            .sr(N__51668));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_7_LC_11_13_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_7_LC_11_13_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_7_LC_11_13_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_7_LC_11_13_7  (
            .in0(N__25400),
            .in1(N__27926),
            .in2(_gnd_net_),
            .in3(N__25403),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48472),
            .ce(N__27968),
            .sr(N__51668));
    defparam sEEPoff_0_LC_11_14_0.C_ON=1'b0;
    defparam sEEPoff_0_LC_11_14_0.SEQ_MODE=4'b1010;
    defparam sEEPoff_0_LC_11_14_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPoff_0_LC_11_14_0 (
            .in0(N__46342),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPoffZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52284),
            .ce(N__25496),
            .sr(N__51662));
    defparam sEEPoff_1_LC_11_14_1.C_ON=1'b0;
    defparam sEEPoff_1_LC_11_14_1.SEQ_MODE=4'b1010;
    defparam sEEPoff_1_LC_11_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_1_LC_11_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50879),
            .lcout(sEEPoffZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52284),
            .ce(N__25496),
            .sr(N__51662));
    defparam sEEPoff_2_LC_11_14_2.C_ON=1'b0;
    defparam sEEPoff_2_LC_11_14_2.SEQ_MODE=4'b1010;
    defparam sEEPoff_2_LC_11_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_2_LC_11_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47501),
            .lcout(sEEPoffZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52284),
            .ce(N__25496),
            .sr(N__51662));
    defparam sEEPoff_3_LC_11_14_3.C_ON=1'b0;
    defparam sEEPoff_3_LC_11_14_3.SEQ_MODE=4'b1011;
    defparam sEEPoff_3_LC_11_14_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPoff_3_LC_11_14_3 (
            .in0(N__46914),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPoffZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52284),
            .ce(N__25496),
            .sr(N__51662));
    defparam sEEPoff_4_LC_11_14_4.C_ON=1'b0;
    defparam sEEPoff_4_LC_11_14_4.SEQ_MODE=4'b1010;
    defparam sEEPoff_4_LC_11_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_4_LC_11_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45567),
            .lcout(sEEPoffZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52284),
            .ce(N__25496),
            .sr(N__51662));
    defparam sEEPoff_5_LC_11_14_5.C_ON=1'b0;
    defparam sEEPoff_5_LC_11_14_5.SEQ_MODE=4'b1010;
    defparam sEEPoff_5_LC_11_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_5_LC_11_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45089),
            .lcout(sEEPoffZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52284),
            .ce(N__25496),
            .sr(N__51662));
    defparam sEEPoff_6_LC_11_14_6.C_ON=1'b0;
    defparam sEEPoff_6_LC_11_14_6.SEQ_MODE=4'b1011;
    defparam sEEPoff_6_LC_11_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_6_LC_11_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50530),
            .lcout(sEEPoffZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52284),
            .ce(N__25496),
            .sr(N__51662));
    defparam sEEPoff_7_LC_11_14_7.C_ON=1'b0;
    defparam sEEPoff_7_LC_11_14_7.SEQ_MODE=4'b1011;
    defparam sEEPoff_7_LC_11_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_7_LC_11_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50030),
            .lcout(sEEPoffZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52284),
            .ce(N__25496),
            .sr(N__51662));
    defparam sAddress_RNIA6242_0_0_LC_11_15_0.C_ON=1'b0;
    defparam sAddress_RNIA6242_0_0_LC_11_15_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_0_0_LC_11_15_0.LUT_INIT=16'b0000000010000000;
    LogicCell40 sAddress_RNIA6242_0_0_LC_11_15_0 (
            .in0(N__40190),
            .in1(N__25521),
            .in2(N__40669),
            .in3(N__40433),
            .lcout(sAddress_RNIA6242_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_1_0_LC_11_15_1.C_ON=1'b0;
    defparam sAddress_RNIA6242_1_0_LC_11_15_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_1_0_LC_11_15_1.LUT_INIT=16'b0000000000001000;
    LogicCell40 sAddress_RNIA6242_1_0_LC_11_15_1 (
            .in0(N__25520),
            .in1(N__40654),
            .in2(N__40438),
            .in3(N__40189),
            .lcout(sAddress_RNIA6242_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_2_0_LC_11_15_2.C_ON=1'b0;
    defparam sAddress_RNIA6242_2_0_LC_11_15_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_2_0_LC_11_15_2.LUT_INIT=16'b0000000000100000;
    LogicCell40 sAddress_RNIA6242_2_0_LC_11_15_2 (
            .in0(N__25523),
            .in1(N__40659),
            .in2(N__40199),
            .in3(N__40437),
            .lcout(sAddress_RNIA6242_2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_3_0_LC_11_15_3.C_ON=1'b0;
    defparam sAddress_RNIA6242_3_0_LC_11_15_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_3_0_LC_11_15_3.LUT_INIT=16'b0000000000000010;
    LogicCell40 sAddress_RNIA6242_3_0_LC_11_15_3 (
            .in0(N__25522),
            .in1(N__40658),
            .in2(N__40439),
            .in3(N__40191),
            .lcout(sAddress_RNIA6242_3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI6VH7_4_1_LC_11_15_4.C_ON=1'b0;
    defparam sAddress_RNI6VH7_4_1_LC_11_15_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI6VH7_4_1_LC_11_15_4.LUT_INIT=16'b0000001000000010;
    LogicCell40 sAddress_RNI6VH7_4_1_LC_11_15_4 (
            .in0(N__40653),
            .in1(N__40545),
            .in2(N__40198),
            .in3(_gnd_net_),
            .lcout(sAddress_RNI6VH7_4Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPoff_10_LC_11_15_5.C_ON=1'b0;
    defparam sEEPoff_10_LC_11_15_5.SEQ_MODE=4'b1010;
    defparam sEEPoff_10_LC_11_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_10_LC_11_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47459),
            .lcout(sEEPoffZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52296),
            .ce(N__26755),
            .sr(N__51656));
    defparam sbuttonModeStatus_RNO_3_LC_11_16_2.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_3_LC_11_16_2.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_3_LC_11_16_2.LUT_INIT=16'b1010101000000000;
    LogicCell40 sbuttonModeStatus_RNO_3_LC_11_16_2 (
            .in0(N__49095),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35312),
            .lcout(sbuttonModeStatus_0_sqmuxa_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_0_c_inv_LC_11_17_0.C_ON=1'b1;
    defparam un4_sacqtime_cry_0_c_inv_LC_11_17_0.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_0_c_inv_LC_11_17_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_0_c_inv_LC_11_17_0 (
            .in0(_gnd_net_),
            .in1(N__25592),
            .in2(N__30229),
            .in3(N__25598),
            .lcout(sEEDelayACQ_i_0),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(un4_sacqtime_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_1_c_inv_LC_11_17_1.C_ON=1'b1;
    defparam un4_sacqtime_cry_1_c_inv_LC_11_17_1.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_1_c_inv_LC_11_17_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_sacqtime_cry_1_c_inv_LC_11_17_1 (
            .in0(N__25586),
            .in1(N__25580),
            .in2(N__30109),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQ_i_1),
            .ltout(),
            .carryin(un4_sacqtime_cry_0),
            .carryout(un4_sacqtime_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_2_c_inv_LC_11_17_2.C_ON=1'b1;
    defparam un4_sacqtime_cry_2_c_inv_LC_11_17_2.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_2_c_inv_LC_11_17_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_sacqtime_cry_2_c_inv_LC_11_17_2 (
            .in0(N__25574),
            .in1(N__25568),
            .in2(N__29996),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQ_i_2),
            .ltout(),
            .carryin(un4_sacqtime_cry_1),
            .carryout(un4_sacqtime_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_3_c_inv_LC_11_17_3.C_ON=1'b1;
    defparam un4_sacqtime_cry_3_c_inv_LC_11_17_3.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_3_c_inv_LC_11_17_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_3_c_inv_LC_11_17_3 (
            .in0(_gnd_net_),
            .in1(N__29867),
            .in2(N__25556),
            .in3(N__25562),
            .lcout(sEEDelayACQ_i_3),
            .ltout(),
            .carryin(un4_sacqtime_cry_2),
            .carryout(un4_sacqtime_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_4_c_inv_LC_11_17_4.C_ON=1'b1;
    defparam un4_sacqtime_cry_4_c_inv_LC_11_17_4.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_4_c_inv_LC_11_17_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_4_c_inv_LC_11_17_4 (
            .in0(_gnd_net_),
            .in1(N__25541),
            .in2(N__31038),
            .in3(N__25547),
            .lcout(sEEDelayACQ_i_4),
            .ltout(),
            .carryin(un4_sacqtime_cry_3),
            .carryout(un4_sacqtime_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_5_c_inv_LC_11_17_5.C_ON=1'b1;
    defparam un4_sacqtime_cry_5_c_inv_LC_11_17_5.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_5_c_inv_LC_11_17_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_5_c_inv_LC_11_17_5 (
            .in0(_gnd_net_),
            .in1(N__25529),
            .in2(N__30900),
            .in3(N__25535),
            .lcout(sEEDelayACQ_i_5),
            .ltout(),
            .carryin(un4_sacqtime_cry_4),
            .carryout(un4_sacqtime_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_6_c_inv_LC_11_17_6.C_ON=1'b1;
    defparam un4_sacqtime_cry_6_c_inv_LC_11_17_6.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_6_c_inv_LC_11_17_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_6_c_inv_LC_11_17_6 (
            .in0(_gnd_net_),
            .in1(N__25691),
            .in2(N__30786),
            .in3(N__25697),
            .lcout(sEEDelayACQ_i_6),
            .ltout(),
            .carryin(un4_sacqtime_cry_5),
            .carryout(un4_sacqtime_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_7_c_inv_LC_11_17_7.C_ON=1'b1;
    defparam un4_sacqtime_cry_7_c_inv_LC_11_17_7.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_7_c_inv_LC_11_17_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_7_c_inv_LC_11_17_7 (
            .in0(_gnd_net_),
            .in1(N__30651),
            .in2(N__25679),
            .in3(N__25685),
            .lcout(sEEDelayACQ_i_7),
            .ltout(),
            .carryin(un4_sacqtime_cry_6),
            .carryout(un4_sacqtime_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_8_c_inv_LC_11_18_0.C_ON=1'b1;
    defparam un4_sacqtime_cry_8_c_inv_LC_11_18_0.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_8_c_inv_LC_11_18_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_8_c_inv_LC_11_18_0 (
            .in0(_gnd_net_),
            .in1(N__25664),
            .in2(N__30562),
            .in3(N__25670),
            .lcout(sEEDelayACQ_i_8),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(un4_sacqtime_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_9_c_inv_LC_11_18_1.C_ON=1'b1;
    defparam un4_sacqtime_cry_9_c_inv_LC_11_18_1.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_9_c_inv_LC_11_18_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_9_c_inv_LC_11_18_1 (
            .in0(_gnd_net_),
            .in1(N__25652),
            .in2(N__30456),
            .in3(N__25658),
            .lcout(sEEDelayACQ_i_9),
            .ltout(),
            .carryin(un4_sacqtime_cry_8),
            .carryout(un4_sacqtime_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_10_c_inv_LC_11_18_2.C_ON=1'b1;
    defparam un4_sacqtime_cry_10_c_inv_LC_11_18_2.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_10_c_inv_LC_11_18_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_10_c_inv_LC_11_18_2 (
            .in0(_gnd_net_),
            .in1(N__25640),
            .in2(N__30341),
            .in3(N__25646),
            .lcout(sEEDelayACQ_i_10),
            .ltout(),
            .carryin(un4_sacqtime_cry_9),
            .carryout(un4_sacqtime_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_11_c_inv_LC_11_18_3.C_ON=1'b1;
    defparam un4_sacqtime_cry_11_c_inv_LC_11_18_3.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_11_c_inv_LC_11_18_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_11_c_inv_LC_11_18_3 (
            .in0(_gnd_net_),
            .in1(N__25628),
            .in2(N__33046),
            .in3(N__25634),
            .lcout(sEEDelayACQ_i_11),
            .ltout(),
            .carryin(un4_sacqtime_cry_10),
            .carryout(un4_sacqtime_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_12_c_inv_LC_11_18_4.C_ON=1'b1;
    defparam un4_sacqtime_cry_12_c_inv_LC_11_18_4.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_12_c_inv_LC_11_18_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_sacqtime_cry_12_c_inv_LC_11_18_4 (
            .in0(N__25622),
            .in1(N__25616),
            .in2(N__31743),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQ_i_12),
            .ltout(),
            .carryin(un4_sacqtime_cry_11),
            .carryout(un4_sacqtime_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_13_c_inv_LC_11_18_5.C_ON=1'b1;
    defparam un4_sacqtime_cry_13_c_inv_LC_11_18_5.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_13_c_inv_LC_11_18_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_sacqtime_cry_13_c_inv_LC_11_18_5 (
            .in0(N__25610),
            .in1(N__25604),
            .in2(N__31659),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQ_i_13),
            .ltout(),
            .carryin(un4_sacqtime_cry_12),
            .carryout(un4_sacqtime_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_14_c_inv_LC_11_18_6.C_ON=1'b1;
    defparam un4_sacqtime_cry_14_c_inv_LC_11_18_6.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_14_c_inv_LC_11_18_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_14_c_inv_LC_11_18_6 (
            .in0(_gnd_net_),
            .in1(N__25733),
            .in2(N__31574),
            .in3(N__25739),
            .lcout(sEEDelayACQ_i_14),
            .ltout(),
            .carryin(un4_sacqtime_cry_13),
            .carryout(un4_sacqtime_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_15_c_inv_LC_11_18_7.C_ON=1'b1;
    defparam un4_sacqtime_cry_15_c_inv_LC_11_18_7.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_15_c_inv_LC_11_18_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_sacqtime_cry_15_c_inv_LC_11_18_7 (
            .in0(N__25727),
            .in1(N__31472),
            .in2(N__25721),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQ_i_15),
            .ltout(),
            .carryin(un4_sacqtime_cry_14),
            .carryout(un4_sacqtime_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_16_c_LC_11_19_0.C_ON=1'b1;
    defparam un4_sacqtime_cry_16_c_LC_11_19_0.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_16_c_LC_11_19_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_16_c_LC_11_19_0 (
            .in0(_gnd_net_),
            .in1(N__31388),
            .in2(N__52709),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(un4_sacqtime_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_17_c_LC_11_19_1.C_ON=1'b1;
    defparam un4_sacqtime_cry_17_c_LC_11_19_1.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_17_c_LC_11_19_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_17_c_LC_11_19_1 (
            .in0(_gnd_net_),
            .in1(N__31266),
            .in2(N__52707),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_sacqtime_cry_16),
            .carryout(un4_sacqtime_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_18_c_LC_11_19_2.C_ON=1'b1;
    defparam un4_sacqtime_cry_18_c_LC_11_19_2.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_18_c_LC_11_19_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_18_c_LC_11_19_2 (
            .in0(_gnd_net_),
            .in1(N__31149),
            .in2(N__52710),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_sacqtime_cry_17),
            .carryout(un4_sacqtime_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_19_c_LC_11_19_3.C_ON=1'b1;
    defparam un4_sacqtime_cry_19_c_LC_11_19_3.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_19_c_LC_11_19_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_19_c_LC_11_19_3 (
            .in0(_gnd_net_),
            .in1(N__33249),
            .in2(N__52708),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_sacqtime_cry_18),
            .carryout(un4_sacqtime_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_20_c_LC_11_19_4.C_ON=1'b1;
    defparam un4_sacqtime_cry_20_c_LC_11_19_4.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_20_c_LC_11_19_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_20_c_LC_11_19_4 (
            .in0(_gnd_net_),
            .in1(N__52639),
            .in2(N__33381),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_sacqtime_cry_19),
            .carryout(un4_sacqtime_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIR3KA_20_LC_11_19_5.C_ON=1'b1;
    defparam sCounter_RNIR3KA_20_LC_11_19_5.SEQ_MODE=4'b0000;
    defparam sCounter_RNIR3KA_20_LC_11_19_5.LUT_INIT=16'b0000000000110011;
    LogicCell40 sCounter_RNIR3KA_20_LC_11_19_5 (
            .in0(_gnd_net_),
            .in1(N__33150),
            .in2(N__52705),
            .in3(N__33366),
            .lcout(g1_i_a4_4),
            .ltout(),
            .carryin(un4_sacqtime_cry_20),
            .carryout(un4_sacqtime_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_22_c_LC_11_19_6.C_ON=1'b1;
    defparam un4_sacqtime_cry_22_c_LC_11_19_6.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_22_c_LC_11_19_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_22_c_LC_11_19_6 (
            .in0(_gnd_net_),
            .in1(N__32020),
            .in2(N__52711),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_sacqtime_cry_21),
            .carryout(un4_sacqtime_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIV7KA_23_LC_11_19_7.C_ON=1'b1;
    defparam sCounter_RNIV7KA_23_LC_11_19_7.SEQ_MODE=4'b0000;
    defparam sCounter_RNIV7KA_23_LC_11_19_7.LUT_INIT=16'b0000000000110011;
    LogicCell40 sCounter_RNIV7KA_23_LC_11_19_7 (
            .in0(_gnd_net_),
            .in1(N__31909),
            .in2(N__52706),
            .in3(N__32019),
            .lcout(g0_4_0),
            .ltout(),
            .carryin(un4_sacqtime_cry_22),
            .carryout(un4_sacqtime_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_23_THRU_LUT4_0_LC_11_20_0.C_ON=1'b0;
    defparam un4_sacqtime_cry_23_THRU_LUT4_0_LC_11_20_0.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_23_THRU_LUT4_0_LC_11_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un4_sacqtime_cry_23_THRU_LUT4_0_LC_11_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25835),
            .lcout(un4_sacqtime_cry_23_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam spi_sclk_inferred_clock_RNO_LC_12_1_2.C_ON=1'b0;
    defparam spi_sclk_inferred_clock_RNO_LC_12_1_2.SEQ_MODE=4'b0000;
    defparam spi_sclk_inferred_clock_RNO_LC_12_1_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 spi_sclk_inferred_clock_RNO_LC_12_1_2 (
            .in0(N__48032),
            .in1(N__25832),
            .in2(_gnd_net_),
            .in3(N__25817),
            .lcout(spi_sclk),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_3_LC_12_3_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_3_LC_12_3_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_3_LC_12_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_3_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31802),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48444),
            .ce(),
            .sr(N__51750));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_12_LC_12_3_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_12_LC_12_3_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_12_LC_12_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_12_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25778),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48444),
            .ce(),
            .sr(N__51750));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_7_LC_12_3_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_7_LC_12_3_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_7_LC_12_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_7_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31769),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48444),
            .ce(),
            .sr(N__51750));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_9_LC_12_3_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_9_LC_12_3_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_9_LC_12_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_9_LC_12_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32120),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48444),
            .ce(),
            .sr(N__51750));
    defparam sDAC_mem_8_0_LC_12_4_0.C_ON=1'b0;
    defparam sDAC_mem_8_0_LC_12_4_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_0_LC_12_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_0_LC_12_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46147),
            .lcout(sDAC_mem_8Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52320),
            .ce(N__27116),
            .sr(N__51737));
    defparam sDAC_mem_8_1_LC_12_4_1.C_ON=1'b0;
    defparam sDAC_mem_8_1_LC_12_4_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_1_LC_12_4_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_8_1_LC_12_4_1 (
            .in0(N__50939),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_8Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52320),
            .ce(N__27116),
            .sr(N__51737));
    defparam sDAC_mem_8_2_LC_12_4_2.C_ON=1'b0;
    defparam sDAC_mem_8_2_LC_12_4_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_2_LC_12_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_2_LC_12_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47251),
            .lcout(sDAC_mem_8Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52320),
            .ce(N__27116),
            .sr(N__51737));
    defparam sDAC_mem_8_3_LC_12_4_3.C_ON=1'b0;
    defparam sDAC_mem_8_3_LC_12_4_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_3_LC_12_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_3_LC_12_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46707),
            .lcout(sDAC_mem_8Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52320),
            .ce(N__27116),
            .sr(N__51737));
    defparam sDAC_mem_8_4_LC_12_4_4.C_ON=1'b0;
    defparam sDAC_mem_8_4_LC_12_4_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_4_LC_12_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_4_LC_12_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45397),
            .lcout(sDAC_mem_8Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52320),
            .ce(N__27116),
            .sr(N__51737));
    defparam sDAC_mem_8_5_LC_12_4_5.C_ON=1'b0;
    defparam sDAC_mem_8_5_LC_12_4_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_5_LC_12_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_5_LC_12_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45005),
            .lcout(sDAC_mem_8Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52320),
            .ce(N__27116),
            .sr(N__51737));
    defparam sDAC_mem_8_6_LC_12_4_6.C_ON=1'b0;
    defparam sDAC_mem_8_6_LC_12_4_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_6_LC_12_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_6_LC_12_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50413),
            .lcout(sDAC_mem_8Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52320),
            .ce(N__27116),
            .sr(N__51737));
    defparam sDAC_mem_8_7_LC_12_4_7.C_ON=1'b0;
    defparam sDAC_mem_8_7_LC_12_4_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_7_LC_12_4_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_7_LC_12_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49893),
            .lcout(sDAC_mem_8Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52320),
            .ce(N__27116),
            .sr(N__51737));
    defparam sDAC_mem_3_3_LC_12_5_0.C_ON=1'b0;
    defparam sDAC_mem_3_3_LC_12_5_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_3_LC_12_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_3_3_LC_12_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46689),
            .lcout(sDAC_mem_3Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52308),
            .ce(N__44238),
            .sr(N__51723));
    defparam sDAC_data_RNO_27_6_LC_12_5_1.C_ON=1'b0;
    defparam sDAC_data_RNO_27_6_LC_12_5_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_6_LC_12_5_1.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_27_6_LC_12_5_1 (
            .in0(N__42588),
            .in1(N__25991),
            .in2(N__42249),
            .in3(N__25877),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_6_LC_12_5_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_6_LC_12_5_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_6_LC_12_5_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_6_LC_12_5_2 (
            .in0(N__42229),
            .in1(N__25871),
            .in2(N__25859),
            .in3(N__25856),
            .lcout(sDAC_data_RNO_15Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_6_LC_12_5_3.C_ON=1'b0;
    defparam sDAC_data_RNO_16_6_LC_12_5_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_6_LC_12_5_3.LUT_INIT=16'b0000110100111101;
    LogicCell40 sDAC_data_RNO_16_6_LC_12_5_3 (
            .in0(N__25928),
            .in1(N__42230),
            .in2(N__42595),
            .in3(N__26804),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_6_LC_12_5_4.C_ON=1'b0;
    defparam sDAC_data_RNO_7_6_LC_12_5_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_6_LC_12_5_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_7_6_LC_12_5_4 (
            .in0(N__42231),
            .in1(N__39872),
            .in2(N__25922),
            .in3(N__36815),
            .lcout(sDAC_data_RNO_7Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_6_LC_12_5_5.C_ON=1'b0;
    defparam sDAC_data_RNO_17_6_LC_12_5_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_6_LC_12_5_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 sDAC_data_RNO_17_6_LC_12_5_5 (
            .in0(N__25919),
            .in1(_gnd_net_),
            .in2(N__42596),
            .in3(N__25910),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_6_LC_12_5_6.C_ON=1'b0;
    defparam sDAC_data_RNO_8_6_LC_12_5_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_6_LC_12_5_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_8_6_LC_12_5_6 (
            .in0(_gnd_net_),
            .in1(N__42218),
            .in2(N__25901),
            .in3(N__25898),
            .lcout(),
            .ltout(sDAC_data_RNO_8Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_6_LC_12_5_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_6_LC_12_5_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_6_LC_12_5_7.LUT_INIT=16'b0111011000110010;
    LogicCell40 sDAC_data_RNO_2_6_LC_12_5_7 (
            .in0(N__38252),
            .in1(N__28859),
            .in2(N__25886),
            .in3(N__25883),
            .lcout(sDAC_data_RNO_2Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_2_0_LC_12_6_0.C_ON=1'b0;
    defparam sDAC_mem_2_0_LC_12_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_0_LC_12_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_0_LC_12_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46146),
            .lcout(sDAC_mem_2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52297),
            .ce(N__32851),
            .sr(N__51713));
    defparam sDAC_mem_2_1_LC_12_6_1.C_ON=1'b0;
    defparam sDAC_mem_2_1_LC_12_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_1_LC_12_6_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_2_1_LC_12_6_1 (
            .in0(N__50938),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_2Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52297),
            .ce(N__32851),
            .sr(N__51713));
    defparam sDAC_mem_2_2_LC_12_6_2.C_ON=1'b0;
    defparam sDAC_mem_2_2_LC_12_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_2_LC_12_6_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_2_2_LC_12_6_2 (
            .in0(N__47245),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52297),
            .ce(N__32851),
            .sr(N__51713));
    defparam sDAC_mem_2_3_LC_12_6_3.C_ON=1'b0;
    defparam sDAC_mem_2_3_LC_12_6_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_3_LC_12_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_3_LC_12_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46709),
            .lcout(sDAC_mem_2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52297),
            .ce(N__32851),
            .sr(N__51713));
    defparam sDAC_mem_2_4_LC_12_6_4.C_ON=1'b0;
    defparam sDAC_mem_2_4_LC_12_6_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_4_LC_12_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_4_LC_12_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45372),
            .lcout(sDAC_mem_2Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52297),
            .ce(N__32851),
            .sr(N__51713));
    defparam sDAC_mem_2_5_LC_12_6_5.C_ON=1'b0;
    defparam sDAC_mem_2_5_LC_12_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_5_LC_12_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_5_LC_12_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44840),
            .lcout(sDAC_mem_2Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52297),
            .ce(N__32851),
            .sr(N__51713));
    defparam sDAC_mem_2_6_LC_12_6_6.C_ON=1'b0;
    defparam sDAC_mem_2_6_LC_12_6_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_6_LC_12_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_6_LC_12_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50334),
            .lcout(sDAC_mem_2Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52297),
            .ce(N__32851),
            .sr(N__51713));
    defparam sDAC_data_RNO_5_4_LC_12_7_0.C_ON=1'b0;
    defparam sDAC_data_RNO_5_4_LC_12_7_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_4_LC_12_7_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_5_4_LC_12_7_0 (
            .in0(N__26249),
            .in1(N__25970),
            .in2(N__42266),
            .in3(N__32564),
            .lcout(sDAC_data_RNO_5Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_7_1_LC_12_7_1.C_ON=1'b0;
    defparam sDAC_mem_7_1_LC_12_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_1_LC_12_7_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_7_1_LC_12_7_1 (
            .in0(N__50816),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_7Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52285),
            .ce(N__44278),
            .sr(N__51702));
    defparam sPointer_RNO_2_0_LC_12_7_2.C_ON=1'b0;
    defparam sPointer_RNO_2_0_LC_12_7_2.SEQ_MODE=4'b0000;
    defparam sPointer_RNO_2_0_LC_12_7_2.LUT_INIT=16'b0000000010000000;
    LogicCell40 sPointer_RNO_2_0_LC_12_7_2 (
            .in0(N__44833),
            .in1(N__50815),
            .in2(N__49994),
            .in3(N__46051),
            .lcout(un1_spointer11_2_0_0_a2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_7_0_LC_12_7_3.C_ON=1'b0;
    defparam sDAC_mem_7_0_LC_12_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_0_LC_12_7_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_7_0_LC_12_7_3 (
            .in0(N__46053),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_7Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52285),
            .ce(N__44278),
            .sr(N__51702));
    defparam sDAC_mem_7_5_LC_12_7_4.C_ON=1'b0;
    defparam sDAC_mem_7_5_LC_12_7_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_5_LC_12_7_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_7_5_LC_12_7_4 (
            .in0(N__44834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_7Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52285),
            .ce(N__44278),
            .sr(N__51702));
    defparam sDAC_mem_7_7_LC_12_7_5.C_ON=1'b0;
    defparam sDAC_mem_7_7_LC_12_7_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_7_LC_12_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_7_7_LC_12_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49892),
            .lcout(sDAC_mem_7Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52285),
            .ce(N__44278),
            .sr(N__51702));
    defparam sPointer_RNIV9N7_1_LC_12_7_6.C_ON=1'b0;
    defparam sPointer_RNIV9N7_1_LC_12_7_6.SEQ_MODE=4'b0000;
    defparam sPointer_RNIV9N7_1_LC_12_7_6.LUT_INIT=16'b0011001111111111;
    LogicCell40 sPointer_RNIV9N7_1_LC_12_7_6 (
            .in0(_gnd_net_),
            .in1(N__46052),
            .in2(_gnd_net_),
            .in3(N__26194),
            .lcout(N_183),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPointerReset_RNO_1_LC_12_7_7.C_ON=1'b0;
    defparam sEEPointerReset_RNO_1_LC_12_7_7.SEQ_MODE=4'b0000;
    defparam sEEPointerReset_RNO_1_LC_12_7_7.LUT_INIT=16'b0100000000000000;
    LogicCell40 sEEPointerReset_RNO_1_LC_12_7_7 (
            .in0(N__26195),
            .in1(N__26099),
            .in2(N__49362),
            .in3(N__26048),
            .lcout(N_1624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_34_0_LC_12_8_0.C_ON=1'b0;
    defparam sDAC_mem_34_0_LC_12_8_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_0_LC_12_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_0_LC_12_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46141),
            .lcout(sDAC_mem_34Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52273),
            .ce(N__25982),
            .sr(N__51694));
    defparam sDAC_mem_34_1_LC_12_8_1.C_ON=1'b0;
    defparam sDAC_mem_34_1_LC_12_8_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_1_LC_12_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_1_LC_12_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50929),
            .lcout(sDAC_mem_34Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52273),
            .ce(N__25982),
            .sr(N__51694));
    defparam sDAC_mem_34_2_LC_12_8_2.C_ON=1'b0;
    defparam sDAC_mem_34_2_LC_12_8_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_2_LC_12_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_2_LC_12_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47246),
            .lcout(sDAC_mem_34Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52273),
            .ce(N__25982),
            .sr(N__51694));
    defparam sDAC_mem_34_3_LC_12_8_3.C_ON=1'b0;
    defparam sDAC_mem_34_3_LC_12_8_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_3_LC_12_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_3_LC_12_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46774),
            .lcout(sDAC_mem_34Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52273),
            .ce(N__25982),
            .sr(N__51694));
    defparam sDAC_mem_34_4_LC_12_8_4.C_ON=1'b0;
    defparam sDAC_mem_34_4_LC_12_8_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_4_LC_12_8_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_34_4_LC_12_8_4 (
            .in0(N__45373),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_34Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52273),
            .ce(N__25982),
            .sr(N__51694));
    defparam sDAC_mem_34_5_LC_12_8_5.C_ON=1'b0;
    defparam sDAC_mem_34_5_LC_12_8_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_5_LC_12_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_5_LC_12_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44841),
            .lcout(sDAC_mem_34Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52273),
            .ce(N__25982),
            .sr(N__51694));
    defparam sDAC_mem_34_6_LC_12_8_6.C_ON=1'b0;
    defparam sDAC_mem_34_6_LC_12_8_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_6_LC_12_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_6_LC_12_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50481),
            .lcout(sDAC_mem_34Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52273),
            .ce(N__25982),
            .sr(N__51694));
    defparam sDAC_mem_34_7_LC_12_8_7.C_ON=1'b0;
    defparam sDAC_mem_34_7_LC_12_8_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_7_LC_12_8_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_34_7_LC_12_8_7 (
            .in0(N__49910),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_34Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52273),
            .ce(N__25982),
            .sr(N__51694));
    defparam sDAC_mem_39_0_LC_12_9_0.C_ON=1'b0;
    defparam sDAC_mem_39_0_LC_12_9_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_0_LC_12_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_39_0_LC_12_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46142),
            .lcout(sDAC_mem_39Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52264),
            .ce(N__26240),
            .sr(N__51688));
    defparam sDAC_mem_39_1_LC_12_9_1.C_ON=1'b0;
    defparam sDAC_mem_39_1_LC_12_9_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_1_LC_12_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_39_1_LC_12_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50930),
            .lcout(sDAC_mem_39Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52264),
            .ce(N__26240),
            .sr(N__51688));
    defparam sDAC_mem_39_2_LC_12_9_2.C_ON=1'b0;
    defparam sDAC_mem_39_2_LC_12_9_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_2_LC_12_9_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_39_2_LC_12_9_2 (
            .in0(_gnd_net_),
            .in1(N__47247),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_39Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52264),
            .ce(N__26240),
            .sr(N__51688));
    defparam sDAC_mem_39_3_LC_12_9_3.C_ON=1'b0;
    defparam sDAC_mem_39_3_LC_12_9_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_3_LC_12_9_3.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_39_3_LC_12_9_3 (
            .in0(_gnd_net_),
            .in1(N__46775),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_39Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52264),
            .ce(N__26240),
            .sr(N__51688));
    defparam sDAC_mem_39_4_LC_12_9_4.C_ON=1'b0;
    defparam sDAC_mem_39_4_LC_12_9_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_4_LC_12_9_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_39_4_LC_12_9_4 (
            .in0(N__45374),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_39Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52264),
            .ce(N__26240),
            .sr(N__51688));
    defparam sDAC_mem_39_5_LC_12_9_5.C_ON=1'b0;
    defparam sDAC_mem_39_5_LC_12_9_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_5_LC_12_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_39_5_LC_12_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45078),
            .lcout(sDAC_mem_39Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52264),
            .ce(N__26240),
            .sr(N__51688));
    defparam sDAC_mem_39_6_LC_12_9_6.C_ON=1'b0;
    defparam sDAC_mem_39_6_LC_12_9_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_6_LC_12_9_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_39_6_LC_12_9_6 (
            .in0(N__50482),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_39Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52264),
            .ce(N__26240),
            .sr(N__51688));
    defparam sDAC_mem_39_7_LC_12_9_7.C_ON=1'b0;
    defparam sDAC_mem_39_7_LC_12_9_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_7_LC_12_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_39_7_LC_12_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49911),
            .lcout(sDAC_mem_39Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52264),
            .ce(N__26240),
            .sr(N__51688));
    defparam un1_spoff_cry_0_c_inv_LC_12_10_0.C_ON=1'b1;
    defparam un1_spoff_cry_0_c_inv_LC_12_10_0.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_0_c_inv_LC_12_10_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_0_c_inv_LC_12_10_0 (
            .in0(_gnd_net_),
            .in1(N__27892),
            .in2(N__26225),
            .in3(N__30188),
            .lcout(sCounter_i_0),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(un1_spoff_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_1_c_inv_LC_12_10_1.C_ON=1'b1;
    defparam un1_spoff_cry_1_c_inv_LC_12_10_1.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_1_c_inv_LC_12_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_1_c_inv_LC_12_10_1 (
            .in0(_gnd_net_),
            .in1(N__26210),
            .in2(N__27877),
            .in3(N__30070),
            .lcout(sCounter_i_1),
            .ltout(),
            .carryin(un1_spoff_cry_0),
            .carryout(un1_spoff_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_2_c_inv_LC_12_10_2.C_ON=1'b1;
    defparam un1_spoff_cry_2_c_inv_LC_12_10_2.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_2_c_inv_LC_12_10_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_2_c_inv_LC_12_10_2 (
            .in0(_gnd_net_),
            .in1(N__26339),
            .in2(N__27856),
            .in3(N__29945),
            .lcout(sCounter_i_2),
            .ltout(),
            .carryin(un1_spoff_cry_1),
            .carryout(un1_spoff_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_3_c_inv_LC_12_10_3.C_ON=1'b1;
    defparam un1_spoff_cry_3_c_inv_LC_12_10_3.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_3_c_inv_LC_12_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_3_c_inv_LC_12_10_3 (
            .in0(_gnd_net_),
            .in1(N__26327),
            .in2(N__28234),
            .in3(N__29818),
            .lcout(sCounter_i_3),
            .ltout(),
            .carryin(un1_spoff_cry_2),
            .carryout(un1_spoff_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_4_c_inv_LC_12_10_4.C_ON=1'b1;
    defparam un1_spoff_cry_4_c_inv_LC_12_10_4.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_4_c_inv_LC_12_10_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_4_c_inv_LC_12_10_4 (
            .in0(_gnd_net_),
            .in1(N__26315),
            .in2(N__28213),
            .in3(N__30955),
            .lcout(sCounter_i_4),
            .ltout(),
            .carryin(un1_spoff_cry_3),
            .carryout(un1_spoff_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_5_c_inv_LC_12_10_5.C_ON=1'b1;
    defparam un1_spoff_cry_5_c_inv_LC_12_10_5.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_5_c_inv_LC_12_10_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_5_c_inv_LC_12_10_5 (
            .in0(_gnd_net_),
            .in1(N__28189),
            .in2(N__26303),
            .in3(N__30838),
            .lcout(sCounter_i_5),
            .ltout(),
            .carryin(un1_spoff_cry_4),
            .carryout(un1_spoff_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_6_c_inv_LC_12_10_6.C_ON=1'b1;
    defparam un1_spoff_cry_6_c_inv_LC_12_10_6.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_6_c_inv_LC_12_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_6_c_inv_LC_12_10_6 (
            .in0(_gnd_net_),
            .in1(N__26288),
            .in2(N__28174),
            .in3(N__30727),
            .lcout(sCounter_i_6),
            .ltout(),
            .carryin(un1_spoff_cry_5),
            .carryout(un1_spoff_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_7_c_inv_LC_12_10_7.C_ON=1'b1;
    defparam un1_spoff_cry_7_c_inv_LC_12_10_7.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_7_c_inv_LC_12_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_7_c_inv_LC_12_10_7 (
            .in0(_gnd_net_),
            .in1(N__28150),
            .in2(N__26276),
            .in3(N__30627),
            .lcout(sCounter_i_7),
            .ltout(),
            .carryin(un1_spoff_cry_6),
            .carryout(un1_spoff_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_8_c_inv_LC_12_11_0.C_ON=1'b1;
    defparam un1_spoff_cry_8_c_inv_LC_12_11_0.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_8_c_inv_LC_12_11_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_8_c_inv_LC_12_11_0 (
            .in0(_gnd_net_),
            .in1(N__26780),
            .in2(N__28135),
            .in3(N__30517),
            .lcout(sCounter_i_8),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(un1_spoff_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_9_c_inv_LC_12_11_1.C_ON=1'b1;
    defparam un1_spoff_cry_9_c_inv_LC_12_11_1.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_9_c_inv_LC_12_11_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_9_c_inv_LC_12_11_1 (
            .in0(_gnd_net_),
            .in1(N__28111),
            .in2(N__26768),
            .in3(N__30407),
            .lcout(sCounter_i_9),
            .ltout(),
            .carryin(un1_spoff_cry_8),
            .carryout(un1_spoff_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_10_c_inv_LC_12_11_2.C_ON=1'b1;
    defparam un1_spoff_cry_10_c_inv_LC_12_11_2.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_10_c_inv_LC_12_11_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_10_c_inv_LC_12_11_2 (
            .in0(_gnd_net_),
            .in1(N__26261),
            .in2(N__28096),
            .in3(N__30290),
            .lcout(sCounter_i_10),
            .ltout(),
            .carryin(un1_spoff_cry_9),
            .carryout(un1_spoff_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_11_c_inv_LC_12_11_3.C_ON=1'b1;
    defparam un1_spoff_cry_11_c_inv_LC_12_11_3.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_11_c_inv_LC_12_11_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_11_c_inv_LC_12_11_3 (
            .in0(_gnd_net_),
            .in1(N__26516),
            .in2(N__28357),
            .in3(N__32990),
            .lcout(sCounter_i_11),
            .ltout(),
            .carryin(un1_spoff_cry_10),
            .carryout(un1_spoff_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_12_c_inv_LC_12_11_4.C_ON=1'b1;
    defparam un1_spoff_cry_12_c_inv_LC_12_11_4.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_12_c_inv_LC_12_11_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_12_c_inv_LC_12_11_4 (
            .in0(_gnd_net_),
            .in1(N__28336),
            .in2(N__26504),
            .in3(N__31700),
            .lcout(sCounter_i_12),
            .ltout(),
            .carryin(un1_spoff_cry_11),
            .carryout(un1_spoff_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_13_c_inv_LC_12_11_5.C_ON=1'b1;
    defparam un1_spoff_cry_13_c_inv_LC_12_11_5.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_13_c_inv_LC_12_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_13_c_inv_LC_12_11_5 (
            .in0(_gnd_net_),
            .in1(N__26492),
            .in2(N__28318),
            .in3(N__31610),
            .lcout(sCounter_i_13),
            .ltout(),
            .carryin(un1_spoff_cry_12),
            .carryout(un1_spoff_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_14_c_inv_LC_12_11_6.C_ON=1'b1;
    defparam un1_spoff_cry_14_c_inv_LC_12_11_6.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_14_c_inv_LC_12_11_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_spoff_cry_14_c_inv_LC_12_11_6 (
            .in0(N__31517),
            .in1(N__26480),
            .in2(N__28297),
            .in3(_gnd_net_),
            .lcout(sCounter_i_14),
            .ltout(),
            .carryin(un1_spoff_cry_13),
            .carryout(un1_spoff_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_15_c_inv_LC_12_11_7.C_ON=1'b1;
    defparam un1_spoff_cry_15_c_inv_LC_12_11_7.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_15_c_inv_LC_12_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_15_c_inv_LC_12_11_7 (
            .in0(_gnd_net_),
            .in1(N__28273),
            .in2(N__26795),
            .in3(N__31430),
            .lcout(sCounter_i_15),
            .ltout(),
            .carryin(un1_spoff_cry_14),
            .carryout(un1_spoff_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_16_c_inv_LC_12_12_0.C_ON=1'b1;
    defparam un1_spoff_cry_16_c_inv_LC_12_12_0.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_16_c_inv_LC_12_12_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_16_c_inv_LC_12_12_0 (
            .in0(_gnd_net_),
            .in1(N__26357),
            .in2(_gnd_net_),
            .in3(N__31338),
            .lcout(sCounter_i_16),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(un1_spoff_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_17_c_inv_LC_12_12_1.C_ON=1'b1;
    defparam un1_spoff_cry_17_c_inv_LC_12_12_1.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_17_c_inv_LC_12_12_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_spoff_cry_17_c_inv_LC_12_12_1 (
            .in0(N__31262),
            .in1(N__26351),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sCounter_i_17),
            .ltout(),
            .carryin(un1_spoff_cry_16),
            .carryout(un1_spoff_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_18_c_inv_LC_12_12_2.C_ON=1'b1;
    defparam un1_spoff_cry_18_c_inv_LC_12_12_2.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_18_c_inv_LC_12_12_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_18_c_inv_LC_12_12_2 (
            .in0(_gnd_net_),
            .in1(N__26345),
            .in2(_gnd_net_),
            .in3(N__31148),
            .lcout(sCounter_i_18),
            .ltout(),
            .carryin(un1_spoff_cry_17),
            .carryout(un1_spoff_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_19_c_inv_LC_12_12_3.C_ON=1'b1;
    defparam un1_spoff_cry_19_c_inv_LC_12_12_3.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_19_c_inv_LC_12_12_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_spoff_cry_19_c_inv_LC_12_12_3 (
            .in0(N__33225),
            .in1(N__26456),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sCounter_i_19),
            .ltout(),
            .carryin(un1_spoff_cry_18),
            .carryout(un1_spoff_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_20_c_inv_LC_12_12_4.C_ON=1'b1;
    defparam un1_spoff_cry_20_c_inv_LC_12_12_4.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_20_c_inv_LC_12_12_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_20_c_inv_LC_12_12_4 (
            .in0(_gnd_net_),
            .in1(N__26450),
            .in2(_gnd_net_),
            .in3(N__33332),
            .lcout(sCounter_i_20),
            .ltout(),
            .carryin(un1_spoff_cry_19),
            .carryout(un1_spoff_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_21_c_inv_LC_12_12_5.C_ON=1'b1;
    defparam un1_spoff_cry_21_c_inv_LC_12_12_5.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_21_c_inv_LC_12_12_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_spoff_cry_21_c_inv_LC_12_12_5 (
            .in0(N__33116),
            .in1(N__26444),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sCounter_i_21),
            .ltout(),
            .carryin(un1_spoff_cry_20),
            .carryout(un1_spoff_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_22_c_inv_LC_12_12_6.C_ON=1'b1;
    defparam un1_spoff_cry_22_c_inv_LC_12_12_6.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_22_c_inv_LC_12_12_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_spoff_cry_22_c_inv_LC_12_12_6 (
            .in0(N__32018),
            .in1(N__26438),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sCounter_i_22),
            .ltout(),
            .carryin(un1_spoff_cry_21),
            .carryout(un1_spoff_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_23_c_inv_LC_12_12_7.C_ON=1'b1;
    defparam un1_spoff_cry_23_c_inv_LC_12_12_7.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_23_c_inv_LC_12_12_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_23_c_inv_LC_12_12_7 (
            .in0(_gnd_net_),
            .in1(N__26432),
            .in2(_gnd_net_),
            .in3(N__31883),
            .lcout(sCounter_i_23),
            .ltout(),
            .carryin(un1_spoff_cry_22),
            .carryout(un1_spoff_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam poff_obuf_RNO_LC_12_13_0.C_ON=1'b0;
    defparam poff_obuf_RNO_LC_12_13_0.SEQ_MODE=4'b0000;
    defparam poff_obuf_RNO_LC_12_13_0.LUT_INIT=16'b0101010111111111;
    LogicCell40 poff_obuf_RNO_LC_12_13_0 (
            .in0(N__31817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26426),
            .lcout(N_1683_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_LC_12_13_1.C_ON=1'b0;
    defparam sbuttonModeStatus_LC_12_13_1.SEQ_MODE=4'b1000;
    defparam sbuttonModeStatus_LC_12_13_1.LUT_INIT=16'b0111100011110000;
    LogicCell40 sbuttonModeStatus_LC_12_13_1 (
            .in0(N__32921),
            .in1(N__26363),
            .in2(N__26389),
            .in3(N__33803),
            .lcout(sbuttonModeStatusZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48468),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_1_LC_12_13_7.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_1_LC_12_13_7.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_1_LC_12_13_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_1_LC_12_13_7 (
            .in0(N__45752),
            .in1(N__45776),
            .in2(N__35108),
            .in3(N__26372),
            .lcout(sbuttonModeStatus_0_sqmuxa_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEACQ_0_LC_12_14_0.C_ON=1'b0;
    defparam sEEACQ_0_LC_12_14_0.SEQ_MODE=4'b1010;
    defparam sEEACQ_0_LC_12_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_0_LC_12_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46381),
            .lcout(sEEACQZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52274),
            .ce(N__26471),
            .sr(N__51654));
    defparam sEEACQ_1_LC_12_14_1.C_ON=1'b0;
    defparam sEEACQ_1_LC_12_14_1.SEQ_MODE=4'b1010;
    defparam sEEACQ_1_LC_12_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_1_LC_12_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50877),
            .lcout(sEEACQZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52274),
            .ce(N__26471),
            .sr(N__51654));
    defparam sEEACQ_2_LC_12_14_2.C_ON=1'b0;
    defparam sEEACQ_2_LC_12_14_2.SEQ_MODE=4'b1010;
    defparam sEEACQ_2_LC_12_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_2_LC_12_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47458),
            .lcout(sEEACQZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52274),
            .ce(N__26471),
            .sr(N__51654));
    defparam sEEACQ_3_LC_12_14_3.C_ON=1'b0;
    defparam sEEACQ_3_LC_12_14_3.SEQ_MODE=4'b1011;
    defparam sEEACQ_3_LC_12_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_3_LC_12_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46915),
            .lcout(sEEACQZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52274),
            .ce(N__26471),
            .sr(N__51654));
    defparam sEEACQ_4_LC_12_14_4.C_ON=1'b0;
    defparam sEEACQ_4_LC_12_14_4.SEQ_MODE=4'b1010;
    defparam sEEACQ_4_LC_12_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_4_LC_12_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45568),
            .lcout(sEEACQZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52274),
            .ce(N__26471),
            .sr(N__51654));
    defparam sEEACQ_5_LC_12_14_5.C_ON=1'b0;
    defparam sEEACQ_5_LC_12_14_5.SEQ_MODE=4'b1010;
    defparam sEEACQ_5_LC_12_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_5_LC_12_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45080),
            .lcout(sEEACQZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52274),
            .ce(N__26471),
            .sr(N__51654));
    defparam sEEACQ_6_LC_12_14_6.C_ON=1'b0;
    defparam sEEACQ_6_LC_12_14_6.SEQ_MODE=4'b1011;
    defparam sEEACQ_6_LC_12_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_6_LC_12_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50531),
            .lcout(sEEACQZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52274),
            .ce(N__26471),
            .sr(N__51654));
    defparam sEEACQ_7_LC_12_14_7.C_ON=1'b0;
    defparam sEEACQ_7_LC_12_14_7.SEQ_MODE=4'b1011;
    defparam sEEACQ_7_LC_12_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_7_LC_12_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50050),
            .lcout(sEEACQZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52274),
            .ce(N__26471),
            .sr(N__51654));
    defparam sEEACQ_10_LC_12_15_0.C_ON=1'b0;
    defparam sEEACQ_10_LC_12_15_0.SEQ_MODE=4'b1010;
    defparam sEEACQ_10_LC_12_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_10_LC_12_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47460),
            .lcout(sEEACQZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52286),
            .ce(N__26525),
            .sr(N__51651));
    defparam sEEACQ_11_LC_12_15_1.C_ON=1'b0;
    defparam sEEACQ_11_LC_12_15_1.SEQ_MODE=4'b1010;
    defparam sEEACQ_11_LC_12_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_11_LC_12_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46925),
            .lcout(sEEACQZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52286),
            .ce(N__26525),
            .sr(N__51651));
    defparam sEEACQ_12_LC_12_15_2.C_ON=1'b0;
    defparam sEEACQ_12_LC_12_15_2.SEQ_MODE=4'b1011;
    defparam sEEACQ_12_LC_12_15_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEACQ_12_LC_12_15_2 (
            .in0(N__45569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEACQZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52286),
            .ce(N__26525),
            .sr(N__51651));
    defparam sEEACQ_13_LC_12_15_3.C_ON=1'b0;
    defparam sEEACQ_13_LC_12_15_3.SEQ_MODE=4'b1011;
    defparam sEEACQ_13_LC_12_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_13_LC_12_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45057),
            .lcout(sEEACQZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52286),
            .ce(N__26525),
            .sr(N__51651));
    defparam sEEACQ_14_LC_12_15_4.C_ON=1'b0;
    defparam sEEACQ_14_LC_12_15_4.SEQ_MODE=4'b1010;
    defparam sEEACQ_14_LC_12_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_14_LC_12_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50544),
            .lcout(sEEACQZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52286),
            .ce(N__26525),
            .sr(N__51651));
    defparam sEEACQ_15_LC_12_15_5.C_ON=1'b0;
    defparam sEEACQ_15_LC_12_15_5.SEQ_MODE=4'b1010;
    defparam sEEACQ_15_LC_12_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_15_LC_12_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50016),
            .lcout(sEEACQZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52286),
            .ce(N__26525),
            .sr(N__51651));
    defparam sEEACQ_8_LC_12_15_6.C_ON=1'b0;
    defparam sEEACQ_8_LC_12_15_6.SEQ_MODE=4'b1010;
    defparam sEEACQ_8_LC_12_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_8_LC_12_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46380),
            .lcout(sEEACQZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52286),
            .ce(N__26525),
            .sr(N__51651));
    defparam sEEACQ_9_LC_12_15_7.C_ON=1'b0;
    defparam sEEACQ_9_LC_12_15_7.SEQ_MODE=4'b1011;
    defparam sEEACQ_9_LC_12_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_9_LC_12_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51018),
            .lcout(sEEACQZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52286),
            .ce(N__26525),
            .sr(N__51651));
    defparam sEEPoff_11_LC_12_16_0.C_ON=1'b0;
    defparam sEEPoff_11_LC_12_16_0.SEQ_MODE=4'b1010;
    defparam sEEPoff_11_LC_12_16_0.LUT_INIT=16'b1100110011001100;
    LogicCell40 sEEPoff_11_LC_12_16_0 (
            .in0(_gnd_net_),
            .in1(N__46763),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPoffZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52298),
            .ce(N__26756),
            .sr(N__51648));
    defparam sEEPoff_12_LC_12_16_1.C_ON=1'b0;
    defparam sEEPoff_12_LC_12_16_1.SEQ_MODE=4'b1010;
    defparam sEEPoff_12_LC_12_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_12_LC_12_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45570),
            .lcout(sEEPoffZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52298),
            .ce(N__26756),
            .sr(N__51648));
    defparam sEEPoff_13_LC_12_16_2.C_ON=1'b0;
    defparam sEEPoff_13_LC_12_16_2.SEQ_MODE=4'b1010;
    defparam sEEPoff_13_LC_12_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_13_LC_12_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45056),
            .lcout(sEEPoffZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52298),
            .ce(N__26756),
            .sr(N__51648));
    defparam sEEPoff_14_LC_12_16_3.C_ON=1'b0;
    defparam sEEPoff_14_LC_12_16_3.SEQ_MODE=4'b1010;
    defparam sEEPoff_14_LC_12_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_14_LC_12_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50545),
            .lcout(sEEPoffZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52298),
            .ce(N__26756),
            .sr(N__51648));
    defparam sEEPoff_15_LC_12_16_4.C_ON=1'b0;
    defparam sEEPoff_15_LC_12_16_4.SEQ_MODE=4'b1010;
    defparam sEEPoff_15_LC_12_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_15_LC_12_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50058),
            .lcout(sEEPoffZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52298),
            .ce(N__26756),
            .sr(N__51648));
    defparam sEEPoff_8_LC_12_16_5.C_ON=1'b0;
    defparam sEEPoff_8_LC_12_16_5.SEQ_MODE=4'b1010;
    defparam sEEPoff_8_LC_12_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_8_LC_12_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46379),
            .lcout(sEEPoffZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52298),
            .ce(N__26756),
            .sr(N__51648));
    defparam sEEPoff_9_LC_12_16_6.C_ON=1'b0;
    defparam sEEPoff_9_LC_12_16_6.SEQ_MODE=4'b1010;
    defparam sEEPoff_9_LC_12_16_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPoff_9_LC_12_16_6 (
            .in0(N__51062),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPoffZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52298),
            .ce(N__26756),
            .sr(N__51648));
    defparam un4_sacqtime_cry_23_c_RNI2CQM_LC_12_17_3.C_ON=1'b0;
    defparam un4_sacqtime_cry_23_c_RNI2CQM_LC_12_17_3.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_23_c_RNI2CQM_LC_12_17_3.LUT_INIT=16'b1111010011110000;
    LogicCell40 un4_sacqtime_cry_23_c_RNI2CQM_LC_12_17_3 (
            .in0(N__49462),
            .in1(N__43315),
            .in2(N__39387),
            .in3(N__43438),
            .lcout(un4_sacqtime_cry_23_c_RNI2CQMZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_1_5_LC_12_18_0.C_ON=1'b0;
    defparam RAM_DATA_1_5_LC_12_18_0.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_5_LC_12_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_5_LC_12_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26720),
            .lcout(RAM_DATA_1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52321),
            .ce(N__51872),
            .sr(N__51644));
    defparam RAM_DATA_1_1_LC_12_18_1.C_ON=1'b0;
    defparam RAM_DATA_1_1_LC_12_18_1.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_1_LC_12_18_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 RAM_DATA_1_1_LC_12_18_1 (
            .in0(N__26678),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RAM_DATA_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52321),
            .ce(N__51872),
            .sr(N__51644));
    defparam RAM_DATA_1_10_LC_12_18_2.C_ON=1'b0;
    defparam RAM_DATA_1_10_LC_12_18_2.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_10_LC_12_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_10_LC_12_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26645),
            .lcout(RAM_DATA_1Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52321),
            .ce(N__51872),
            .sr(N__51644));
    defparam RAM_DATA_1_11_LC_12_18_3.C_ON=1'b0;
    defparam RAM_DATA_1_11_LC_12_18_3.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_11_LC_12_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_11_LC_12_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26609),
            .lcout(RAM_DATA_1Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52321),
            .ce(N__51872),
            .sr(N__51644));
    defparam RAM_DATA_1_13_LC_12_18_5.C_ON=1'b0;
    defparam RAM_DATA_1_13_LC_12_18_5.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_13_LC_12_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_13_LC_12_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26573),
            .lcout(RAM_DATA_1Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52321),
            .ce(N__51872),
            .sr(N__51644));
    defparam RAM_DATA_1_14_LC_12_18_6.C_ON=1'b0;
    defparam RAM_DATA_1_14_LC_12_18_6.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_14_LC_12_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_14_LC_12_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26960),
            .lcout(RAM_DATA_1Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52321),
            .ce(N__51872),
            .sr(N__51644));
    defparam RAM_DATA_1_2_LC_12_18_7.C_ON=1'b0;
    defparam RAM_DATA_1_2_LC_12_18_7.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_2_LC_12_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_2_LC_12_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26912),
            .lcout(RAM_DATA_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52321),
            .ce(N__51872),
            .sr(N__51644));
    defparam RAM_DATA_1_6_LC_12_20_4.C_ON=1'b0;
    defparam RAM_DATA_1_6_LC_12_20_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_6_LC_12_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_6_LC_12_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26879),
            .lcout(RAM_DATA_1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52339),
            .ce(N__51889),
            .sr(N__51642));
    defparam RAM_DATA_1_0_LC_12_20_6.C_ON=1'b0;
    defparam RAM_DATA_1_0_LC_12_20_6.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_0_LC_12_20_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_0_LC_12_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26840),
            .lcout(RAM_DATA_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52339),
            .ce(N__51889),
            .sr(N__51642));
    defparam sDAC_mem_40_0_LC_13_3_0.C_ON=1'b0;
    defparam sDAC_mem_40_0_LC_13_3_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_0_LC_13_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_0_LC_13_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46144),
            .lcout(sDAC_mem_40Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52323),
            .ce(N__27125),
            .sr(N__51768));
    defparam sDAC_mem_40_1_LC_13_3_1.C_ON=1'b0;
    defparam sDAC_mem_40_1_LC_13_3_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_1_LC_13_3_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_1_LC_13_3_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51075),
            .lcout(sDAC_mem_40Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52323),
            .ce(N__27125),
            .sr(N__51768));
    defparam sDAC_mem_40_2_LC_13_3_2.C_ON=1'b0;
    defparam sDAC_mem_40_2_LC_13_3_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_2_LC_13_3_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_2_LC_13_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47346),
            .lcout(sDAC_mem_40Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52323),
            .ce(N__27125),
            .sr(N__51768));
    defparam sDAC_mem_40_3_LC_13_3_3.C_ON=1'b0;
    defparam sDAC_mem_40_3_LC_13_3_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_3_LC_13_3_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_3_LC_13_3_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46793),
            .lcout(sDAC_mem_40Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52323),
            .ce(N__27125),
            .sr(N__51768));
    defparam sDAC_mem_40_4_LC_13_3_4.C_ON=1'b0;
    defparam sDAC_mem_40_4_LC_13_3_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_4_LC_13_3_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_4_LC_13_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45529),
            .lcout(sDAC_mem_40Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52323),
            .ce(N__27125),
            .sr(N__51768));
    defparam sDAC_mem_40_5_LC_13_3_5.C_ON=1'b0;
    defparam sDAC_mem_40_5_LC_13_3_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_5_LC_13_3_5.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_40_5_LC_13_3_5 (
            .in0(_gnd_net_),
            .in1(N__45053),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_40Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52323),
            .ce(N__27125),
            .sr(N__51768));
    defparam sDAC_mem_40_6_LC_13_3_6.C_ON=1'b0;
    defparam sDAC_mem_40_6_LC_13_3_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_6_LC_13_3_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_6_LC_13_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50420),
            .lcout(sDAC_mem_40Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52323),
            .ce(N__27125),
            .sr(N__51768));
    defparam sDAC_mem_40_7_LC_13_3_7.C_ON=1'b0;
    defparam sDAC_mem_40_7_LC_13_3_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_7_LC_13_3_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_40_7_LC_13_3_7 (
            .in0(N__49995),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_40Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52323),
            .ce(N__27125),
            .sr(N__51768));
    defparam sAddress_RNI9IH12_0_2_LC_13_4_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_0_2_LC_13_4_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_0_2_LC_13_4_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 sAddress_RNI9IH12_0_2_LC_13_4_0 (
            .in0(N__40673),
            .in1(N__27020),
            .in2(N__41010),
            .in3(N__40809),
            .lcout(sDAC_mem_40_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_3_2_LC_13_4_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_3_2_LC_13_4_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_3_2_LC_13_4_2.LUT_INIT=16'b0100000000000000;
    LogicCell40 sAddress_RNI9IH12_3_2_LC_13_4_2 (
            .in0(N__40674),
            .in1(N__27022),
            .in2(N__41011),
            .in3(N__40810),
            .lcout(sDAC_mem_36_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_4_2_LC_13_4_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_4_2_LC_13_4_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_4_2_LC_13_4_3.LUT_INIT=16'b0000100000000000;
    LogicCell40 sAddress_RNI9IH12_4_2_LC_13_4_3 (
            .in0(N__27021),
            .in1(N__40811),
            .in2(N__41012),
            .in3(N__40675),
            .lcout(sDAC_mem_8_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_rpi_ibuf_RNIRGF52_0_LC_13_4_5.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNIRGF52_0_LC_13_4_5.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNIRGF52_0_LC_13_4_5.LUT_INIT=16'b0100000000000000;
    LogicCell40 reset_rpi_ibuf_RNIRGF52_0_LC_13_4_5 (
            .in0(N__27110),
            .in1(N__27062),
            .in2(N__49260),
            .in3(N__33769),
            .lcout(sEEDAC_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_2_2_LC_13_4_6.C_ON=1'b0;
    defparam sAddress_RNI9IH12_2_2_LC_13_4_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_2_2_LC_13_4_6.LUT_INIT=16'b0000101000000000;
    LogicCell40 sAddress_RNI9IH12_2_2_LC_13_4_6 (
            .in0(N__40025),
            .in1(_gnd_net_),
            .in2(N__40676),
            .in3(N__27019),
            .lcout(sDAC_mem_20_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_1_LC_13_4_7.C_ON=1'b0;
    defparam sAddress_RNI9IH12_1_LC_13_4_7.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_1_LC_13_4_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 sAddress_RNI9IH12_1_LC_13_4_7 (
            .in0(_gnd_net_),
            .in1(N__26984),
            .in2(_gnd_net_),
            .in3(N__40024),
            .lcout(sDAC_mem_21_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_6_LC_13_5_0.C_ON=1'b0;
    defparam sDAC_data_RNO_22_6_LC_13_5_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_6_LC_13_5_0.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_22_6_LC_13_5_0 (
            .in0(N__38556),
            .in1(N__28478),
            .in2(N__38207),
            .in3(N__28679),
            .lcout(),
            .ltout(sDAC_data_2_32_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_6_LC_13_5_1.C_ON=1'b0;
    defparam sDAC_data_RNO_10_6_LC_13_5_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_6_LC_13_5_1.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_10_6_LC_13_5_1 (
            .in0(N__38301),
            .in1(N__32354),
            .in2(N__27206),
            .in3(N__34406),
            .lcout(sDAC_data_RNO_10Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_6_LC_13_5_2.C_ON=1'b0;
    defparam sDAC_data_RNO_6_6_LC_13_5_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_6_LC_13_5_2.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_6_6_LC_13_5_2 (
            .in0(N__38557),
            .in1(N__27203),
            .in2(N__38208),
            .in3(N__36674),
            .lcout(),
            .ltout(sDAC_data_2_14_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_6_LC_13_5_3.C_ON=1'b0;
    defparam sDAC_data_RNO_1_6_LC_13_5_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_6_LC_13_5_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_1_6_LC_13_5_3 (
            .in0(N__38302),
            .in1(N__28718),
            .in2(N__27197),
            .in3(N__39641),
            .lcout(sDAC_data_RNO_1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_6_LC_13_5_4.C_ON=1'b0;
    defparam sDAC_data_RNO_3_6_LC_13_5_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_6_LC_13_5_4.LUT_INIT=16'b0010010101110101;
    LogicCell40 sDAC_data_RNO_3_6_LC_13_5_4 (
            .in0(N__37355),
            .in1(N__37829),
            .in2(N__37472),
            .in3(N__27194),
            .lcout(),
            .ltout(sDAC_data_2_41_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_6_LC_13_5_5.C_ON=1'b0;
    defparam sDAC_data_RNO_0_6_LC_13_5_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_6_LC_13_5_5.LUT_INIT=16'b0101111000001110;
    LogicCell40 sDAC_data_RNO_0_6_LC_13_5_5 (
            .in0(N__37461),
            .in1(N__27188),
            .in2(N__27182),
            .in3(N__27179),
            .lcout(),
            .ltout(sDAC_data_2_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_6_LC_13_5_6.C_ON=1'b0;
    defparam sDAC_data_6_LC_13_5_6.SEQ_MODE=4'b1010;
    defparam sDAC_data_6_LC_13_5_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 sDAC_data_6_LC_13_5_6 (
            .in0(N__32099),
            .in1(_gnd_net_),
            .in2(N__27173),
            .in3(N__37636),
            .lcout(sDAC_dataZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48445),
            .ce(N__43956),
            .sr(N__51743));
    defparam sDAC_mem_3_5_LC_13_6_0.C_ON=1'b0;
    defparam sDAC_mem_3_5_LC_13_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_5_LC_13_6_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_3_5_LC_13_6_0 (
            .in0(N__45001),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_3Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52287),
            .ce(N__44243),
            .sr(N__51728));
    defparam sDAC_data_RNO_27_8_LC_13_6_1.C_ON=1'b0;
    defparam sDAC_data_RNO_27_8_LC_13_6_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_8_LC_13_6_1.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_27_8_LC_13_6_1 (
            .in0(N__42570),
            .in1(N__27161),
            .in2(N__42204),
            .in3(N__27149),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_8_LC_13_6_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_8_LC_13_6_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_8_LC_13_6_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_8_LC_13_6_2 (
            .in0(N__42242),
            .in1(N__27143),
            .in2(N__27134),
            .in3(N__27131),
            .lcout(sDAC_data_RNO_15Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_8_LC_13_6_3.C_ON=1'b0;
    defparam sDAC_data_RNO_17_8_LC_13_6_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_8_LC_13_6_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_8_LC_13_6_3 (
            .in0(N__42569),
            .in1(N__27290),
            .in2(_gnd_net_),
            .in3(N__27278),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_8_LC_13_6_4.C_ON=1'b0;
    defparam sDAC_data_RNO_8_8_LC_13_6_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_8_LC_13_6_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_8_8_LC_13_6_4 (
            .in0(_gnd_net_),
            .in1(N__42072),
            .in2(N__27266),
            .in3(N__27263),
            .lcout(sDAC_data_RNO_8Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_8_LC_13_6_5.C_ON=1'b0;
    defparam sDAC_data_RNO_16_8_LC_13_6_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_8_LC_13_6_5.LUT_INIT=16'b0001110000011111;
    LogicCell40 sDAC_data_RNO_16_8_LC_13_6_5 (
            .in0(N__27254),
            .in1(N__42243),
            .in2(N__42580),
            .in3(N__27245),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_8_LC_13_6_6.C_ON=1'b0;
    defparam sDAC_data_RNO_7_8_LC_13_6_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_8_LC_13_6_6.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_7_8_LC_13_6_6 (
            .in0(N__36788),
            .in1(N__42073),
            .in2(N__27236),
            .in3(N__39857),
            .lcout(),
            .ltout(sDAC_data_RNO_7Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_8_LC_13_6_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_8_LC_13_6_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_8_LC_13_6_7.LUT_INIT=16'b0111010101100100;
    LogicCell40 sDAC_data_RNO_2_8_LC_13_6_7 (
            .in0(N__28655),
            .in1(N__38303),
            .in2(N__27233),
            .in3(N__27230),
            .lcout(sDAC_data_RNO_2Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_8_LC_13_7_0.C_ON=1'b0;
    defparam sDAC_data_RNO_6_8_LC_13_7_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_8_LC_13_7_0.LUT_INIT=16'b0101010100100111;
    LogicCell40 sDAC_data_RNO_6_8_LC_13_7_0 (
            .in0(N__38476),
            .in1(N__27224),
            .in2(N__36860),
            .in3(N__38288),
            .lcout(),
            .ltout(sDAC_data_2_14_ns_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_8_LC_13_7_1.C_ON=1'b0;
    defparam sDAC_data_RNO_1_8_LC_13_7_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_8_LC_13_7_1.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_1_8_LC_13_7_1 (
            .in0(N__38289),
            .in1(N__32498),
            .in2(N__27218),
            .in3(N__32549),
            .lcout(),
            .ltout(sDAC_data_RNO_1Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_8_LC_13_7_2.C_ON=1'b0;
    defparam sDAC_data_RNO_0_8_LC_13_7_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_8_LC_13_7_2.LUT_INIT=16'b0101000011101110;
    LogicCell40 sDAC_data_RNO_0_8_LC_13_7_2 (
            .in0(N__37457),
            .in1(N__27215),
            .in2(N__27209),
            .in3(N__27377),
            .lcout(),
            .ltout(sDAC_data_2_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_8_LC_13_7_3.C_ON=1'b0;
    defparam sDAC_data_8_LC_13_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_data_8_LC_13_7_3.LUT_INIT=16'b1110010011100100;
    LogicCell40 sDAC_data_8_LC_13_7_3 (
            .in0(N__37627),
            .in1(N__32087),
            .in2(N__27386),
            .in3(_gnd_net_),
            .lcout(sDAC_dataZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48450),
            .ce(N__43953),
            .sr(N__51716));
    defparam sDAC_data_RNO_22_8_LC_13_7_4.C_ON=1'b0;
    defparam sDAC_data_RNO_22_8_LC_13_7_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_8_LC_13_7_4.LUT_INIT=16'b0001110000011111;
    LogicCell40 sDAC_data_RNO_22_8_LC_13_7_4 (
            .in0(N__28565),
            .in1(N__38286),
            .in2(N__38510),
            .in3(N__28814),
            .lcout(),
            .ltout(sDAC_data_2_32_ns_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_8_LC_13_7_5.C_ON=1'b0;
    defparam sDAC_data_RNO_10_8_LC_13_7_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_8_LC_13_7_5.LUT_INIT=16'b1000111110000101;
    LogicCell40 sDAC_data_RNO_10_8_LC_13_7_5 (
            .in0(N__38287),
            .in1(N__32231),
            .in2(N__27383),
            .in3(N__33581),
            .lcout(),
            .ltout(sDAC_data_RNO_10Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_8_LC_13_7_6.C_ON=1'b0;
    defparam sDAC_data_RNO_3_8_LC_13_7_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_8_LC_13_7_6.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_3_8_LC_13_7_6 (
            .in0(N__37456),
            .in1(N__37351),
            .in2(N__27380),
            .in3(N__27521),
            .lcout(sDAC_data_2_41_ns_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_3_1_LC_13_8_0.C_ON=1'b0;
    defparam sDAC_mem_3_1_LC_13_8_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_1_LC_13_8_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_3_1_LC_13_8_0 (
            .in0(N__50928),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_3Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52265),
            .ce(N__44224),
            .sr(N__51705));
    defparam sDAC_data_RNO_27_4_LC_13_8_1.C_ON=1'b0;
    defparam sDAC_data_RNO_27_4_LC_13_8_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_4_LC_13_8_1.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_27_4_LC_13_8_1 (
            .in0(N__42545),
            .in1(N__27371),
            .in2(N__42246),
            .in3(N__27365),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_4_LC_13_8_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_4_LC_13_8_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_4_LC_13_8_2.LUT_INIT=16'b1010110000001111;
    LogicCell40 sDAC_data_RNO_15_4_LC_13_8_2 (
            .in0(N__27356),
            .in1(N__27350),
            .in2(N__27335),
            .in3(N__42197),
            .lcout(sDAC_data_RNO_15Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_4_LC_13_8_3.C_ON=1'b0;
    defparam sDAC_data_RNO_17_4_LC_13_8_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_4_LC_13_8_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 sDAC_data_RNO_17_4_LC_13_8_3 (
            .in0(N__27332),
            .in1(_gnd_net_),
            .in2(N__42574),
            .in3(N__27320),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_4_LC_13_8_4.C_ON=1'b0;
    defparam sDAC_data_RNO_8_4_LC_13_8_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_4_LC_13_8_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_8_4_LC_13_8_4 (
            .in0(_gnd_net_),
            .in1(N__42198),
            .in2(N__27308),
            .in3(N__27305),
            .lcout(sDAC_data_RNO_8Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_4_LC_13_8_5.C_ON=1'b0;
    defparam sDAC_data_RNO_16_4_LC_13_8_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_4_LC_13_8_5.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_16_4_LC_13_8_5 (
            .in0(N__42549),
            .in1(N__27485),
            .in2(N__42247),
            .in3(N__27476),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_4_LC_13_8_6.C_ON=1'b0;
    defparam sDAC_data_RNO_7_4_LC_13_8_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_4_LC_13_8_6.LUT_INIT=16'b1010110000001111;
    LogicCell40 sDAC_data_RNO_7_4_LC_13_8_6 (
            .in0(N__36833),
            .in1(N__39896),
            .in2(N__27464),
            .in3(N__42202),
            .lcout(),
            .ltout(sDAC_data_RNO_7Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_4_LC_13_8_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_4_LC_13_8_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_4_LC_13_8_7.LUT_INIT=16'b0111010101100100;
    LogicCell40 sDAC_data_RNO_2_4_LC_13_8_7 (
            .in0(N__27419),
            .in1(N__38111),
            .in2(N__27461),
            .in3(N__27458),
            .lcout(sDAC_data_RNO_2Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_19_3_LC_13_9_0.C_ON=1'b0;
    defparam sDAC_data_RNO_19_3_LC_13_9_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_3_LC_13_9_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_19_3_LC_13_9_0 (
            .in0(N__27452),
            .in1(N__42075),
            .in2(_gnd_net_),
            .in3(N__27443),
            .lcout(sDAC_data_RNO_19Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_3_LC_13_9_1.C_ON=1'b0;
    defparam sDAC_data_RNO_18_3_LC_13_9_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_3_LC_13_9_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_3_LC_13_9_1 (
            .in0(N__42076),
            .in1(N__45668),
            .in2(_gnd_net_),
            .in3(N__27584),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_3_LC_13_9_2.C_ON=1'b0;
    defparam sDAC_data_RNO_9_3_LC_13_9_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_3_LC_13_9_2.LUT_INIT=16'b0001010110011101;
    LogicCell40 sDAC_data_RNO_9_3_LC_13_9_2 (
            .in0(N__38489),
            .in1(N__38290),
            .in2(N__27431),
            .in3(N__27428),
            .lcout(sDAC_data_2_24_ns_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_4_LC_13_9_3.C_ON=1'b0;
    defparam sDAC_data_RNO_18_4_LC_13_9_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_4_LC_13_9_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_4_LC_13_9_3 (
            .in0(N__42080),
            .in1(N__45653),
            .in2(_gnd_net_),
            .in3(N__27578),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_4_LC_13_9_4.C_ON=1'b0;
    defparam sDAC_data_RNO_9_4_LC_13_9_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_4_LC_13_9_4.LUT_INIT=16'b0001010110011101;
    LogicCell40 sDAC_data_RNO_9_4_LC_13_9_4 (
            .in0(N__38490),
            .in1(N__38291),
            .in2(N__27422),
            .in3(N__27392),
            .lcout(sDAC_data_2_24_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_19_4_LC_13_9_5.C_ON=1'b0;
    defparam sDAC_data_RNO_19_4_LC_13_9_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_4_LC_13_9_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 sDAC_data_RNO_19_4_LC_13_9_5 (
            .in0(N__27413),
            .in1(_gnd_net_),
            .in2(N__42205),
            .in3(N__27404),
            .lcout(sDAC_data_RNO_19Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_12_0_LC_13_9_6.C_ON=1'b0;
    defparam sDAC_mem_12_0_LC_13_9_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_0_LC_13_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_0_LC_13_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46143),
            .lcout(sDAC_mem_12Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52252),
            .ce(N__36952),
            .sr(N__51698));
    defparam sDAC_mem_12_1_LC_13_9_7.C_ON=1'b0;
    defparam sDAC_mem_12_1_LC_13_9_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_1_LC_13_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_1_LC_13_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50931),
            .lcout(sDAC_mem_12Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52252),
            .ce(N__36952),
            .sr(N__51698));
    defparam sDAC_data_RNO_24_8_LC_13_10_0.C_ON=1'b0;
    defparam sDAC_data_RNO_24_8_LC_13_10_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_8_LC_13_10_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_8_LC_13_10_0 (
            .in0(N__41990),
            .in1(N__27572),
            .in2(_gnd_net_),
            .in3(N__27560),
            .lcout(sDAC_data_RNO_24Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_8_LC_13_10_1.C_ON=1'b0;
    defparam sDAC_data_RNO_23_8_LC_13_10_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_8_LC_13_10_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_8_LC_13_10_1 (
            .in0(N__42014),
            .in1(N__27545),
            .in2(_gnd_net_),
            .in3(N__27512),
            .lcout(),
            .ltout(sDAC_data_RNO_23Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_8_LC_13_10_2.C_ON=1'b0;
    defparam sDAC_data_RNO_11_8_LC_13_10_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_8_LC_13_10_2.LUT_INIT=16'b1010000011011101;
    LogicCell40 sDAC_data_RNO_11_8_LC_13_10_2 (
            .in0(N__38300),
            .in1(N__27530),
            .in2(N__27524),
            .in3(N__27590),
            .lcout(sDAC_data_RNO_11Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_28_5_LC_13_10_3.C_ON=1'b0;
    defparam sDAC_mem_28_5_LC_13_10_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_5_LC_13_10_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_28_5_LC_13_10_3 (
            .in0(N__45077),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_28Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52242),
            .ce(N__37796),
            .sr(N__51690));
    defparam sDAC_data_RNO_30_9_LC_13_10_4.C_ON=1'b0;
    defparam sDAC_data_RNO_30_9_LC_13_10_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_9_LC_13_10_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_30_9_LC_13_10_4 (
            .in0(N__41989),
            .in1(N__41312),
            .in2(_gnd_net_),
            .in3(N__27506),
            .lcout(),
            .ltout(sDAC_data_RNO_30Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_25_9_LC_13_10_5.C_ON=1'b0;
    defparam sDAC_data_RNO_25_9_LC_13_10_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_9_LC_13_10_5.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_25_9_LC_13_10_5 (
            .in0(N__38249),
            .in1(N__38477),
            .in2(N__27491),
            .in3(N__27695),
            .lcout(),
            .ltout(sDAC_data_2_39_ns_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_9_LC_13_10_6.C_ON=1'b0;
    defparam sDAC_data_RNO_11_9_LC_13_10_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_9_LC_13_10_6.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_11_9_LC_13_10_6 (
            .in0(N__29423),
            .in1(N__38250),
            .in2(N__27488),
            .in3(N__29636),
            .lcout(sDAC_data_RNO_11Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_31_9_LC_13_10_7.C_ON=1'b0;
    defparam sDAC_data_RNO_31_9_LC_13_10_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_9_LC_13_10_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_31_9_LC_13_10_7 (
            .in0(N__42013),
            .in1(N__29747),
            .in2(_gnd_net_),
            .in3(N__27710),
            .lcout(sDAC_data_RNO_31Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_30_7_LC_13_11_0.C_ON=1'b0;
    defparam sDAC_data_RNO_30_7_LC_13_11_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_7_LC_13_11_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_30_7_LC_13_11_0 (
            .in0(N__42018),
            .in1(N__41339),
            .in2(_gnd_net_),
            .in3(N__27596),
            .lcout(),
            .ltout(sDAC_data_RNO_30Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_25_7_LC_13_11_1.C_ON=1'b0;
    defparam sDAC_data_RNO_25_7_LC_13_11_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_7_LC_13_11_1.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_25_7_LC_13_11_1 (
            .in0(N__38262),
            .in1(N__38425),
            .in2(N__27689),
            .in3(N__27671),
            .lcout(),
            .ltout(sDAC_data_2_39_ns_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_7_LC_13_11_2.C_ON=1'b0;
    defparam sDAC_data_RNO_11_7_LC_13_11_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_7_LC_13_11_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_11_7_LC_13_11_2 (
            .in0(N__38202),
            .in1(N__27602),
            .in2(N__27686),
            .in3(N__27635),
            .lcout(sDAC_data_RNO_11Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_31_7_LC_13_11_3.C_ON=1'b0;
    defparam sDAC_data_RNO_31_7_LC_13_11_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_7_LC_13_11_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_31_7_LC_13_11_3 (
            .in0(N__29768),
            .in1(N__42015),
            .in2(_gnd_net_),
            .in3(N__27683),
            .lcout(sDAC_data_RNO_31Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_7_LC_13_11_4.C_ON=1'b0;
    defparam sDAC_data_RNO_23_7_LC_13_11_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_7_LC_13_11_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_7_LC_13_11_4 (
            .in0(N__42017),
            .in1(N__27665),
            .in2(_gnd_net_),
            .in3(N__27650),
            .lcout(sDAC_data_RNO_23Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_7_LC_13_11_5.C_ON=1'b0;
    defparam sDAC_data_RNO_24_7_LC_13_11_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_7_LC_13_11_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_24_7_LC_13_11_5 (
            .in0(N__27629),
            .in1(N__42016),
            .in2(_gnd_net_),
            .in3(N__27617),
            .lcout(sDAC_data_RNO_24Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_24_4_LC_13_11_6.C_ON=1'b0;
    defparam sDAC_mem_24_4_LC_13_11_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_4_LC_13_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_4_LC_13_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45585),
            .lcout(sDAC_mem_24Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52233),
            .ce(N__27741),
            .sr(N__51683));
    defparam sDAC_data_RNO_25_8_LC_13_11_7.C_ON=1'b0;
    defparam sDAC_data_RNO_25_8_LC_13_11_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_8_LC_13_11_7.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_25_8_LC_13_11_7 (
            .in0(N__38414),
            .in1(N__28064),
            .in2(N__38285),
            .in3(N__29450),
            .lcout(sDAC_data_2_39_ns_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_31_4_LC_13_12_0.C_ON=1'b0;
    defparam sDAC_data_RNO_31_4_LC_13_12_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_4_LC_13_12_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_31_4_LC_13_12_0 (
            .in0(N__41607),
            .in1(N__29570),
            .in2(_gnd_net_),
            .in3(N__27836),
            .lcout(sDAC_data_RNO_31Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_30_4_LC_13_12_1.C_ON=1'b0;
    defparam sDAC_data_RNO_30_4_LC_13_12_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_4_LC_13_12_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_30_4_LC_13_12_1 (
            .in0(N__42012),
            .in1(N__50609),
            .in2(_gnd_net_),
            .in3(N__27752),
            .lcout(),
            .ltout(sDAC_data_RNO_30Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_25_4_LC_13_12_2.C_ON=1'b0;
    defparam sDAC_data_RNO_25_4_LC_13_12_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_4_LC_13_12_2.LUT_INIT=16'b0100010101100111;
    LogicCell40 sDAC_data_RNO_25_4_LC_13_12_2 (
            .in0(N__38426),
            .in1(N__38216),
            .in2(N__27824),
            .in3(N__27821),
            .lcout(),
            .ltout(sDAC_data_2_39_ns_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_4_LC_13_12_3.C_ON=1'b0;
    defparam sDAC_data_RNO_11_4_LC_13_12_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_4_LC_13_12_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_11_4_LC_13_12_3 (
            .in0(N__38217),
            .in1(N__27758),
            .in2(N__27815),
            .in3(N__27788),
            .lcout(sDAC_data_RNO_11Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_4_LC_13_12_4.C_ON=1'b0;
    defparam sDAC_data_RNO_23_4_LC_13_12_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_4_LC_13_12_4.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_23_4_LC_13_12_4 (
            .in0(N__27812),
            .in1(N__42011),
            .in2(_gnd_net_),
            .in3(N__27800),
            .lcout(sDAC_data_RNO_23Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_4_LC_13_12_5.C_ON=1'b0;
    defparam sDAC_data_RNO_24_4_LC_13_12_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_4_LC_13_12_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_4_LC_13_12_5 (
            .in0(N__42010),
            .in1(N__27782),
            .in2(_gnd_net_),
            .in3(N__27770),
            .lcout(sDAC_data_RNO_24Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_24_1_LC_13_12_6.C_ON=1'b0;
    defparam sDAC_mem_24_1_LC_13_12_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_1_LC_13_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_1_LC_13_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51017),
            .lcout(sDAC_mem_24Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52243),
            .ce(N__27746),
            .sr(N__51677));
    defparam sDAC_data_RNO_25_5_LC_13_12_7.C_ON=1'b0;
    defparam sDAC_data_RNO_25_5_LC_13_12_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_5_LC_13_12_7.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_25_5_LC_13_12_7 (
            .in0(N__38387),
            .in1(N__28076),
            .in2(N__38254),
            .in3(N__29468),
            .lcout(sDAC_data_2_39_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_31_5_LC_13_13_0.C_ON=1'b0;
    defparam sDAC_data_RNO_31_5_LC_13_13_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_5_LC_13_13_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_31_5_LC_13_13_0 (
            .in0(N__41536),
            .in1(N__29777),
            .in2(_gnd_net_),
            .in3(N__28070),
            .lcout(sDAC_data_RNO_31Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_26_2_LC_13_13_1.C_ON=1'b0;
    defparam sDAC_mem_26_2_LC_13_13_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_2_LC_13_13_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_26_2_LC_13_13_1 (
            .in0(N__47506),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_26Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52253),
            .ce(N__28049),
            .sr(N__51669));
    defparam sDAC_data_RNO_31_8_LC_13_13_2.C_ON=1'b0;
    defparam sDAC_data_RNO_31_8_LC_13_13_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_8_LC_13_13_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_31_8_LC_13_13_2 (
            .in0(N__41537),
            .in1(N__29756),
            .in2(_gnd_net_),
            .in3(N__28055),
            .lcout(sDAC_data_RNO_31Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_26_5_LC_13_13_3.C_ON=1'b0;
    defparam sDAC_mem_26_5_LC_13_13_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_5_LC_13_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_26_5_LC_13_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45079),
            .lcout(sDAC_mem_26Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52253),
            .ce(N__28049),
            .sr(N__51669));
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_RNISHDJ_LC_13_13_5 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_RNISHDJ_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_RNISHDJ_LC_13_13_5 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_clk_i_RNISHDJ_LC_13_13_5  (
            .in0(N__27959),
            .in1(N__28025),
            .in2(_gnd_net_),
            .in3(N__28007),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNIK09A_LC_13_13_6 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNIK09A_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNIK09A_LC_13_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNIK09A_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27958),
            .lcout(\spi_master_inst.sclk_gen_u0.falling_count_start_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_0_c_LC_13_14_0.C_ON=1'b1;
    defparam un1_sacqtime_cry_0_c_LC_13_14_0.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_0_c_LC_13_14_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_0_c_LC_13_14_0 (
            .in0(_gnd_net_),
            .in1(N__27896),
            .in2(N__29119),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_14_0_),
            .carryout(un1_sacqtime_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_1_c_LC_13_14_1.C_ON=1'b1;
    defparam un1_sacqtime_cry_1_c_LC_13_14_1.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_1_c_LC_13_14_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_1_c_LC_13_14_1 (
            .in0(_gnd_net_),
            .in1(N__27878),
            .in2(N__29086),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_0),
            .carryout(un1_sacqtime_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_2_c_LC_13_14_2.C_ON=1'b1;
    defparam un1_sacqtime_cry_2_c_LC_13_14_2.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_2_c_LC_13_14_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_2_c_LC_13_14_2 (
            .in0(_gnd_net_),
            .in1(N__27857),
            .in2(N__29050),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_1),
            .carryout(un1_sacqtime_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_3_c_LC_13_14_3.C_ON=1'b1;
    defparam un1_sacqtime_cry_3_c_LC_13_14_3.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_3_c_LC_13_14_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_3_c_LC_13_14_3 (
            .in0(_gnd_net_),
            .in1(N__28235),
            .in2(N__29023),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_2),
            .carryout(un1_sacqtime_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_4_c_LC_13_14_4.C_ON=1'b1;
    defparam un1_sacqtime_cry_4_c_LC_13_14_4.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_4_c_LC_13_14_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_4_c_LC_13_14_4 (
            .in0(_gnd_net_),
            .in1(N__28214),
            .in2(N__28996),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_3),
            .carryout(un1_sacqtime_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_5_c_LC_13_14_5.C_ON=1'b1;
    defparam un1_sacqtime_cry_5_c_LC_13_14_5.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_5_c_LC_13_14_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_5_c_LC_13_14_5 (
            .in0(_gnd_net_),
            .in1(N__28193),
            .in2(N__28960),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_4),
            .carryout(un1_sacqtime_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_6_c_LC_13_14_6.C_ON=1'b1;
    defparam un1_sacqtime_cry_6_c_LC_13_14_6.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_6_c_LC_13_14_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_6_c_LC_13_14_6 (
            .in0(_gnd_net_),
            .in1(N__28175),
            .in2(N__28930),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_5),
            .carryout(un1_sacqtime_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_7_c_LC_13_14_7.C_ON=1'b1;
    defparam un1_sacqtime_cry_7_c_LC_13_14_7.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_7_c_LC_13_14_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_7_c_LC_13_14_7 (
            .in0(_gnd_net_),
            .in1(N__28154),
            .in2(N__29377),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_6),
            .carryout(un1_sacqtime_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_8_c_LC_13_15_0.C_ON=1'b1;
    defparam un1_sacqtime_cry_8_c_LC_13_15_0.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_8_c_LC_13_15_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_8_c_LC_13_15_0 (
            .in0(_gnd_net_),
            .in1(N__28136),
            .in2(N__29341),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(un1_sacqtime_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_9_c_LC_13_15_1.C_ON=1'b1;
    defparam un1_sacqtime_cry_9_c_LC_13_15_1.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_9_c_LC_13_15_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_9_c_LC_13_15_1 (
            .in0(_gnd_net_),
            .in1(N__28115),
            .in2(N__29308),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_8),
            .carryout(un1_sacqtime_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_10_c_LC_13_15_2.C_ON=1'b1;
    defparam un1_sacqtime_cry_10_c_LC_13_15_2.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_10_c_LC_13_15_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_10_c_LC_13_15_2 (
            .in0(_gnd_net_),
            .in1(N__28097),
            .in2(N__29278),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_9),
            .carryout(un1_sacqtime_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_11_c_LC_13_15_3.C_ON=1'b1;
    defparam un1_sacqtime_cry_11_c_LC_13_15_3.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_11_c_LC_13_15_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_11_c_LC_13_15_3 (
            .in0(_gnd_net_),
            .in1(N__28358),
            .in2(N__29248),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_10),
            .carryout(un1_sacqtime_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_12_c_LC_13_15_4.C_ON=1'b1;
    defparam un1_sacqtime_cry_12_c_LC_13_15_4.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_12_c_LC_13_15_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_12_c_LC_13_15_4 (
            .in0(_gnd_net_),
            .in1(N__28337),
            .in2(N__29212),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_11),
            .carryout(un1_sacqtime_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_13_c_LC_13_15_5.C_ON=1'b1;
    defparam un1_sacqtime_cry_13_c_LC_13_15_5.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_13_c_LC_13_15_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_13_c_LC_13_15_5 (
            .in0(_gnd_net_),
            .in1(N__28319),
            .in2(N__29182),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_12),
            .carryout(un1_sacqtime_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_14_c_LC_13_15_6.C_ON=1'b1;
    defparam un1_sacqtime_cry_14_c_LC_13_15_6.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_14_c_LC_13_15_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_14_c_LC_13_15_6 (
            .in0(_gnd_net_),
            .in1(N__28298),
            .in2(N__29155),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_13),
            .carryout(un1_sacqtime_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_15_c_LC_13_15_7.C_ON=1'b1;
    defparam un1_sacqtime_cry_15_c_LC_13_15_7.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_15_c_LC_13_15_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_15_c_LC_13_15_7 (
            .in0(_gnd_net_),
            .in1(N__28277),
            .in2(N__29407),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_14),
            .carryout(un1_sacqtime_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_16_c_inv_LC_13_16_0.C_ON=1'b1;
    defparam un1_sacqtime_cry_16_c_inv_LC_13_16_0.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_16_c_inv_LC_13_16_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_sacqtime_cry_16_c_inv_LC_13_16_0 (
            .in0(_gnd_net_),
            .in1(N__28259),
            .in2(_gnd_net_),
            .in3(N__31365),
            .lcout(un1_sacqtime_cry_16_sf),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(un1_sacqtime_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_17_c_inv_LC_13_16_1.C_ON=1'b1;
    defparam un1_sacqtime_cry_17_c_inv_LC_13_16_1.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_17_c_inv_LC_13_16_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_sacqtime_cry_17_c_inv_LC_13_16_1 (
            .in0(_gnd_net_),
            .in1(N__28253),
            .in2(_gnd_net_),
            .in3(N__31269),
            .lcout(un1_sacqtime_cry_17_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_16),
            .carryout(un1_sacqtime_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_18_c_inv_LC_13_16_2.C_ON=1'b1;
    defparam un1_sacqtime_cry_18_c_inv_LC_13_16_2.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_18_c_inv_LC_13_16_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_sacqtime_cry_18_c_inv_LC_13_16_2 (
            .in0(_gnd_net_),
            .in1(N__28247),
            .in2(_gnd_net_),
            .in3(N__31150),
            .lcout(un1_sacqtime_cry_18_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_17),
            .carryout(un1_sacqtime_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_19_c_inv_LC_13_16_3.C_ON=1'b1;
    defparam un1_sacqtime_cry_19_c_inv_LC_13_16_3.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_19_c_inv_LC_13_16_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_sacqtime_cry_19_c_inv_LC_13_16_3 (
            .in0(N__33253),
            .in1(N__28241),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_sacqtime_cry_19_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_18),
            .carryout(un1_sacqtime_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_20_c_inv_LC_13_16_4.C_ON=1'b1;
    defparam un1_sacqtime_cry_20_c_inv_LC_13_16_4.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_20_c_inv_LC_13_16_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_sacqtime_cry_20_c_inv_LC_13_16_4 (
            .in0(_gnd_net_),
            .in1(N__28403),
            .in2(_gnd_net_),
            .in3(N__33373),
            .lcout(un1_sacqtime_cry_20_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_19),
            .carryout(un1_sacqtime_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_21_c_inv_LC_13_16_5.C_ON=1'b1;
    defparam un1_sacqtime_cry_21_c_inv_LC_13_16_5.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_21_c_inv_LC_13_16_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_sacqtime_cry_21_c_inv_LC_13_16_5 (
            .in0(_gnd_net_),
            .in1(N__28397),
            .in2(_gnd_net_),
            .in3(N__33154),
            .lcout(un1_sacqtime_cry_21_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_20),
            .carryout(un1_sacqtime_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_22_c_inv_LC_13_16_6.C_ON=1'b1;
    defparam un1_sacqtime_cry_22_c_inv_LC_13_16_6.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_22_c_inv_LC_13_16_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_sacqtime_cry_22_c_inv_LC_13_16_6 (
            .in0(N__32027),
            .in1(N__28391),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_sacqtime_cry_22_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_21),
            .carryout(un1_sacqtime_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_23_c_inv_LC_13_16_7.C_ON=1'b1;
    defparam un1_sacqtime_cry_23_c_inv_LC_13_16_7.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_23_c_inv_LC_13_16_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_sacqtime_cry_23_c_inv_LC_13_16_7 (
            .in0(_gnd_net_),
            .in1(N__28385),
            .in2(_gnd_net_),
            .in3(N__31913),
            .lcout(un1_sacqtime_cry_23_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_22),
            .carryout(un1_sacqtime_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_23_THRU_LUT4_0_LC_13_17_0.C_ON=1'b0;
    defparam un1_sacqtime_cry_23_THRU_LUT4_0_LC_13_17_0.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_23_THRU_LUT4_0_LC_13_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_sacqtime_cry_23_THRU_LUT4_0_LC_13_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28379),
            .lcout(un1_sacqtime_cry_23_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sADC_clk_prev_LC_13_17_1.C_ON=1'b0;
    defparam sADC_clk_prev_LC_13_17_1.SEQ_MODE=4'b1000;
    defparam sADC_clk_prev_LC_13_17_1.LUT_INIT=16'b1011100011110000;
    LogicCell40 sADC_clk_prev_LC_13_17_1 (
            .in0(N__34014),
            .in1(N__49381),
            .in2(N__28376),
            .in3(N__48962),
            .lcout(sADC_clk_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52299),
            .ce(),
            .sr(_gnd_net_));
    defparam sADC_clk_prev_RNI4BVG_LC_13_17_6.C_ON=1'b0;
    defparam sADC_clk_prev_RNI4BVG_LC_13_17_6.SEQ_MODE=4'b0000;
    defparam sADC_clk_prev_RNI4BVG_LC_13_17_6.LUT_INIT=16'b1100110011111111;
    LogicCell40 sADC_clk_prev_RNI4BVG_LC_13_17_6 (
            .in0(_gnd_net_),
            .in1(N__28372),
            .in2(_gnd_net_),
            .in3(N__34013),
            .lcout(N_71),
            .ltout(N_71_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_23_c_RNIJ7QO_LC_13_17_7.C_ON=1'b0;
    defparam un4_sacqtime_cry_23_c_RNIJ7QO_LC_13_17_7.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_23_c_RNIJ7QO_LC_13_17_7.LUT_INIT=16'b0000100000000000;
    LogicCell40 un4_sacqtime_cry_23_c_RNIJ7QO_LC_13_17_7 (
            .in0(N__49382),
            .in1(N__43439),
            .in2(N__28364),
            .in3(N__43316),
            .lcout(N_31_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sRAM_pointer_read_0_LC_13_18_0.C_ON=1'b1;
    defparam sRAM_pointer_read_0_LC_13_18_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_0_LC_13_18_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_0_LC_13_18_0 (
            .in0(N__39344),
            .in1(N__35902),
            .in2(_gnd_net_),
            .in3(N__28361),
            .lcout(sRAM_pointer_readZ0Z_0),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(sRAM_pointer_read_cry_0),
            .clk(N__52309),
            .ce(N__28445),
            .sr(N__51646));
    defparam sRAM_pointer_read_1_LC_13_18_1.C_ON=1'b1;
    defparam sRAM_pointer_read_1_LC_13_18_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_1_LC_13_18_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_1_LC_13_18_1 (
            .in0(N__39340),
            .in1(N__36040),
            .in2(_gnd_net_),
            .in3(N__28430),
            .lcout(sRAM_pointer_readZ0Z_1),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_0),
            .carryout(sRAM_pointer_read_cry_1),
            .clk(N__52309),
            .ce(N__28445),
            .sr(N__51646));
    defparam sRAM_pointer_read_2_LC_13_18_2.C_ON=1'b1;
    defparam sRAM_pointer_read_2_LC_13_18_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_2_LC_13_18_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_2_LC_13_18_2 (
            .in0(N__39345),
            .in1(N__36130),
            .in2(_gnd_net_),
            .in3(N__28427),
            .lcout(sRAM_pointer_readZ0Z_2),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_1),
            .carryout(sRAM_pointer_read_cry_2),
            .clk(N__52309),
            .ce(N__28445),
            .sr(N__51646));
    defparam sRAM_pointer_read_3_LC_13_18_3.C_ON=1'b1;
    defparam sRAM_pointer_read_3_LC_13_18_3.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_3_LC_13_18_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_3_LC_13_18_3 (
            .in0(N__39341),
            .in1(N__43366),
            .in2(_gnd_net_),
            .in3(N__28424),
            .lcout(sRAM_pointer_readZ0Z_3),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_2),
            .carryout(sRAM_pointer_read_cry_3),
            .clk(N__52309),
            .ce(N__28445),
            .sr(N__51646));
    defparam sRAM_pointer_read_4_LC_13_18_4.C_ON=1'b1;
    defparam sRAM_pointer_read_4_LC_13_18_4.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_4_LC_13_18_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_4_LC_13_18_4 (
            .in0(N__39346),
            .in1(N__43549),
            .in2(_gnd_net_),
            .in3(N__28421),
            .lcout(sRAM_pointer_readZ0Z_4),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_3),
            .carryout(sRAM_pointer_read_cry_4),
            .clk(N__52309),
            .ce(N__28445),
            .sr(N__51646));
    defparam sRAM_pointer_read_5_LC_13_18_5.C_ON=1'b1;
    defparam sRAM_pointer_read_5_LC_13_18_5.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_5_LC_13_18_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_5_LC_13_18_5 (
            .in0(N__39342),
            .in1(N__35248),
            .in2(_gnd_net_),
            .in3(N__28418),
            .lcout(sRAM_pointer_readZ0Z_5),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_4),
            .carryout(sRAM_pointer_read_cry_5),
            .clk(N__52309),
            .ce(N__28445),
            .sr(N__51646));
    defparam sRAM_pointer_read_6_LC_13_18_6.C_ON=1'b1;
    defparam sRAM_pointer_read_6_LC_13_18_6.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_6_LC_13_18_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_6_LC_13_18_6 (
            .in0(N__39347),
            .in1(N__35983),
            .in2(_gnd_net_),
            .in3(N__28415),
            .lcout(sRAM_pointer_readZ0Z_6),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_5),
            .carryout(sRAM_pointer_read_cry_6),
            .clk(N__52309),
            .ce(N__28445),
            .sr(N__51646));
    defparam sRAM_pointer_read_7_LC_13_18_7.C_ON=1'b1;
    defparam sRAM_pointer_read_7_LC_13_18_7.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_7_LC_13_18_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_7_LC_13_18_7 (
            .in0(N__39343),
            .in1(N__36163),
            .in2(_gnd_net_),
            .in3(N__28412),
            .lcout(sRAM_pointer_readZ0Z_7),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_6),
            .carryout(sRAM_pointer_read_cry_7),
            .clk(N__52309),
            .ce(N__28445),
            .sr(N__51646));
    defparam sRAM_pointer_read_8_LC_13_19_0.C_ON=1'b1;
    defparam sRAM_pointer_read_8_LC_13_19_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_8_LC_13_19_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_8_LC_13_19_0 (
            .in0(N__39395),
            .in1(N__43621),
            .in2(_gnd_net_),
            .in3(N__28409),
            .lcout(sRAM_pointer_readZ0Z_8),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(sRAM_pointer_read_cry_8),
            .clk(N__52322),
            .ce(N__28444),
            .sr(N__51645));
    defparam sRAM_pointer_read_9_LC_13_19_1.C_ON=1'b1;
    defparam sRAM_pointer_read_9_LC_13_19_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_9_LC_13_19_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_9_LC_13_19_1 (
            .in0(N__39391),
            .in1(N__36229),
            .in2(_gnd_net_),
            .in3(N__28406),
            .lcout(sRAM_pointer_readZ0Z_9),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_8),
            .carryout(sRAM_pointer_read_cry_9),
            .clk(N__52322),
            .ce(N__28444),
            .sr(N__51645));
    defparam sRAM_pointer_read_10_LC_13_19_2.C_ON=1'b1;
    defparam sRAM_pointer_read_10_LC_13_19_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_10_LC_13_19_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_10_LC_13_19_2 (
            .in0(N__39392),
            .in1(N__35839),
            .in2(_gnd_net_),
            .in3(N__28472),
            .lcout(sRAM_pointer_readZ0Z_10),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_9),
            .carryout(sRAM_pointer_read_cry_10),
            .clk(N__52322),
            .ce(N__28444),
            .sr(N__51645));
    defparam sRAM_pointer_read_11_LC_13_19_3.C_ON=1'b1;
    defparam sRAM_pointer_read_11_LC_13_19_3.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_11_LC_13_19_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_11_LC_13_19_3 (
            .in0(N__39388),
            .in1(N__35767),
            .in2(_gnd_net_),
            .in3(N__28469),
            .lcout(sRAM_pointer_readZ0Z_11),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_10),
            .carryout(sRAM_pointer_read_cry_11),
            .clk(N__52322),
            .ce(N__28444),
            .sr(N__51645));
    defparam sRAM_pointer_read_12_LC_13_19_4.C_ON=1'b1;
    defparam sRAM_pointer_read_12_LC_13_19_4.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_12_LC_13_19_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_12_LC_13_19_4 (
            .in0(N__39393),
            .in1(N__35671),
            .in2(_gnd_net_),
            .in3(N__28466),
            .lcout(sRAM_pointer_readZ0Z_12),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_11),
            .carryout(sRAM_pointer_read_cry_12),
            .clk(N__52322),
            .ce(N__28444),
            .sr(N__51645));
    defparam sRAM_pointer_read_13_LC_13_19_5.C_ON=1'b1;
    defparam sRAM_pointer_read_13_LC_13_19_5.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_13_LC_13_19_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_13_LC_13_19_5 (
            .in0(N__39389),
            .in1(N__35632),
            .in2(_gnd_net_),
            .in3(N__28463),
            .lcout(sRAM_pointer_readZ0Z_13),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_12),
            .carryout(sRAM_pointer_read_cry_13),
            .clk(N__52322),
            .ce(N__28444),
            .sr(N__51645));
    defparam sRAM_pointer_read_14_LC_13_19_6.C_ON=1'b1;
    defparam sRAM_pointer_read_14_LC_13_19_6.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_14_LC_13_19_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_14_LC_13_19_6 (
            .in0(N__39394),
            .in1(N__35539),
            .in2(_gnd_net_),
            .in3(N__28460),
            .lcout(sRAM_pointer_readZ0Z_14),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_13),
            .carryout(sRAM_pointer_read_cry_14),
            .clk(N__52322),
            .ce(N__28444),
            .sr(N__51645));
    defparam sRAM_pointer_read_15_LC_13_19_7.C_ON=1'b1;
    defparam sRAM_pointer_read_15_LC_13_19_7.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_15_LC_13_19_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_15_LC_13_19_7 (
            .in0(N__39390),
            .in1(N__35497),
            .in2(_gnd_net_),
            .in3(N__28457),
            .lcout(sRAM_pointer_readZ0Z_15),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_14),
            .carryout(sRAM_pointer_read_cry_15),
            .clk(N__52322),
            .ce(N__28444),
            .sr(N__51645));
    defparam sRAM_pointer_read_16_LC_13_20_0.C_ON=1'b1;
    defparam sRAM_pointer_read_16_LC_13_20_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_16_LC_13_20_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_16_LC_13_20_0 (
            .in0(N__39296),
            .in1(N__35425),
            .in2(_gnd_net_),
            .in3(N__28454),
            .lcout(sRAM_pointer_readZ0Z_16),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(sRAM_pointer_read_cry_16),
            .clk(N__52330),
            .ce(N__28443),
            .sr(N__51643));
    defparam sRAM_pointer_read_17_LC_13_20_1.C_ON=1'b1;
    defparam sRAM_pointer_read_17_LC_13_20_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_17_LC_13_20_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_17_LC_13_20_1 (
            .in0(N__39295),
            .in1(N__36367),
            .in2(_gnd_net_),
            .in3(N__28451),
            .lcout(sRAM_pointer_readZ0Z_17),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_16),
            .carryout(sRAM_pointer_read_cry_17),
            .clk(N__52330),
            .ce(N__28443),
            .sr(N__51643));
    defparam sRAM_pointer_read_18_LC_13_20_2.C_ON=1'b0;
    defparam sRAM_pointer_read_18_LC_13_20_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_18_LC_13_20_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_18_LC_13_20_2 (
            .in0(N__39297),
            .in1(N__36301),
            .in2(_gnd_net_),
            .in3(N__28448),
            .lcout(sRAM_pointer_readZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52330),
            .ce(N__28443),
            .sr(N__51643));
    defparam sDAC_mem_36_0_LC_14_3_0.C_ON=1'b0;
    defparam sDAC_mem_36_0_LC_14_3_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_0_LC_14_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_0_LC_14_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46145),
            .lcout(sDAC_mem_36Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52310),
            .ce(N__28484),
            .sr(N__51782));
    defparam sDAC_mem_36_1_LC_14_3_1.C_ON=1'b0;
    defparam sDAC_mem_36_1_LC_14_3_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_1_LC_14_3_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_1_LC_14_3_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51074),
            .lcout(sDAC_mem_36Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52310),
            .ce(N__28484),
            .sr(N__51782));
    defparam sDAC_mem_36_2_LC_14_3_2.C_ON=1'b0;
    defparam sDAC_mem_36_2_LC_14_3_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_2_LC_14_3_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_2_LC_14_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47328),
            .lcout(sDAC_mem_36Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52310),
            .ce(N__28484),
            .sr(N__51782));
    defparam sDAC_mem_36_3_LC_14_3_3.C_ON=1'b0;
    defparam sDAC_mem_36_3_LC_14_3_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_3_LC_14_3_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_3_LC_14_3_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46901),
            .lcout(sDAC_mem_36Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52310),
            .ce(N__28484),
            .sr(N__51782));
    defparam sDAC_mem_36_4_LC_14_3_4.C_ON=1'b0;
    defparam sDAC_mem_36_4_LC_14_3_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_4_LC_14_3_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_4_LC_14_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45530),
            .lcout(sDAC_mem_36Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52310),
            .ce(N__28484),
            .sr(N__51782));
    defparam sDAC_mem_36_5_LC_14_3_5.C_ON=1'b0;
    defparam sDAC_mem_36_5_LC_14_3_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_5_LC_14_3_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_5_LC_14_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45055),
            .lcout(sDAC_mem_36Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52310),
            .ce(N__28484),
            .sr(N__51782));
    defparam sDAC_mem_36_6_LC_14_3_6.C_ON=1'b0;
    defparam sDAC_mem_36_6_LC_14_3_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_6_LC_14_3_6.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_36_6_LC_14_3_6 (
            .in0(_gnd_net_),
            .in1(N__50408),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_36Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52310),
            .ce(N__28484),
            .sr(N__51782));
    defparam sDAC_mem_36_7_LC_14_3_7.C_ON=1'b0;
    defparam sDAC_mem_36_7_LC_14_3_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_7_LC_14_3_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_7_LC_14_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49996),
            .lcout(sDAC_mem_36Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52310),
            .ce(N__28484),
            .sr(N__51782));
    defparam sDAC_data_RNO_29_6_LC_14_4_0.C_ON=1'b0;
    defparam sDAC_data_RNO_29_6_LC_14_4_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_6_LC_14_4_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_29_6_LC_14_4_0 (
            .in0(N__41813),
            .in1(N__35012),
            .in2(_gnd_net_),
            .in3(N__28577),
            .lcout(sDAC_data_RNO_29Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_18_3_LC_14_4_1.C_ON=1'b0;
    defparam sDAC_mem_18_3_LC_14_4_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_3_LC_14_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_3_LC_14_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46746),
            .lcout(sDAC_mem_18Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52300),
            .ce(N__28544),
            .sr(N__51769));
    defparam sDAC_data_RNO_29_7_LC_14_4_2.C_ON=1'b0;
    defparam sDAC_data_RNO_29_7_LC_14_4_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_7_LC_14_4_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_29_7_LC_14_4_2 (
            .in0(N__41810),
            .in1(N__33923),
            .in2(_gnd_net_),
            .in3(N__28571),
            .lcout(sDAC_data_RNO_29Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_18_4_LC_14_4_3.C_ON=1'b0;
    defparam sDAC_mem_18_4_LC_14_4_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_4_LC_14_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_4_LC_14_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45528),
            .lcout(sDAC_mem_18Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52300),
            .ce(N__28544),
            .sr(N__51769));
    defparam sDAC_data_RNO_29_8_LC_14_4_4.C_ON=1'b0;
    defparam sDAC_data_RNO_29_8_LC_14_4_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_8_LC_14_4_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_29_8_LC_14_4_4 (
            .in0(N__41811),
            .in1(N__33911),
            .in2(_gnd_net_),
            .in3(N__28556),
            .lcout(sDAC_data_RNO_29Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_18_5_LC_14_4_5.C_ON=1'b0;
    defparam sDAC_mem_18_5_LC_14_4_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_5_LC_14_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_5_LC_14_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45054),
            .lcout(sDAC_mem_18Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52300),
            .ce(N__28544),
            .sr(N__51769));
    defparam sDAC_data_RNO_29_9_LC_14_4_6.C_ON=1'b0;
    defparam sDAC_data_RNO_29_9_LC_14_4_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_9_LC_14_4_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_29_9_LC_14_4_6 (
            .in0(N__41812),
            .in1(N__34091),
            .in2(_gnd_net_),
            .in3(N__28550),
            .lcout(sDAC_data_RNO_29Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_18_6_LC_14_4_7.C_ON=1'b0;
    defparam sDAC_mem_18_6_LC_14_4_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_6_LC_14_4_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_6_LC_14_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50407),
            .lcout(sDAC_mem_18Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52300),
            .ce(N__28544),
            .sr(N__51769));
    defparam sDAC_data_RNO_19_7_LC_14_5_0.C_ON=1'b0;
    defparam sDAC_data_RNO_19_7_LC_14_5_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_7_LC_14_5_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_7_LC_14_5_0 (
            .in0(N__42093),
            .in1(N__28517),
            .in2(_gnd_net_),
            .in3(N__28505),
            .lcout(sDAC_data_RNO_19Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_7_LC_14_5_1.C_ON=1'b0;
    defparam sDAC_data_RNO_18_7_LC_14_5_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_7_LC_14_5_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_7_LC_14_5_1 (
            .in0(N__42233),
            .in1(N__45134),
            .in2(_gnd_net_),
            .in3(N__28619),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_7_LC_14_5_2.C_ON=1'b0;
    defparam sDAC_data_RNO_9_7_LC_14_5_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_7_LC_14_5_2.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_9_7_LC_14_5_2 (
            .in0(N__38129),
            .in1(N__38553),
            .in2(N__28493),
            .in3(N__28490),
            .lcout(sDAC_data_2_24_ns_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_8_LC_14_5_3.C_ON=1'b0;
    defparam sDAC_data_RNO_18_8_LC_14_5_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_8_LC_14_5_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_8_LC_14_5_3 (
            .in0(N__42234),
            .in1(N__44624),
            .in2(_gnd_net_),
            .in3(N__28613),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_8_LC_14_5_4.C_ON=1'b0;
    defparam sDAC_data_RNO_9_8_LC_14_5_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_8_LC_14_5_4.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_9_8_LC_14_5_4 (
            .in0(N__38130),
            .in1(N__38554),
            .in2(N__28658),
            .in3(N__28625),
            .lcout(sDAC_data_2_24_ns_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_19_8_LC_14_5_5.C_ON=1'b0;
    defparam sDAC_data_RNO_19_8_LC_14_5_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_8_LC_14_5_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_8_LC_14_5_5 (
            .in0(N__42232),
            .in1(N__28649),
            .in2(_gnd_net_),
            .in3(N__28637),
            .lcout(sDAC_data_RNO_19Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_12_4_LC_14_5_6.C_ON=1'b0;
    defparam sDAC_mem_12_4_LC_14_5_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_4_LC_14_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_4_LC_14_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45348),
            .lcout(sDAC_mem_12Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52288),
            .ce(N__36960),
            .sr(N__51756));
    defparam sDAC_mem_12_5_LC_14_5_7.C_ON=1'b0;
    defparam sDAC_mem_12_5_LC_14_5_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_5_LC_14_5_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_12_5_LC_14_5_7 (
            .in0(N__44867),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_12Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52288),
            .ce(N__36960),
            .sr(N__51756));
    defparam sDAC_data_RNO_13_5_LC_14_6_0.C_ON=1'b0;
    defparam sDAC_data_RNO_13_5_LC_14_6_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_5_LC_14_6_0.LUT_INIT=16'b0011010000110111;
    LogicCell40 sDAC_data_RNO_13_5_LC_14_6_0 (
            .in0(N__28607),
            .in1(N__42567),
            .in2(N__42192),
            .in3(N__28583),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_5_LC_14_6_1.C_ON=1'b0;
    defparam sDAC_data_RNO_5_5_LC_14_6_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_5_LC_14_6_1.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_5_5_LC_14_6_1 (
            .in0(N__42067),
            .in1(N__28598),
            .in2(N__28586),
            .in3(N__43835),
            .lcout(sDAC_data_RNO_5Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_6_2_LC_14_6_2.C_ON=1'b0;
    defparam sDAC_mem_6_2_LC_14_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_2_LC_14_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_2_LC_14_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47364),
            .lcout(sDAC_mem_6Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52275),
            .ce(N__36549),
            .sr(N__51744));
    defparam sDAC_data_RNO_13_6_LC_14_6_3.C_ON=1'b0;
    defparam sDAC_data_RNO_13_6_LC_14_6_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_6_LC_14_6_3.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_13_6_LC_14_6_3 (
            .in0(N__42568),
            .in1(N__28745),
            .in2(N__42203),
            .in3(N__28712),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_6_LC_14_6_4.C_ON=1'b0;
    defparam sDAC_data_RNO_5_6_LC_14_6_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_6_LC_14_6_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_5_6_LC_14_6_4 (
            .in0(N__42052),
            .in1(N__28733),
            .in2(N__28721),
            .in3(N__43820),
            .lcout(sDAC_data_RNO_5Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_6_3_LC_14_6_5.C_ON=1'b0;
    defparam sDAC_mem_6_3_LC_14_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_3_LC_14_6_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_6_3_LC_14_6_5 (
            .in0(N__46794),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_6Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52275),
            .ce(N__36549),
            .sr(N__51744));
    defparam sDAC_data_RNO_13_7_LC_14_6_6.C_ON=1'b0;
    defparam sDAC_data_RNO_13_7_LC_14_6_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_7_LC_14_6_6.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_13_7_LC_14_6_6 (
            .in0(N__42559),
            .in1(N__28706),
            .in2(N__42193),
            .in3(N__36581),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_7_LC_14_6_7.C_ON=1'b0;
    defparam sDAC_data_RNO_5_7_LC_14_6_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_7_LC_14_6_7.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_5_7_LC_14_6_7 (
            .in0(N__42068),
            .in1(N__28697),
            .in2(N__28682),
            .in3(N__44312),
            .lcout(sDAC_data_RNO_5Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_28_6_LC_14_7_0.C_ON=1'b0;
    defparam sDAC_data_RNO_28_6_LC_14_7_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_6_LC_14_7_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_28_6_LC_14_7_0 (
            .in0(N__41873),
            .in1(N__38612),
            .in2(_gnd_net_),
            .in3(N__28670),
            .lcout(sDAC_data_RNO_28Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_16_3_LC_14_7_1.C_ON=1'b0;
    defparam sDAC_mem_16_3_LC_14_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_3_LC_14_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_3_LC_14_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46891),
            .lcout(sDAC_mem_16Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52266),
            .ce(N__33508),
            .sr(N__51729));
    defparam sDAC_data_RNO_28_7_LC_14_7_2.C_ON=1'b0;
    defparam sDAC_data_RNO_28_7_LC_14_7_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_7_LC_14_7_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_28_7_LC_14_7_2 (
            .in0(N__41872),
            .in1(N__39008),
            .in2(_gnd_net_),
            .in3(N__28664),
            .lcout(sDAC_data_RNO_28Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_16_4_LC_14_7_3.C_ON=1'b0;
    defparam sDAC_mem_16_4_LC_14_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_4_LC_14_7_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_16_4_LC_14_7_3 (
            .in0(N__45531),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_16Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52266),
            .ce(N__33508),
            .sr(N__51729));
    defparam sDAC_data_RNO_28_8_LC_14_7_4.C_ON=1'b0;
    defparam sDAC_data_RNO_28_8_LC_14_7_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_8_LC_14_7_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_28_8_LC_14_7_4 (
            .in0(N__41874),
            .in1(N__38993),
            .in2(_gnd_net_),
            .in3(N__28808),
            .lcout(sDAC_data_RNO_28Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_16_5_LC_14_7_5.C_ON=1'b0;
    defparam sDAC_mem_16_5_LC_14_7_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_5_LC_14_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_5_LC_14_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45081),
            .lcout(sDAC_mem_16Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52266),
            .ce(N__33508),
            .sr(N__51729));
    defparam sDAC_data_RNO_28_9_LC_14_7_6.C_ON=1'b0;
    defparam sDAC_data_RNO_28_9_LC_14_7_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_9_LC_14_7_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_28_9_LC_14_7_6 (
            .in0(N__41875),
            .in1(N__38978),
            .in2(_gnd_net_),
            .in3(N__28802),
            .lcout(sDAC_data_RNO_28Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_16_6_LC_14_7_7.C_ON=1'b0;
    defparam sDAC_mem_16_6_LC_14_7_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_6_LC_14_7_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_16_6_LC_14_7_7 (
            .in0(_gnd_net_),
            .in1(N__50468),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_16Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52266),
            .ce(N__33508),
            .sr(N__51729));
    defparam sDAC_data_RNO_10_4_LC_14_8_0.C_ON=1'b0;
    defparam sDAC_data_RNO_10_4_LC_14_8_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_4_LC_14_8_0.LUT_INIT=16'b1010000011001111;
    LogicCell40 sDAC_data_RNO_10_4_LC_14_8_0 (
            .in0(N__34436),
            .in1(N__32384),
            .in2(N__38210),
            .in3(N__28898),
            .lcout(),
            .ltout(sDAC_data_RNO_10Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_4_LC_14_8_1.C_ON=1'b0;
    defparam sDAC_data_RNO_3_4_LC_14_8_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_4_LC_14_8_1.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_3_4_LC_14_8_1 (
            .in0(N__37439),
            .in1(N__37344),
            .in2(N__28796),
            .in3(N__28793),
            .lcout(sDAC_data_2_41_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_4_LC_14_8_2.C_ON=1'b0;
    defparam sDAC_data_RNO_1_4_LC_14_8_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_4_LC_14_8_2.LUT_INIT=16'b1010000011001111;
    LogicCell40 sDAC_data_RNO_1_4_LC_14_8_2 (
            .in0(N__41144),
            .in1(N__28781),
            .in2(N__38211),
            .in3(N__28904),
            .lcout(),
            .ltout(sDAC_data_RNO_1Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_4_LC_14_8_3.C_ON=1'b0;
    defparam sDAC_data_RNO_0_4_LC_14_8_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_4_LC_14_8_3.LUT_INIT=16'b0101000011101110;
    LogicCell40 sDAC_data_RNO_0_4_LC_14_8_3 (
            .in0(N__37440),
            .in1(N__28769),
            .in2(N__28763),
            .in3(N__28760),
            .lcout(),
            .ltout(sDAC_data_2_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_4_LC_14_8_4.C_ON=1'b0;
    defparam sDAC_data_4_LC_14_8_4.SEQ_MODE=4'b1010;
    defparam sDAC_data_4_LC_14_8_4.LUT_INIT=16'b1110010011100100;
    LogicCell40 sDAC_data_4_LC_14_8_4 (
            .in0(N__37628),
            .in1(N__32111),
            .in2(N__28754),
            .in3(_gnd_net_),
            .lcout(sDAC_dataZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48457),
            .ce(N__43950),
            .sr(N__51717));
    defparam sDAC_data_RNO_6_4_LC_14_8_5.C_ON=1'b0;
    defparam sDAC_data_RNO_6_4_LC_14_8_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_4_LC_14_8_5.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_6_4_LC_14_8_5 (
            .in0(N__38558),
            .in1(N__28751),
            .in2(N__38212),
            .in3(N__41045),
            .lcout(sDAC_data_2_14_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_4_LC_14_8_6.C_ON=1'b0;
    defparam sDAC_data_RNO_22_4_LC_14_8_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_4_LC_14_8_6.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_22_4_LC_14_8_6 (
            .in0(N__38555),
            .in1(N__34787),
            .in2(N__38209),
            .in3(N__29594),
            .lcout(sDAC_data_2_32_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_19_5_LC_14_9_0.C_ON=1'b0;
    defparam sDAC_data_RNO_19_5_LC_14_9_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_5_LC_14_9_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_5_LC_14_9_0 (
            .in0(N__42082),
            .in1(N__28892),
            .in2(_gnd_net_),
            .in3(N__28883),
            .lcout(sDAC_data_RNO_19Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_5_LC_14_9_1.C_ON=1'b0;
    defparam sDAC_data_RNO_18_5_LC_14_9_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_5_LC_14_9_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_5_LC_14_9_1 (
            .in0(N__41809),
            .in1(N__45638),
            .in2(_gnd_net_),
            .in3(N__28820),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_5_LC_14_9_2.C_ON=1'b0;
    defparam sDAC_data_RNO_9_5_LC_14_9_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_5_LC_14_9_2.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_9_5_LC_14_9_2 (
            .in0(N__38168),
            .in1(N__38551),
            .in2(N__28871),
            .in3(N__28868),
            .lcout(sDAC_data_2_24_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_6_LC_14_9_3.C_ON=1'b0;
    defparam sDAC_data_RNO_18_6_LC_14_9_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_6_LC_14_9_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_6_LC_14_9_3 (
            .in0(N__41808),
            .in1(N__45623),
            .in2(_gnd_net_),
            .in3(N__29126),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_6_LC_14_9_4.C_ON=1'b0;
    defparam sDAC_data_RNO_9_6_LC_14_9_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_6_LC_14_9_4.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_9_6_LC_14_9_4 (
            .in0(N__38169),
            .in1(N__38550),
            .in2(N__28862),
            .in3(N__28826),
            .lcout(sDAC_data_2_24_ns_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_19_6_LC_14_9_5.C_ON=1'b0;
    defparam sDAC_data_RNO_19_6_LC_14_9_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_6_LC_14_9_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_19_6_LC_14_9_5 (
            .in0(N__28847),
            .in1(N__42081),
            .in2(_gnd_net_),
            .in3(N__28838),
            .lcout(sDAC_data_RNO_19Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_12_2_LC_14_9_6.C_ON=1'b0;
    defparam sDAC_mem_12_2_LC_14_9_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_2_LC_14_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_2_LC_14_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47345),
            .lcout(sDAC_mem_12Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52244),
            .ce(N__36965),
            .sr(N__51706));
    defparam sDAC_mem_12_3_LC_14_9_7.C_ON=1'b0;
    defparam sDAC_mem_12_3_LC_14_9_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_3_LC_14_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_3_LC_14_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46853),
            .lcout(sDAC_mem_12Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52244),
            .ce(N__36965),
            .sr(N__51706));
    defparam un5_sdacdyn_cry_0_c_inv_LC_14_10_0.C_ON=1'b1;
    defparam un5_sdacdyn_cry_0_c_inv_LC_14_10_0.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_0_c_inv_LC_14_10_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_0_c_inv_LC_14_10_0 (
            .in0(_gnd_net_),
            .in1(N__30216),
            .in2(N__29096),
            .in3(N__29120),
            .lcout(sEEACQ_i_0),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(un5_sdacdyn_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_1_c_inv_LC_14_10_1.C_ON=1'b1;
    defparam un5_sdacdyn_cry_1_c_inv_LC_14_10_1.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_1_c_inv_LC_14_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_1_c_inv_LC_14_10_1 (
            .in0(_gnd_net_),
            .in1(N__30096),
            .in2(N__29063),
            .in3(N__29087),
            .lcout(sEEACQ_i_1),
            .ltout(),
            .carryin(un5_sdacdyn_cry_0),
            .carryout(un5_sdacdyn_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_2_c_inv_LC_14_10_2.C_ON=1'b1;
    defparam un5_sdacdyn_cry_2_c_inv_LC_14_10_2.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_2_c_inv_LC_14_10_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_2_c_inv_LC_14_10_2 (
            .in0(_gnd_net_),
            .in1(N__29033),
            .in2(N__29997),
            .in3(N__29054),
            .lcout(sEEACQ_i_2),
            .ltout(),
            .carryin(un5_sdacdyn_cry_1),
            .carryout(un5_sdacdyn_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_3_c_inv_LC_14_10_3.C_ON=1'b1;
    defparam un5_sdacdyn_cry_3_c_inv_LC_14_10_3.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_3_c_inv_LC_14_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_3_c_inv_LC_14_10_3 (
            .in0(_gnd_net_),
            .in1(N__29871),
            .in2(N__29006),
            .in3(N__29027),
            .lcout(sEEACQ_i_3),
            .ltout(),
            .carryin(un5_sdacdyn_cry_2),
            .carryout(un5_sdacdyn_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_4_c_inv_LC_14_10_4.C_ON=1'b1;
    defparam un5_sdacdyn_cry_4_c_inv_LC_14_10_4.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_4_c_inv_LC_14_10_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_4_c_inv_LC_14_10_4 (
            .in0(_gnd_net_),
            .in1(N__31001),
            .in2(N__28973),
            .in3(N__28997),
            .lcout(sEEACQ_i_4),
            .ltout(),
            .carryin(un5_sdacdyn_cry_3),
            .carryout(un5_sdacdyn_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_5_c_inv_LC_14_10_5.C_ON=1'b1;
    defparam un5_sdacdyn_cry_5_c_inv_LC_14_10_5.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_5_c_inv_LC_14_10_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_5_c_inv_LC_14_10_5 (
            .in0(_gnd_net_),
            .in1(N__30881),
            .in2(N__28943),
            .in3(N__28964),
            .lcout(sEEACQ_i_5),
            .ltout(),
            .carryin(un5_sdacdyn_cry_4),
            .carryout(un5_sdacdyn_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_6_c_inv_LC_14_10_6.C_ON=1'b1;
    defparam un5_sdacdyn_cry_6_c_inv_LC_14_10_6.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_6_c_inv_LC_14_10_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_sdacdyn_cry_6_c_inv_LC_14_10_6 (
            .in0(N__28934),
            .in1(N__30762),
            .in2(N__28913),
            .in3(_gnd_net_),
            .lcout(sEEACQ_i_6),
            .ltout(),
            .carryin(un5_sdacdyn_cry_5),
            .carryout(un5_sdacdyn_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_7_c_inv_LC_14_10_7.C_ON=1'b1;
    defparam un5_sdacdyn_cry_7_c_inv_LC_14_10_7.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_7_c_inv_LC_14_10_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_sdacdyn_cry_7_c_inv_LC_14_10_7 (
            .in0(N__29378),
            .in1(N__30652),
            .in2(N__29354),
            .in3(_gnd_net_),
            .lcout(sEEACQ_i_7),
            .ltout(),
            .carryin(un5_sdacdyn_cry_6),
            .carryout(un5_sdacdyn_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_8_c_inv_LC_14_11_0.C_ON=1'b1;
    defparam un5_sdacdyn_cry_8_c_inv_LC_14_11_0.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_8_c_inv_LC_14_11_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_8_c_inv_LC_14_11_0 (
            .in0(_gnd_net_),
            .in1(N__30551),
            .in2(N__29324),
            .in3(N__29345),
            .lcout(sEEACQ_i_8),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(un5_sdacdyn_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_9_c_inv_LC_14_11_1.C_ON=1'b1;
    defparam un5_sdacdyn_cry_9_c_inv_LC_14_11_1.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_9_c_inv_LC_14_11_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_9_c_inv_LC_14_11_1 (
            .in0(_gnd_net_),
            .in1(N__30445),
            .in2(N__29291),
            .in3(N__29315),
            .lcout(sEEACQ_i_9),
            .ltout(),
            .carryin(un5_sdacdyn_cry_8),
            .carryout(un5_sdacdyn_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_10_c_inv_LC_14_11_2.C_ON=1'b1;
    defparam un5_sdacdyn_cry_10_c_inv_LC_14_11_2.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_10_c_inv_LC_14_11_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_10_c_inv_LC_14_11_2 (
            .in0(_gnd_net_),
            .in1(N__30337),
            .in2(N__29258),
            .in3(N__29282),
            .lcout(sEEACQ_i_10),
            .ltout(),
            .carryin(un5_sdacdyn_cry_9),
            .carryout(un5_sdacdyn_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_11_c_inv_LC_14_11_3.C_ON=1'b1;
    defparam un5_sdacdyn_cry_11_c_inv_LC_14_11_3.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_11_c_inv_LC_14_11_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_11_c_inv_LC_14_11_3 (
            .in0(_gnd_net_),
            .in1(N__33052),
            .in2(N__29225),
            .in3(N__29249),
            .lcout(sEEACQ_i_11),
            .ltout(),
            .carryin(un5_sdacdyn_cry_10),
            .carryout(un5_sdacdyn_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_12_c_inv_LC_14_11_4.C_ON=1'b1;
    defparam un5_sdacdyn_cry_12_c_inv_LC_14_11_4.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_12_c_inv_LC_14_11_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_12_c_inv_LC_14_11_4 (
            .in0(_gnd_net_),
            .in1(N__31732),
            .in2(N__29195),
            .in3(N__29216),
            .lcout(sEEACQ_i_12),
            .ltout(),
            .carryin(un5_sdacdyn_cry_11),
            .carryout(un5_sdacdyn_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_13_c_inv_LC_14_11_5.C_ON=1'b1;
    defparam un5_sdacdyn_cry_13_c_inv_LC_14_11_5.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_13_c_inv_LC_14_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_13_c_inv_LC_14_11_5 (
            .in0(_gnd_net_),
            .in1(N__31644),
            .in2(N__29165),
            .in3(N__29186),
            .lcout(sEEACQ_i_13),
            .ltout(),
            .carryin(un5_sdacdyn_cry_12),
            .carryout(un5_sdacdyn_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_14_c_inv_LC_14_11_6.C_ON=1'b1;
    defparam un5_sdacdyn_cry_14_c_inv_LC_14_11_6.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_14_c_inv_LC_14_11_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_14_c_inv_LC_14_11_6 (
            .in0(_gnd_net_),
            .in1(N__29132),
            .in2(N__31579),
            .in3(N__29156),
            .lcout(sEEACQ_i_14),
            .ltout(),
            .carryin(un5_sdacdyn_cry_13),
            .carryout(un5_sdacdyn_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_15_c_inv_LC_14_11_7.C_ON=1'b1;
    defparam un5_sdacdyn_cry_15_c_inv_LC_14_11_7.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_15_c_inv_LC_14_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_15_c_inv_LC_14_11_7 (
            .in0(_gnd_net_),
            .in1(N__31454),
            .in2(N__29390),
            .in3(N__29411),
            .lcout(sEEACQ_i_15),
            .ltout(),
            .carryin(un5_sdacdyn_cry_14),
            .carryout(un5_sdacdyn_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_16_c_LC_14_12_0.C_ON=1'b1;
    defparam un5_sdacdyn_cry_16_c_LC_14_12_0.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_16_c_LC_14_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_16_c_LC_14_12_0 (
            .in0(_gnd_net_),
            .in1(N__31389),
            .in2(N__52570),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(un5_sdacdyn_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_17_c_LC_14_12_1.C_ON=1'b1;
    defparam un5_sdacdyn_cry_17_c_LC_14_12_1.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_17_c_LC_14_12_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_17_c_LC_14_12_1 (
            .in0(_gnd_net_),
            .in1(N__52491),
            .in2(N__31284),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_16),
            .carryout(un5_sdacdyn_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_18_c_LC_14_12_2.C_ON=1'b1;
    defparam un5_sdacdyn_cry_18_c_LC_14_12_2.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_18_c_LC_14_12_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_18_c_LC_14_12_2 (
            .in0(_gnd_net_),
            .in1(N__31162),
            .in2(N__52571),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_17),
            .carryout(un5_sdacdyn_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_19_c_LC_14_12_3.C_ON=1'b1;
    defparam un5_sdacdyn_cry_19_c_LC_14_12_3.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_19_c_LC_14_12_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_19_c_LC_14_12_3 (
            .in0(_gnd_net_),
            .in1(N__52495),
            .in2(N__33274),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_18),
            .carryout(un5_sdacdyn_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_20_c_LC_14_12_4.C_ON=1'b1;
    defparam un5_sdacdyn_cry_20_c_LC_14_12_4.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_20_c_LC_14_12_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_20_c_LC_14_12_4 (
            .in0(_gnd_net_),
            .in1(N__33375),
            .in2(N__52572),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_19),
            .carryout(un5_sdacdyn_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_21_c_LC_14_12_5.C_ON=1'b1;
    defparam un5_sdacdyn_cry_21_c_LC_14_12_5.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_21_c_LC_14_12_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_21_c_LC_14_12_5 (
            .in0(_gnd_net_),
            .in1(N__52499),
            .in2(N__33169),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_20),
            .carryout(un5_sdacdyn_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_22_c_LC_14_12_6.C_ON=1'b1;
    defparam un5_sdacdyn_cry_22_c_LC_14_12_6.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_22_c_LC_14_12_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_22_c_LC_14_12_6 (
            .in0(_gnd_net_),
            .in1(N__32037),
            .in2(N__52573),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_21),
            .carryout(un5_sdacdyn_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_23_c_LC_14_12_7.C_ON=1'b1;
    defparam un5_sdacdyn_cry_23_c_LC_14_12_7.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_23_c_LC_14_12_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_23_c_LC_14_12_7 (
            .in0(_gnd_net_),
            .in1(N__52503),
            .in2(N__31936),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_22),
            .carryout(un5_sdacdyn_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_23_c_RNIELG28_LC_14_13_0.C_ON=1'b0;
    defparam un5_sdacdyn_cry_23_c_RNIELG28_LC_14_13_0.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_23_c_RNIELG28_LC_14_13_0.LUT_INIT=16'b0000000011001000;
    LogicCell40 un5_sdacdyn_cry_23_c_RNIELG28_LC_14_13_0 (
            .in0(N__29557),
            .in1(N__36899),
            .in2(N__31052),
            .in3(N__29528),
            .lcout(un5_sdacdyn_cry_23_c_RNIELGZ0Z28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_pointer_0_LC_14_13_1.C_ON=1'b0;
    defparam sDAC_mem_pointer_0_LC_14_13_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_0_LC_14_13_1.LUT_INIT=16'b0011001111111111;
    LogicCell40 sDAC_mem_pointer_0_LC_14_13_1 (
            .in0(_gnd_net_),
            .in1(N__41566),
            .in2(_gnd_net_),
            .in3(N__37584),
            .lcout(sDAC_mem_pointerZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48469),
            .ce(N__43951),
            .sr(N__51678));
    defparam sDAC_data_RNO_30_10_LC_14_13_2.C_ON=1'b0;
    defparam sDAC_data_RNO_30_10_LC_14_13_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_10_LC_14_13_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_30_10_LC_14_13_2 (
            .in0(N__41565),
            .in1(N__42803),
            .in2(_gnd_net_),
            .in3(N__29525),
            .lcout(sDAC_data_RNO_30Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_31_10_LC_14_13_3.C_ON=1'b0;
    defparam sDAC_data_RNO_31_10_LC_14_13_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_10_LC_14_13_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_31_10_LC_14_13_3 (
            .in0(N__29735),
            .in1(N__41564),
            .in2(_gnd_net_),
            .in3(N__29513),
            .lcout(sDAC_data_RNO_31Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_pointer_1_LC_14_13_4.C_ON=1'b0;
    defparam sDAC_mem_pointer_1_LC_14_13_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_1_LC_14_13_4.LUT_INIT=16'b0010001010001000;
    LogicCell40 sDAC_mem_pointer_1_LC_14_13_4 (
            .in0(N__37582),
            .in1(N__38403),
            .in2(_gnd_net_),
            .in3(N__41658),
            .lcout(sDAC_mem_pointerZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48469),
            .ce(N__43951),
            .sr(N__51678));
    defparam sDAC_data_10_LC_14_13_5.C_ON=1'b0;
    defparam sDAC_data_10_LC_14_13_5.SEQ_MODE=4'b1010;
    defparam sDAC_data_10_LC_14_13_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_10_LC_14_13_5 (
            .in0(N__32072),
            .in1(N__37583),
            .in2(_gnd_net_),
            .in3(N__32927),
            .lcout(sDAC_dataZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48469),
            .ce(N__43951),
            .sr(N__51678));
    defparam sDAC_data_RNO_30_5_LC_14_13_6.C_ON=1'b0;
    defparam sDAC_data_RNO_30_5_LC_14_13_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_5_LC_14_13_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_30_5_LC_14_13_6 (
            .in0(N__41563),
            .in1(N__41357),
            .in2(_gnd_net_),
            .in3(N__29480),
            .lcout(sDAC_data_RNO_30Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_30_8_LC_14_13_7.C_ON=1'b0;
    defparam sDAC_data_RNO_30_8_LC_14_13_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_8_LC_14_13_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_30_8_LC_14_13_7 (
            .in0(N__41657),
            .in1(N__41369),
            .in2(_gnd_net_),
            .in3(N__29462),
            .lcout(sDAC_data_RNO_30Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_9_LC_14_14_0.C_ON=1'b0;
    defparam sDAC_data_RNO_23_9_LC_14_14_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_9_LC_14_14_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_9_LC_14_14_0 (
            .in0(N__41861),
            .in1(N__29438),
            .in2(_gnd_net_),
            .in3(N__29714),
            .lcout(sDAC_data_RNO_23Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_28_6_LC_14_14_1.C_ON=1'b0;
    defparam sDAC_mem_28_6_LC_14_14_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_6_LC_14_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_6_LC_14_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50546),
            .lcout(sDAC_mem_28Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52254),
            .ce(N__37807),
            .sr(N__51670));
    defparam sDAC_data_RNO_24_3_LC_14_14_2.C_ON=1'b0;
    defparam sDAC_data_RNO_24_3_LC_14_14_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_3_LC_14_14_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_3_LC_14_14_2 (
            .in0(N__41864),
            .in1(N__29708),
            .in2(_gnd_net_),
            .in3(N__29699),
            .lcout(sDAC_data_RNO_24Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_6_LC_14_14_3.C_ON=1'b0;
    defparam sDAC_data_RNO_24_6_LC_14_14_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_6_LC_14_14_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_6_LC_14_14_3 (
            .in0(N__41720),
            .in1(N__29684),
            .in2(_gnd_net_),
            .in3(N__29675),
            .lcout(sDAC_data_RNO_24Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_9_LC_14_14_4.C_ON=1'b0;
    defparam sDAC_data_RNO_24_9_LC_14_14_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_9_LC_14_14_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_9_LC_14_14_4 (
            .in0(N__41862),
            .in1(N__29663),
            .in2(_gnd_net_),
            .in3(N__29651),
            .lcout(sDAC_data_RNO_24Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_28_3_LC_14_14_5.C_ON=1'b0;
    defparam sDAC_data_RNO_28_3_LC_14_14_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_3_LC_14_14_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_28_3_LC_14_14_5 (
            .in0(N__41721),
            .in1(N__38639),
            .in2(_gnd_net_),
            .in3(N__29624),
            .lcout(sDAC_data_RNO_28Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_28_4_LC_14_14_6.C_ON=1'b0;
    defparam sDAC_data_RNO_28_4_LC_14_14_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_4_LC_14_14_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_28_4_LC_14_14_6 (
            .in0(N__41863),
            .in1(N__38630),
            .in2(_gnd_net_),
            .in3(N__29609),
            .lcout(sDAC_data_RNO_28Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_28_5_LC_14_14_7.C_ON=1'b0;
    defparam sDAC_data_RNO_28_5_LC_14_14_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_5_LC_14_14_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_28_5_LC_14_14_7 (
            .in0(N__41722),
            .in1(N__38621),
            .in2(_gnd_net_),
            .in3(N__29582),
            .lcout(sDAC_data_RNO_28Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_27_0_LC_14_15_0.C_ON=1'b0;
    defparam sDAC_mem_27_0_LC_14_15_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_0_LC_14_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_0_LC_14_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46235),
            .lcout(sDAC_mem_27Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52267),
            .ce(N__29726),
            .sr(N__51663));
    defparam sDAC_mem_27_1_LC_14_15_1.C_ON=1'b0;
    defparam sDAC_mem_27_1_LC_14_15_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_1_LC_14_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_1_LC_14_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51041),
            .lcout(sDAC_mem_27Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52267),
            .ce(N__29726),
            .sr(N__51663));
    defparam sDAC_mem_27_2_LC_14_15_2.C_ON=1'b0;
    defparam sDAC_mem_27_2_LC_14_15_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_2_LC_14_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_2_LC_14_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47343),
            .lcout(sDAC_mem_27Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52267),
            .ce(N__29726),
            .sr(N__51663));
    defparam sDAC_mem_27_3_LC_14_15_3.C_ON=1'b0;
    defparam sDAC_mem_27_3_LC_14_15_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_3_LC_14_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_3_LC_14_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46905),
            .lcout(sDAC_mem_27Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52267),
            .ce(N__29726),
            .sr(N__51663));
    defparam sDAC_mem_27_4_LC_14_15_4.C_ON=1'b0;
    defparam sDAC_mem_27_4_LC_14_15_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_4_LC_14_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_4_LC_14_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45605),
            .lcout(sDAC_mem_27Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52267),
            .ce(N__29726),
            .sr(N__51663));
    defparam sDAC_mem_27_5_LC_14_15_5.C_ON=1'b0;
    defparam sDAC_mem_27_5_LC_14_15_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_5_LC_14_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_5_LC_14_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45119),
            .lcout(sDAC_mem_27Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52267),
            .ce(N__29726),
            .sr(N__51663));
    defparam sDAC_mem_27_6_LC_14_15_6.C_ON=1'b0;
    defparam sDAC_mem_27_6_LC_14_15_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_6_LC_14_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_6_LC_14_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50541),
            .lcout(sDAC_mem_27Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52267),
            .ce(N__29726),
            .sr(N__51663));
    defparam sDAC_mem_27_7_LC_14_15_7.C_ON=1'b0;
    defparam sDAC_mem_27_7_LC_14_15_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_7_LC_14_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_7_LC_14_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50059),
            .lcout(sDAC_mem_27Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52267),
            .ce(N__29726),
            .sr(N__51663));
    defparam sEEPonPoff_0_LC_14_16_0.C_ON=1'b0;
    defparam sEEPonPoff_0_LC_14_16_0.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_0_LC_14_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_0_LC_14_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46234),
            .lcout(sEEPonPoffZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52276),
            .ce(N__33677),
            .sr(N__51657));
    defparam sEEPonPoff_1_LC_14_16_1.C_ON=1'b0;
    defparam sEEPonPoff_1_LC_14_16_1.SEQ_MODE=4'b1011;
    defparam sEEPonPoff_1_LC_14_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_1_LC_14_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51040),
            .lcout(sEEPonPoffZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52276),
            .ce(N__33677),
            .sr(N__51657));
    defparam sEEPonPoff_2_LC_14_16_2.C_ON=1'b0;
    defparam sEEPonPoff_2_LC_14_16_2.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_2_LC_14_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_2_LC_14_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47344),
            .lcout(sEEPonPoffZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52276),
            .ce(N__33677),
            .sr(N__51657));
    defparam sEEPonPoff_3_LC_14_16_3.C_ON=1'b0;
    defparam sEEPonPoff_3_LC_14_16_3.SEQ_MODE=4'b1011;
    defparam sEEPonPoff_3_LC_14_16_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPonPoff_3_LC_14_16_3 (
            .in0(N__46764),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPonPoffZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52276),
            .ce(N__33677),
            .sr(N__51657));
    defparam sEEPonPoff_4_LC_14_16_4.C_ON=1'b0;
    defparam sEEPonPoff_4_LC_14_16_4.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_4_LC_14_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_4_LC_14_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45606),
            .lcout(sEEPonPoffZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52276),
            .ce(N__33677),
            .sr(N__51657));
    defparam sEEPonPoff_5_LC_14_16_5.C_ON=1'b0;
    defparam sEEPonPoff_5_LC_14_16_5.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_5_LC_14_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_5_LC_14_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45114),
            .lcout(sEEPonPoffZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52276),
            .ce(N__33677),
            .sr(N__51657));
    defparam sEEPonPoff_6_LC_14_16_6.C_ON=1'b0;
    defparam sEEPonPoff_6_LC_14_16_6.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_6_LC_14_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_6_LC_14_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50543),
            .lcout(sEEPonPoffZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52276),
            .ce(N__33677),
            .sr(N__51657));
    defparam sEEPonPoff_7_LC_14_16_7.C_ON=1'b0;
    defparam sEEPonPoff_7_LC_14_16_7.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_7_LC_14_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_7_LC_14_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50047),
            .lcout(sEEPonPoffZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52276),
            .ce(N__33677),
            .sr(N__51657));
    defparam un4_spoff_cry_0_c_inv_LC_14_17_0.C_ON=1'b1;
    defparam un4_spoff_cry_0_c_inv_LC_14_17_0.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_0_c_inv_LC_14_17_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_spoff_cry_0_c_inv_LC_14_17_0 (
            .in0(N__30248),
            .in1(N__30143),
            .in2(N__30242),
            .in3(_gnd_net_),
            .lcout(sEEPonPoff_i_0),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(un4_spoff_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_1_c_inv_LC_14_17_1.C_ON=1'b1;
    defparam un4_spoff_cry_1_c_inv_LC_14_17_1.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_1_c_inv_LC_14_17_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_spoff_cry_1_c_inv_LC_14_17_1 (
            .in0(_gnd_net_),
            .in1(N__30026),
            .in2(N__30137),
            .in3(N__30032),
            .lcout(sEEPonPoff_i_1),
            .ltout(),
            .carryin(un4_spoff_cry_0),
            .carryout(un4_spoff_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_2_c_inv_LC_14_17_2.C_ON=1'b1;
    defparam un4_spoff_cry_2_c_inv_LC_14_17_2.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_2_c_inv_LC_14_17_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_spoff_cry_2_c_inv_LC_14_17_2 (
            .in0(N__30020),
            .in1(N__29897),
            .in2(N__30014),
            .in3(_gnd_net_),
            .lcout(sEEPonPoff_i_2),
            .ltout(),
            .carryin(un4_spoff_cry_1),
            .carryout(un4_spoff_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_3_c_inv_LC_14_17_3.C_ON=1'b1;
    defparam un4_spoff_cry_3_c_inv_LC_14_17_3.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_3_c_inv_LC_14_17_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_spoff_cry_3_c_inv_LC_14_17_3 (
            .in0(N__29891),
            .in1(N__29783),
            .in2(N__29884),
            .in3(_gnd_net_),
            .lcout(sEEPonPoff_i_3),
            .ltout(),
            .carryin(un4_spoff_cry_2),
            .carryout(un4_spoff_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_4_c_inv_LC_14_17_4.C_ON=1'b1;
    defparam un4_spoff_cry_4_c_inv_LC_14_17_4.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_4_c_inv_LC_14_17_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_spoff_cry_4_c_inv_LC_14_17_4 (
            .in0(N__31067),
            .in1(N__30920),
            .in2(N__31060),
            .in3(_gnd_net_),
            .lcout(sEEPonPoff_i_4),
            .ltout(),
            .carryin(un4_spoff_cry_3),
            .carryout(un4_spoff_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_5_c_inv_LC_14_17_5.C_ON=1'b1;
    defparam un4_spoff_cry_5_c_inv_LC_14_17_5.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_5_c_inv_LC_14_17_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_spoff_cry_5_c_inv_LC_14_17_5 (
            .in0(N__30914),
            .in1(N__30803),
            .in2(N__30908),
            .in3(_gnd_net_),
            .lcout(sEEPonPoff_i_5),
            .ltout(),
            .carryin(un4_spoff_cry_4),
            .carryout(un4_spoff_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_6_c_inv_LC_14_17_6.C_ON=1'b1;
    defparam un4_spoff_cry_6_c_inv_LC_14_17_6.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_6_c_inv_LC_14_17_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_spoff_cry_6_c_inv_LC_14_17_6 (
            .in0(N__30797),
            .in1(N__30692),
            .in2(N__30791),
            .in3(_gnd_net_),
            .lcout(sEEPonPoff_i_6),
            .ltout(),
            .carryin(un4_spoff_cry_5),
            .carryout(un4_spoff_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_7_c_inv_LC_14_17_7.C_ON=1'b1;
    defparam un4_spoff_cry_7_c_inv_LC_14_17_7.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_7_c_inv_LC_14_17_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_spoff_cry_7_c_inv_LC_14_17_7 (
            .in0(_gnd_net_),
            .in1(N__30581),
            .in2(N__30686),
            .in3(N__30587),
            .lcout(sEEPonPoff_i_7),
            .ltout(),
            .carryin(un4_spoff_cry_6),
            .carryout(un4_spoff_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_8_c_LC_14_18_0.C_ON=1'b1;
    defparam un4_spoff_cry_8_c_LC_14_18_0.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_8_c_LC_14_18_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_8_c_LC_14_18_0 (
            .in0(_gnd_net_),
            .in1(N__30571),
            .in2(N__52671),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(un4_spoff_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_9_c_LC_14_18_1.C_ON=1'b1;
    defparam un4_spoff_cry_9_c_LC_14_18_1.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_9_c_LC_14_18_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_9_c_LC_14_18_1 (
            .in0(_gnd_net_),
            .in1(N__52602),
            .in2(N__30470),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_8),
            .carryout(un4_spoff_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_10_c_LC_14_18_2.C_ON=1'b1;
    defparam un4_spoff_cry_10_c_LC_14_18_2.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_10_c_LC_14_18_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_10_c_LC_14_18_2 (
            .in0(_gnd_net_),
            .in1(N__30360),
            .in2(N__52668),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_9),
            .carryout(un4_spoff_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_11_c_LC_14_18_3.C_ON=1'b1;
    defparam un4_spoff_cry_11_c_LC_14_18_3.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_11_c_LC_14_18_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_11_c_LC_14_18_3 (
            .in0(_gnd_net_),
            .in1(N__52590),
            .in2(N__33062),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_10),
            .carryout(un4_spoff_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_12_c_LC_14_18_4.C_ON=1'b1;
    defparam un4_spoff_cry_12_c_LC_14_18_4.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_12_c_LC_14_18_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_12_c_LC_14_18_4 (
            .in0(_gnd_net_),
            .in1(N__31747),
            .in2(N__52669),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_11),
            .carryout(un4_spoff_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_13_c_LC_14_18_5.C_ON=1'b1;
    defparam un4_spoff_cry_13_c_LC_14_18_5.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_13_c_LC_14_18_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_13_c_LC_14_18_5 (
            .in0(_gnd_net_),
            .in1(N__52594),
            .in2(N__31664),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_12),
            .carryout(un4_spoff_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_14_c_LC_14_18_6.C_ON=1'b1;
    defparam un4_spoff_cry_14_c_LC_14_18_6.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_14_c_LC_14_18_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_14_c_LC_14_18_6 (
            .in0(_gnd_net_),
            .in1(N__31578),
            .in2(N__52670),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_13),
            .carryout(un4_spoff_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_15_c_LC_14_18_7.C_ON=1'b1;
    defparam un4_spoff_cry_15_c_LC_14_18_7.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_15_c_LC_14_18_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_15_c_LC_14_18_7 (
            .in0(_gnd_net_),
            .in1(N__52598),
            .in2(N__31484),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_14),
            .carryout(un4_spoff_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_16_c_LC_14_19_0.C_ON=1'b1;
    defparam un4_spoff_cry_16_c_LC_14_19_0.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_16_c_LC_14_19_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_16_c_LC_14_19_0 (
            .in0(_gnd_net_),
            .in1(N__52536),
            .in2(N__31397),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(un4_spoff_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_17_c_LC_14_19_1.C_ON=1'b1;
    defparam un4_spoff_cry_17_c_LC_14_19_1.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_17_c_LC_14_19_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_17_c_LC_14_19_1 (
            .in0(_gnd_net_),
            .in1(N__31283),
            .in2(N__52623),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_16),
            .carryout(un4_spoff_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_18_c_LC_14_19_2.C_ON=1'b1;
    defparam un4_spoff_cry_18_c_LC_14_19_2.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_18_c_LC_14_19_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_18_c_LC_14_19_2 (
            .in0(_gnd_net_),
            .in1(N__52540),
            .in2(N__31176),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_17),
            .carryout(un4_spoff_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_19_c_LC_14_19_3.C_ON=1'b1;
    defparam un4_spoff_cry_19_c_LC_14_19_3.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_19_c_LC_14_19_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_19_c_LC_14_19_3 (
            .in0(_gnd_net_),
            .in1(N__33273),
            .in2(N__52624),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_18),
            .carryout(un4_spoff_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_20_c_LC_14_19_4.C_ON=1'b1;
    defparam un4_spoff_cry_20_c_LC_14_19_4.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_20_c_LC_14_19_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_20_c_LC_14_19_4 (
            .in0(_gnd_net_),
            .in1(N__52544),
            .in2(N__33388),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_19),
            .carryout(un4_spoff_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_21_c_LC_14_19_5.C_ON=1'b1;
    defparam un4_spoff_cry_21_c_LC_14_19_5.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_21_c_LC_14_19_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_21_c_LC_14_19_5 (
            .in0(_gnd_net_),
            .in1(N__33167),
            .in2(N__52625),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_20),
            .carryout(un4_spoff_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_22_c_LC_14_19_6.C_ON=1'b1;
    defparam un4_spoff_cry_22_c_LC_14_19_6.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_22_c_LC_14_19_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_22_c_LC_14_19_6 (
            .in0(_gnd_net_),
            .in1(N__52548),
            .in2(N__32048),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_21),
            .carryout(un4_spoff_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_23_c_LC_14_19_7.C_ON=1'b1;
    defparam un4_spoff_cry_23_c_LC_14_19_7.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_23_c_LC_14_19_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_23_c_LC_14_19_7 (
            .in0(_gnd_net_),
            .in1(N__31929),
            .in2(N__52626),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_22),
            .carryout(un4_spoff_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_23_THRU_LUT4_0_LC_14_20_0.C_ON=1'b0;
    defparam un4_spoff_cry_23_THRU_LUT4_0_LC_14_20_0.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_23_THRU_LUT4_0_LC_14_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un4_spoff_cry_23_THRU_LUT4_0_LC_14_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31820),
            .lcout(un4_spoff_cry_23_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.data_in_3_LC_15_3_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_3_LC_15_3_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_3_LC_15_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_3_LC_15_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37526),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48446),
            .ce(N__43903),
            .sr(N__51796));
    defparam \spi_master_inst.spi_data_path_u1.data_in_4_LC_15_3_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_4_LC_15_3_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_4_LC_15_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_4_LC_15_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31793),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48446),
            .ce(N__43903),
            .sr(N__51796));
    defparam \spi_master_inst.spi_data_path_u1.data_in_7_LC_15_3_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_7_LC_15_3_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_7_LC_15_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_7_LC_15_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32132),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48446),
            .ce(N__43903),
            .sr(N__51796));
    defparam \spi_master_inst.spi_data_path_u1.data_in_8_LC_15_3_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_8_LC_15_3_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_8_LC_15_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_8_LC_15_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31760),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48446),
            .ce(N__43903),
            .sr(N__51796));
    defparam \spi_master_inst.spi_data_path_u1.data_in_9_LC_15_3_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_9_LC_15_3_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_9_LC_15_3_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_9_LC_15_3_7  (
            .in0(N__32288),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48446),
            .ce(N__43903),
            .sr(N__51796));
    defparam sEEDAC_0_LC_15_4_0.C_ON=1'b0;
    defparam sEEDAC_0_LC_15_4_0.SEQ_MODE=4'b1000;
    defparam sEEDAC_0_LC_15_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_0_LC_15_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46233),
            .lcout(sEEDACZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52289),
            .ce(N__32057),
            .sr(_gnd_net_));
    defparam sEEDAC_1_LC_15_4_1.C_ON=1'b0;
    defparam sEEDAC_1_LC_15_4_1.SEQ_MODE=4'b1000;
    defparam sEEDAC_1_LC_15_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_1_LC_15_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50982),
            .lcout(sEEDACZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52289),
            .ce(N__32057),
            .sr(_gnd_net_));
    defparam sEEDAC_2_LC_15_4_2.C_ON=1'b0;
    defparam sEEDAC_2_LC_15_4_2.SEQ_MODE=4'b1000;
    defparam sEEDAC_2_LC_15_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_2_LC_15_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47347),
            .lcout(sEEDACZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52289),
            .ce(N__32057),
            .sr(_gnd_net_));
    defparam sEEDAC_3_LC_15_4_3.C_ON=1'b0;
    defparam sEEDAC_3_LC_15_4_3.SEQ_MODE=4'b1000;
    defparam sEEDAC_3_LC_15_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_3_LC_15_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46750),
            .lcout(sEEDACZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52289),
            .ce(N__32057),
            .sr(_gnd_net_));
    defparam sEEDAC_4_LC_15_4_4.C_ON=1'b0;
    defparam sEEDAC_4_LC_15_4_4.SEQ_MODE=4'b1000;
    defparam sEEDAC_4_LC_15_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_4_LC_15_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45506),
            .lcout(sEEDACZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52289),
            .ce(N__32057),
            .sr(_gnd_net_));
    defparam sEEDAC_5_LC_15_4_5.C_ON=1'b0;
    defparam sEEDAC_5_LC_15_4_5.SEQ_MODE=4'b1000;
    defparam sEEDAC_5_LC_15_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_5_LC_15_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44980),
            .lcout(sEEDACZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52289),
            .ce(N__32057),
            .sr(_gnd_net_));
    defparam sEEDAC_6_LC_15_4_6.C_ON=1'b0;
    defparam sEEDAC_6_LC_15_4_6.SEQ_MODE=4'b1000;
    defparam sEEDAC_6_LC_15_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_6_LC_15_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50409),
            .lcout(sEEDACZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52289),
            .ce(N__32057),
            .sr(_gnd_net_));
    defparam sEEDAC_7_LC_15_4_7.C_ON=1'b0;
    defparam sEEDAC_7_LC_15_4_7.SEQ_MODE=4'b1000;
    defparam sEEDAC_7_LC_15_4_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEDAC_7_LC_15_4_7 (
            .in0(N__50052),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEDACZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52289),
            .ce(N__32057),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_7_LC_15_5_0.C_ON=1'b0;
    defparam sDAC_data_RNO_10_7_LC_15_5_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_7_LC_15_5_0.LUT_INIT=16'b1010000011001111;
    LogicCell40 sDAC_data_RNO_10_7_LC_15_5_0 (
            .in0(N__34385),
            .in1(N__33602),
            .in2(N__38258),
            .in3(N__32189),
            .lcout(sDAC_data_RNO_10Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_7_LC_15_5_1.C_ON=1'b0;
    defparam sDAC_data_RNO_22_7_LC_15_5_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_7_LC_15_5_1.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_22_7_LC_15_5_1 (
            .in0(N__38508),
            .in1(N__32204),
            .in2(N__38200),
            .in3(N__32198),
            .lcout(sDAC_data_2_32_ns_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_7_LC_15_5_2.C_ON=1'b0;
    defparam sDAC_data_RNO_6_7_LC_15_5_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_7_LC_15_5_2.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_6_7_LC_15_5_2 (
            .in0(N__38509),
            .in1(N__34187),
            .in2(N__38257),
            .in3(N__36881),
            .lcout(),
            .ltout(sDAC_data_2_14_ns_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_7_LC_15_5_3.C_ON=1'b0;
    defparam sDAC_data_RNO_1_7_LC_15_5_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_7_LC_15_5_3.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_1_7_LC_15_5_3 (
            .in0(N__32327),
            .in1(N__38230),
            .in2(N__32183),
            .in3(N__32180),
            .lcout(sDAC_data_RNO_1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_7_LC_15_5_4.C_ON=1'b0;
    defparam sDAC_data_RNO_3_7_LC_15_5_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_7_LC_15_5_4.LUT_INIT=16'b0010010101110101;
    LogicCell40 sDAC_data_RNO_3_7_LC_15_5_4 (
            .in0(N__37342),
            .in1(N__32174),
            .in2(N__37487),
            .in3(N__32159),
            .lcout(),
            .ltout(sDAC_data_2_41_ns_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_7_LC_15_5_5.C_ON=1'b0;
    defparam sDAC_data_RNO_0_7_LC_15_5_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_7_LC_15_5_5.LUT_INIT=16'b0011111000001110;
    LogicCell40 sDAC_data_RNO_0_7_LC_15_5_5 (
            .in0(N__34142),
            .in1(N__37485),
            .in2(N__32153),
            .in3(N__32150),
            .lcout(),
            .ltout(sDAC_data_2_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_7_LC_15_5_6.C_ON=1'b0;
    defparam sDAC_data_7_LC_15_5_6.SEQ_MODE=4'b1010;
    defparam sDAC_data_7_LC_15_5_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 sDAC_data_7_LC_15_5_6 (
            .in0(N__32144),
            .in1(_gnd_net_),
            .in2(N__32135),
            .in3(N__37637),
            .lcout(sDAC_dataZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48453),
            .ce(N__43954),
            .sr(N__51770));
    defparam sDAC_data_RNO_1_9_LC_15_6_0.C_ON=1'b0;
    defparam sDAC_data_RNO_1_9_LC_15_6_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_9_LC_15_6_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_1_9_LC_15_6_0 (
            .in0(N__32453),
            .in1(N__32684),
            .in2(N__38256),
            .in3(N__32279),
            .lcout(),
            .ltout(sDAC_data_RNO_1Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_9_LC_15_6_1.C_ON=1'b0;
    defparam sDAC_data_RNO_0_9_LC_15_6_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_9_LC_15_6_1.LUT_INIT=16'b0101000011101110;
    LogicCell40 sDAC_data_RNO_0_9_LC_15_6_1 (
            .in0(N__37486),
            .in1(N__34253),
            .in2(N__32123),
            .in3(N__32237),
            .lcout(),
            .ltout(sDAC_data_2_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_9_LC_15_6_2.C_ON=1'b0;
    defparam sDAC_data_9_LC_15_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_data_9_LC_15_6_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 sDAC_data_9_LC_15_6_2 (
            .in0(N__32300),
            .in1(_gnd_net_),
            .in2(N__32291),
            .in3(N__37630),
            .lcout(sDAC_dataZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48456),
            .ce(N__43952),
            .sr(N__51757));
    defparam sDAC_data_RNO_6_9_LC_15_6_3.C_ON=1'b0;
    defparam sDAC_data_RNO_6_9_LC_15_6_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_9_LC_15_6_3.LUT_INIT=16'b0011010000110111;
    LogicCell40 sDAC_data_RNO_6_9_LC_15_6_3 (
            .in0(N__34337),
            .in1(N__38533),
            .in2(N__38201),
            .in3(N__34460),
            .lcout(sDAC_data_2_14_ns_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_9_LC_15_6_4.C_ON=1'b0;
    defparam sDAC_data_RNO_22_9_LC_15_6_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_9_LC_15_6_4.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_22_9_LC_15_6_4 (
            .in0(N__38532),
            .in1(N__32273),
            .in2(N__38255),
            .in3(N__32264),
            .lcout(),
            .ltout(sDAC_data_2_32_ns_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_9_LC_15_6_5.C_ON=1'b0;
    defparam sDAC_data_RNO_10_9_LC_15_6_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_9_LC_15_6_5.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_10_9_LC_15_6_5 (
            .in0(N__38104),
            .in1(N__33560),
            .in2(N__32258),
            .in3(N__32216),
            .lcout(),
            .ltout(sDAC_data_RNO_10Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_9_LC_15_6_6.C_ON=1'b0;
    defparam sDAC_data_RNO_3_9_LC_15_6_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_9_LC_15_6_6.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_3_9_LC_15_6_6 (
            .in0(N__37462),
            .in1(N__37341),
            .in2(N__32255),
            .in3(N__32252),
            .lcout(sDAC_data_2_41_ns_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_20_8_LC_15_7_0.C_ON=1'b0;
    defparam sDAC_data_RNO_20_8_LC_15_7_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_8_LC_15_7_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_20_8_LC_15_7_0 (
            .in0(N__34067),
            .in1(N__42146),
            .in2(_gnd_net_),
            .in3(N__32222),
            .lcout(sDAC_data_RNO_20Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_20_5_LC_15_7_1.C_ON=1'b0;
    defparam sDAC_mem_20_5_LC_15_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_5_LC_15_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_5_LC_15_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45068),
            .lcout(sDAC_mem_20Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52255),
            .ce(N__36637),
            .sr(N__51745));
    defparam sDAC_data_RNO_20_9_LC_15_7_2.C_ON=1'b0;
    defparam sDAC_data_RNO_20_9_LC_15_7_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_9_LC_15_7_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_20_9_LC_15_7_2 (
            .in0(N__42114),
            .in1(N__34058),
            .in2(_gnd_net_),
            .in3(N__32210),
            .lcout(sDAC_data_RNO_20Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_20_6_LC_15_7_3.C_ON=1'b0;
    defparam sDAC_mem_20_6_LC_15_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_6_LC_15_7_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_20_6_LC_15_7_3 (
            .in0(N__50469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_20Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52255),
            .ce(N__36637),
            .sr(N__51745));
    defparam sDAC_data_RNO_21_3_LC_15_7_4.C_ON=1'b0;
    defparam sDAC_data_RNO_21_3_LC_15_7_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_3_LC_15_7_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_3_LC_15_7_4 (
            .in0(N__42112),
            .in1(N__36515),
            .in2(_gnd_net_),
            .in3(N__32408),
            .lcout(sDAC_data_RNO_21Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_21_4_LC_15_7_5.C_ON=1'b0;
    defparam sDAC_data_RNO_21_4_LC_15_7_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_4_LC_15_7_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_4_LC_15_7_5 (
            .in0(N__42147),
            .in1(N__36503),
            .in2(_gnd_net_),
            .in3(N__32396),
            .lcout(sDAC_data_RNO_21Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_21_5_LC_15_7_6.C_ON=1'b0;
    defparam sDAC_data_RNO_21_5_LC_15_7_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_5_LC_15_7_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_5_LC_15_7_6 (
            .in0(N__42113),
            .in1(N__36491),
            .in2(_gnd_net_),
            .in3(N__32378),
            .lcout(sDAC_data_RNO_21Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_21_6_LC_15_7_7.C_ON=1'b0;
    defparam sDAC_data_RNO_21_6_LC_15_7_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_6_LC_15_7_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_6_LC_15_7_7 (
            .in0(N__42145),
            .in1(N__36776),
            .in2(_gnd_net_),
            .in3(N__32366),
            .lcout(sDAC_data_RNO_21Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_4_3_LC_15_8_2.C_ON=1'b0;
    defparam sDAC_mem_4_3_LC_15_8_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_3_LC_15_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_3_LC_15_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46779),
            .lcout(sDAC_mem_4Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52245),
            .ce(N__42640),
            .sr(N__51730));
    defparam sDAC_data_RNO_12_7_LC_15_8_3.C_ON=1'b0;
    defparam sDAC_data_RNO_12_7_LC_15_8_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_7_LC_15_8_3.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_12_7_LC_15_8_3 (
            .in0(N__42426),
            .in1(N__32342),
            .in2(N__42248),
            .in3(N__32318),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_7_LC_15_8_4.C_ON=1'b0;
    defparam sDAC_data_RNO_4_7_LC_15_8_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_7_LC_15_8_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_7_LC_15_8_4 (
            .in0(N__42211),
            .in1(N__41123),
            .in2(N__32330),
            .in3(N__44483),
            .lcout(sDAC_data_RNO_4Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_4_4_LC_15_8_5.C_ON=1'b0;
    defparam sDAC_mem_4_4_LC_15_8_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_4_LC_15_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_4_LC_15_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45509),
            .lcout(sDAC_mem_4Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52245),
            .ce(N__42640),
            .sr(N__51730));
    defparam sDAC_data_RNO_12_8_LC_15_8_6.C_ON=1'b0;
    defparam sDAC_data_RNO_12_8_LC_15_8_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_8_LC_15_8_6.LUT_INIT=16'b0101010100100111;
    LogicCell40 sDAC_data_RNO_12_8_LC_15_8_6 (
            .in0(N__42432),
            .in1(N__32312),
            .in2(N__36479),
            .in3(N__42209),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_8_LC_15_8_7.C_ON=1'b0;
    defparam sDAC_data_RNO_4_8_LC_15_8_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_8_LC_15_8_7.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_8_LC_15_8_7 (
            .in0(N__42210),
            .in1(N__41111),
            .in2(N__32552),
            .in3(N__44471),
            .lcout(sDAC_data_RNO_4Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_13_8_LC_15_9_0.C_ON=1'b0;
    defparam sDAC_data_RNO_13_8_LC_15_9_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_8_LC_15_9_0.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_13_8_LC_15_9_0 (
            .in0(N__42425),
            .in1(N__32537),
            .in2(N__42213),
            .in3(N__32486),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_8_LC_15_9_1.C_ON=1'b0;
    defparam sDAC_data_RNO_5_8_LC_15_9_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_8_LC_15_9_1.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_5_8_LC_15_9_1 (
            .in0(N__42149),
            .in1(N__32522),
            .in2(N__32513),
            .in3(N__32510),
            .lcout(sDAC_data_RNO_5Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_6_5_LC_15_9_2.C_ON=1'b0;
    defparam sDAC_mem_6_5_LC_15_9_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_5_LC_15_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_5_LC_15_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45067),
            .lcout(sDAC_mem_6Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52234),
            .ce(N__36553),
            .sr(N__51718));
    defparam sDAC_data_RNO_13_9_LC_15_9_3.C_ON=1'b0;
    defparam sDAC_data_RNO_13_9_LC_15_9_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_9_LC_15_9_3.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_13_9_LC_15_9_3 (
            .in0(N__42525),
            .in1(N__32480),
            .in2(N__42238),
            .in3(N__32444),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_9_LC_15_9_4.C_ON=1'b0;
    defparam sDAC_data_RNO_5_9_LC_15_9_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_9_LC_15_9_4.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_5_9_LC_15_9_4 (
            .in0(N__44297),
            .in1(N__42153),
            .in2(N__32465),
            .in3(N__32462),
            .lcout(sDAC_data_RNO_5Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_6_6_LC_15_9_5.C_ON=1'b0;
    defparam sDAC_mem_6_6_LC_15_9_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_6_LC_15_9_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_6_6_LC_15_9_5 (
            .in0(N__50463),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_6Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52234),
            .ce(N__36553),
            .sr(N__51718));
    defparam sDAC_data_RNO_16_10_LC_15_9_6.C_ON=1'b0;
    defparam sDAC_data_RNO_16_10_LC_15_9_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_10_LC_15_9_6.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_16_10_LC_15_9_6 (
            .in0(N__42424),
            .in1(N__32438),
            .in2(N__42212),
            .in3(N__32423),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_10_LC_15_9_7.C_ON=1'b0;
    defparam sDAC_data_RNO_7_10_LC_15_9_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_10_LC_15_9_7.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_7_10_LC_15_9_7 (
            .in0(N__42148),
            .in1(N__39830),
            .in2(N__32702),
            .in3(N__37028),
            .lcout(sDAC_data_RNO_7Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_12_9_LC_15_10_0.C_ON=1'b0;
    defparam sDAC_data_RNO_12_9_LC_15_10_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_9_LC_15_10_0.LUT_INIT=16'b0101010100100111;
    LogicCell40 sDAC_data_RNO_12_9_LC_15_10_0 (
            .in0(N__42576),
            .in1(N__32699),
            .in2(N__32672),
            .in3(N__42000),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_9_LC_15_10_1.C_ON=1'b0;
    defparam sDAC_data_RNO_4_9_LC_15_10_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_9_LC_15_10_1.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_4_9_LC_15_10_1 (
            .in0(N__44459),
            .in1(N__41988),
            .in2(N__32687),
            .in3(N__41099),
            .lcout(sDAC_data_RNO_4Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_4_6_LC_15_10_2.C_ON=1'b0;
    defparam sDAC_mem_4_6_LC_15_10_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_6_LC_15_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_6_LC_15_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50516),
            .lcout(sDAC_mem_4Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52224),
            .ce(N__42636),
            .sr(N__51707));
    defparam sDAC_data_RNO_13_10_LC_15_10_3.C_ON=1'b0;
    defparam sDAC_data_RNO_13_10_LC_15_10_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_10_LC_15_10_3.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_13_10_LC_15_10_3 (
            .in0(N__42511),
            .in1(N__32663),
            .in2(N__42172),
            .in3(N__36569),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_10_LC_15_10_4.C_ON=1'b0;
    defparam sDAC_data_RNO_5_10_LC_15_10_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_10_LC_15_10_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_5_10_LC_15_10_4 (
            .in0(N__41986),
            .in1(N__32648),
            .in2(N__32636),
            .in3(N__32633),
            .lcout(sDAC_data_RNO_5Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_13_3_LC_15_10_5.C_ON=1'b0;
    defparam sDAC_data_RNO_13_3_LC_15_10_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_3_LC_15_10_5.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_13_3_LC_15_10_5 (
            .in0(N__42512),
            .in1(N__32621),
            .in2(N__42173),
            .in3(N__36611),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_3_LC_15_10_6.C_ON=1'b0;
    defparam sDAC_data_RNO_5_3_LC_15_10_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_3_LC_15_10_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_5_3_LC_15_10_6 (
            .in0(N__41987),
            .in1(N__32606),
            .in2(N__32594),
            .in3(N__32591),
            .lcout(sDAC_data_RNO_5Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_13_4_LC_15_10_7.C_ON=1'b0;
    defparam sDAC_data_RNO_13_4_LC_15_10_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_4_LC_15_10_7.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_13_4_LC_15_10_7 (
            .in0(N__42510),
            .in1(N__32579),
            .in2(N__42171),
            .in3(N__36596),
            .lcout(sDAC_data_2_13_bm_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_27_10_LC_15_11_0.C_ON=1'b0;
    defparam sDAC_data_RNO_27_10_LC_15_11_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_10_LC_15_11_0.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_27_10_LC_15_11_0 (
            .in0(N__42515),
            .in1(N__32873),
            .in2(N__42097),
            .in3(N__32861),
            .lcout(sDAC_data_2_6_bm_1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_2_7_LC_15_11_1.C_ON=1'b0;
    defparam sDAC_mem_2_7_LC_15_11_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_7_LC_15_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_7_LC_15_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50009),
            .lcout(sDAC_mem_2Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52218),
            .ce(N__32855),
            .sr(N__51699));
    defparam sDAC_data_RNO_18_10_LC_15_11_2.C_ON=1'b0;
    defparam sDAC_data_RNO_18_10_LC_15_11_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_10_LC_15_11_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_10_LC_15_11_2 (
            .in0(N__41891),
            .in1(N__44597),
            .in2(_gnd_net_),
            .in3(N__32828),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_10_LC_15_11_3.C_ON=1'b0;
    defparam sDAC_data_RNO_9_10_LC_15_11_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_10_LC_15_11_3.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_9_10_LC_15_11_3 (
            .in0(N__38166),
            .in1(N__38500),
            .in2(N__32813),
            .in3(N__32780),
            .lcout(sDAC_data_2_24_ns_1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_19_10_LC_15_11_4.C_ON=1'b0;
    defparam sDAC_data_RNO_19_10_LC_15_11_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_10_LC_15_11_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_10_LC_15_11_4 (
            .in0(N__41887),
            .in1(N__32810),
            .in2(_gnd_net_),
            .in3(N__32795),
            .lcout(sDAC_data_RNO_19Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_10_LC_15_11_5.C_ON=1'b0;
    defparam sDAC_data_RNO_17_10_LC_15_11_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_10_LC_15_11_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_10_LC_15_11_5 (
            .in0(N__42521),
            .in1(N__32774),
            .in2(_gnd_net_),
            .in3(N__32759),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_10_LC_15_11_6.C_ON=1'b0;
    defparam sDAC_data_RNO_8_10_LC_15_11_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_10_LC_15_11_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 sDAC_data_RNO_8_10_LC_15_11_6 (
            .in0(N__41892),
            .in1(_gnd_net_),
            .in2(N__32741),
            .in3(N__32738),
            .lcout(),
            .ltout(sDAC_data_RNO_8Z0Z_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_10_LC_15_11_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_10_LC_15_11_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_10_LC_15_11_7.LUT_INIT=16'b0111011000110010;
    LogicCell40 sDAC_data_RNO_2_10_LC_15_11_7 (
            .in0(N__38167),
            .in1(N__32720),
            .in2(N__32714),
            .in3(N__32711),
            .lcout(sDAC_data_RNO_2Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam button_debounce_counter_esr_RNO_0_23_LC_15_12_0.C_ON=1'b0;
    defparam button_debounce_counter_esr_RNO_0_23_LC_15_12_0.SEQ_MODE=4'b0000;
    defparam button_debounce_counter_esr_RNO_0_23_LC_15_12_0.LUT_INIT=16'b1111111110101010;
    LogicCell40 button_debounce_counter_esr_RNO_0_23_LC_15_12_0 (
            .in0(N__45722),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49427),
            .lcout(LED3_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNITC6L_19_LC_15_12_1.C_ON=1'b0;
    defparam sCounter_RNITC6L_19_LC_15_12_1.SEQ_MODE=4'b0000;
    defparam sCounter_RNITC6L_19_LC_15_12_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNITC6L_19_LC_15_12_1 (
            .in0(N__33374),
            .in1(N__33257),
            .in2(N__33168),
            .in3(N__33047),
            .lcout(g0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.spi_cs_i_LC_15_12_2 .C_ON=1'b0;
    defparam \spi_slave_inst.spi_cs_i_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.spi_cs_i_LC_15_12_2 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \spi_slave_inst.spi_cs_i_LC_15_12_2  (
            .in0(N__47903),
            .in1(N__48041),
            .in2(_gnd_net_),
            .in3(N__47947),
            .lcout(\spi_slave_inst.spi_cs_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_10_LC_15_12_4.C_ON=1'b0;
    defparam sDAC_data_RNO_3_10_LC_15_12_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_10_LC_15_12_4.LUT_INIT=16'b0001010110110101;
    LogicCell40 sDAC_data_RNO_3_10_LC_15_12_4 (
            .in0(N__37343),
            .in1(N__32879),
            .in2(N__37481),
            .in3(N__33404),
            .lcout(),
            .ltout(sDAC_data_2_41_ns_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_10_LC_15_12_5.C_ON=1'b0;
    defparam sDAC_data_RNO_0_10_LC_15_12_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_10_LC_15_12_5.LUT_INIT=16'b0011111000001110;
    LogicCell40 sDAC_data_RNO_0_10_LC_15_12_5 (
            .in0(N__32936),
            .in1(N__37471),
            .in2(N__32930),
            .in3(N__34943),
            .lcout(sDAC_data_2_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_0_LC_15_12_6.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_0_LC_15_12_6.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_0_LC_15_12_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_0_LC_15_12_6 (
            .in0(N__35072),
            .in1(N__35039),
            .in2(N__35057),
            .in3(N__35087),
            .lcout(sbuttonModeStatus_0_sqmuxa_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_21_10_LC_15_13_0.C_ON=1'b0;
    defparam sDAC_data_RNO_21_10_LC_15_13_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_10_LC_15_13_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_10_LC_15_13_0 (
            .in0(N__41804),
            .in1(N__36716),
            .in2(_gnd_net_),
            .in3(N__32909),
            .lcout(sDAC_data_RNO_21Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_28_10_LC_15_13_1.C_ON=1'b0;
    defparam sDAC_data_RNO_28_10_LC_15_13_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_10_LC_15_13_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_28_10_LC_15_13_1 (
            .in0(N__41807),
            .in1(N__38963),
            .in2(_gnd_net_),
            .in3(N__33518),
            .lcout(),
            .ltout(sDAC_data_RNO_28Z0Z_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_10_LC_15_13_2.C_ON=1'b0;
    defparam sDAC_data_RNO_22_10_LC_15_13_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_10_LC_15_13_2.LUT_INIT=16'b0100010101100111;
    LogicCell40 sDAC_data_RNO_22_10_LC_15_13_2 (
            .in0(N__38452),
            .in1(N__38115),
            .in2(N__32891),
            .in3(N__33524),
            .lcout(),
            .ltout(sDAC_data_2_32_ns_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_10_LC_15_13_3.C_ON=1'b0;
    defparam sDAC_data_RNO_10_10_LC_15_13_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_10_LC_15_13_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_10_10_LC_15_13_3 (
            .in0(N__38116),
            .in1(N__32888),
            .in2(N__32882),
            .in3(N__33548),
            .lcout(sDAC_data_RNO_10Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_20_10_LC_15_13_4.C_ON=1'b0;
    defparam sDAC_data_RNO_20_10_LC_15_13_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_10_LC_15_13_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_20_10_LC_15_13_4 (
            .in0(N__41805),
            .in1(N__34046),
            .in2(_gnd_net_),
            .in3(N__36653),
            .lcout(sDAC_data_RNO_20Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_29_10_LC_15_13_5.C_ON=1'b0;
    defparam sDAC_data_RNO_29_10_LC_15_13_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_10_LC_15_13_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 sDAC_data_RNO_29_10_LC_15_13_5 (
            .in0(_gnd_net_),
            .in1(N__34079),
            .in2(N__33542),
            .in3(N__41806),
            .lcout(sDAC_data_RNO_29Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_16_7_LC_15_13_6.C_ON=1'b0;
    defparam sDAC_mem_16_7_LC_15_13_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_7_LC_15_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_7_LC_15_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50056),
            .lcout(sDAC_mem_16Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52235),
            .ce(N__33512),
            .sr(N__51684));
    defparam sDAC_data_RNO_25_10_LC_15_13_7.C_ON=1'b0;
    defparam sDAC_data_RNO_25_10_LC_15_13_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_10_LC_15_13_7.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_25_10_LC_15_13_7 (
            .in0(N__38448),
            .in1(N__33470),
            .in2(N__38203),
            .in3(N__33464),
            .lcout(sDAC_data_2_39_ns_1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_10_LC_15_14_0.C_ON=1'b0;
    defparam sDAC_data_RNO_24_10_LC_15_14_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_10_LC_15_14_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_10_LC_15_14_0 (
            .in0(N__41606),
            .in1(N__33458),
            .in2(_gnd_net_),
            .in3(N__33449),
            .lcout(sDAC_data_RNO_24Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_10_LC_15_14_1.C_ON=1'b0;
    defparam sDAC_data_RNO_23_10_LC_15_14_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_10_LC_15_14_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_10_LC_15_14_1 (
            .in0(N__41609),
            .in1(N__33434),
            .in2(_gnd_net_),
            .in3(N__33395),
            .lcout(),
            .ltout(sDAC_data_RNO_23Z0Z_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_10_LC_15_14_2.C_ON=1'b0;
    defparam sDAC_data_RNO_11_10_LC_15_14_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_10_LC_15_14_2.LUT_INIT=16'b1010000011011101;
    LogicCell40 sDAC_data_RNO_11_10_LC_15_14_2 (
            .in0(N__38117),
            .in1(N__33419),
            .in2(N__33413),
            .in3(N__33410),
            .lcout(sDAC_data_RNO_11Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_28_7_LC_15_14_3.C_ON=1'b0;
    defparam sDAC_mem_28_7_LC_15_14_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_7_LC_15_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_7_LC_15_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50057),
            .lcout(sDAC_mem_28Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52246),
            .ce(N__37808),
            .sr(N__51679));
    defparam sDAC_data_RNO_31_3_LC_15_14_4.C_ON=1'b0;
    defparam sDAC_data_RNO_31_3_LC_15_14_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_3_LC_15_14_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_31_3_LC_15_14_4 (
            .in0(N__41605),
            .in1(N__33650),
            .in2(_gnd_net_),
            .in3(N__33644),
            .lcout(sDAC_data_RNO_31Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_30_3_LC_15_14_5.C_ON=1'b0;
    defparam sDAC_data_RNO_30_3_LC_15_14_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_3_LC_15_14_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_30_3_LC_15_14_5 (
            .in0(N__41608),
            .in1(N__41324),
            .in2(_gnd_net_),
            .in3(N__33635),
            .lcout(),
            .ltout(sDAC_data_RNO_30Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_25_3_LC_15_14_6.C_ON=1'b0;
    defparam sDAC_data_RNO_25_3_LC_15_14_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_3_LC_15_14_6.LUT_INIT=16'b0100010101100111;
    LogicCell40 sDAC_data_RNO_25_3_LC_15_14_6 (
            .in0(N__38402),
            .in1(N__38121),
            .in2(N__33620),
            .in3(N__33617),
            .lcout(),
            .ltout(sDAC_data_2_39_ns_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_3_LC_15_14_7.C_ON=1'b0;
    defparam sDAC_data_RNO_11_3_LC_15_14_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_3_LC_15_14_7.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_11_3_LC_15_14_7 (
            .in0(N__38122),
            .in1(N__33611),
            .in2(N__33605),
            .in3(N__33845),
            .lcout(sDAC_data_RNO_11Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_21_7_LC_15_15_0.C_ON=1'b0;
    defparam sDAC_data_RNO_21_7_LC_15_15_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_7_LC_15_15_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_7_LC_15_15_0 (
            .in0(N__41866),
            .in1(N__36764),
            .in2(_gnd_net_),
            .in3(N__33587),
            .lcout(sDAC_data_RNO_21Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_22_4_LC_15_15_1.C_ON=1'b0;
    defparam sDAC_mem_22_4_LC_15_15_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_4_LC_15_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_4_LC_15_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45603),
            .lcout(sDAC_mem_22Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52256),
            .ce(N__33893),
            .sr(N__51671));
    defparam sDAC_data_RNO_21_8_LC_15_15_2.C_ON=1'b0;
    defparam sDAC_data_RNO_21_8_LC_15_15_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_8_LC_15_15_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_8_LC_15_15_2 (
            .in0(N__41868),
            .in1(N__36746),
            .in2(_gnd_net_),
            .in3(N__33566),
            .lcout(sDAC_data_RNO_21Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_22_5_LC_15_15_3.C_ON=1'b0;
    defparam sDAC_mem_22_5_LC_15_15_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_5_LC_15_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_5_LC_15_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45118),
            .lcout(sDAC_mem_22Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52256),
            .ce(N__33893),
            .sr(N__51671));
    defparam sDAC_data_RNO_21_9_LC_15_15_4.C_ON=1'b0;
    defparam sDAC_data_RNO_21_9_LC_15_15_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_9_LC_15_15_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_9_LC_15_15_4 (
            .in0(N__41867),
            .in1(N__36728),
            .in2(_gnd_net_),
            .in3(N__33899),
            .lcout(sDAC_data_RNO_21Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_22_6_LC_15_15_5.C_ON=1'b0;
    defparam sDAC_mem_22_6_LC_15_15_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_6_LC_15_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_6_LC_15_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50542),
            .lcout(sDAC_mem_22Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52256),
            .ce(N__33893),
            .sr(N__51671));
    defparam sDAC_data_RNO_23_3_LC_15_15_6.C_ON=1'b0;
    defparam sDAC_data_RNO_23_3_LC_15_15_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_3_LC_15_15_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_3_LC_15_15_6 (
            .in0(N__41865),
            .in1(N__33869),
            .in2(_gnd_net_),
            .in3(N__33860),
            .lcout(sDAC_data_RNO_23Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_6_LC_15_15_7.C_ON=1'b0;
    defparam sDAC_data_RNO_23_6_LC_15_15_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_6_LC_15_15_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_6_LC_15_15_7 (
            .in0(N__41985),
            .in1(N__33839),
            .in2(_gnd_net_),
            .in3(N__33827),
            .lcout(sDAC_data_RNO_23Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_4_LC_15_16_0.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_4_LC_15_16_0.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_4_LC_15_16_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_4_LC_15_16_0 (
            .in0(N__35344),
            .in1(N__35122),
            .in2(N__35330),
            .in3(N__35359),
            .lcout(sbuttonModeStatus_0_sqmuxa_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_5_LC_15_16_1.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_5_LC_15_16_1.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_5_LC_15_16_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_5_LC_15_16_1 (
            .in0(N__35180),
            .in1(N__35141),
            .in2(N__35285),
            .in3(N__35162),
            .lcout(),
            .ltout(sbuttonModeStatus_0_sqmuxa_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_2_LC_15_16_2.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_2_LC_15_16_2.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_2_LC_15_16_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_2_LC_15_16_2 (
            .in0(N__38843),
            .in1(N__38765),
            .in2(N__33812),
            .in3(N__33809),
            .lcout(sbuttonModeStatus_0_sqmuxa_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_6_LC_15_16_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_6_LC_15_16_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_6_LC_15_16_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 sAddress_RNI9IH12_6_LC_15_16_3 (
            .in0(N__33791),
            .in1(N__40072),
            .in2(_gnd_net_),
            .in3(N__33773),
            .lcout(sEEPonPoff_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_nWE_obuf_RNO_LC_15_16_6.C_ON=1'b0;
    defparam RAM_nWE_obuf_RNO_LC_15_16_6.SEQ_MODE=4'b0000;
    defparam RAM_nWE_obuf_RNO_LC_15_16_6.LUT_INIT=16'b1111111101010101;
    LogicCell40 RAM_nWE_obuf_RNO_LC_15_16_6 (
            .in0(N__48961),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34015),
            .lcout(RAM_nWE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sRead_data_RNO_0_LC_15_17_1.C_ON=1'b0;
    defparam sRead_data_RNO_0_LC_15_17_1.SEQ_MODE=4'b0000;
    defparam sRead_data_RNO_0_LC_15_17_1.LUT_INIT=16'b1100110011111111;
    LogicCell40 sRead_data_RNO_0_LC_15_17_1 (
            .in0(_gnd_net_),
            .in1(N__39163),
            .in2(_gnd_net_),
            .in3(N__39139),
            .lcout(),
            .ltout(sRead_data_RNOZ0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sRead_data_LC_15_17_2.C_ON=1'b0;
    defparam sRead_data_LC_15_17_2.SEQ_MODE=4'b1010;
    defparam sRead_data_LC_15_17_2.LUT_INIT=16'b1010101010001100;
    LogicCell40 sRead_data_LC_15_17_2 (
            .in0(N__33983),
            .in1(N__43735),
            .in2(N__34031),
            .in3(N__48952),
            .lcout(sRead_dataZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52277),
            .ce(),
            .sr(N__51658));
    defparam sCounterRAM_RNIS8L63_1_LC_15_17_4.C_ON=1'b0;
    defparam sCounterRAM_RNIS8L63_1_LC_15_17_4.SEQ_MODE=4'b0000;
    defparam sCounterRAM_RNIS8L63_1_LC_15_17_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounterRAM_RNIS8L63_1_LC_15_17_4 (
            .in0(N__39029),
            .in1(N__33965),
            .in2(N__39608),
            .in3(N__33971),
            .lcout(N_75),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sSPI_MSB0LSB1_LC_15_17_5.C_ON=1'b0;
    defparam sSPI_MSB0LSB1_LC_15_17_5.SEQ_MODE=4'b1010;
    defparam sSPI_MSB0LSB1_LC_15_17_5.LUT_INIT=16'b1001001111001100;
    LogicCell40 sSPI_MSB0LSB1_LC_15_17_5 (
            .in0(N__43336),
            .in1(N__39164),
            .in2(N__43487),
            .in3(N__39140),
            .lcout(sSPI_MSB0LSBZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52277),
            .ce(),
            .sr(N__51658));
    defparam sADC_clk_LC_15_17_6.C_ON=1'b0;
    defparam sADC_clk_LC_15_17_6.SEQ_MODE=4'b1010;
    defparam sADC_clk_LC_15_17_6.LUT_INIT=16'b0100100000000000;
    LogicCell40 sADC_clk_LC_15_17_6 (
            .in0(N__34006),
            .in1(N__43335),
            .in2(N__46970),
            .in3(N__43446),
            .lcout(ADC_clk_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52277),
            .ce(),
            .sr(N__51658));
    defparam sRead_data_RNI74VQ_LC_15_18_6.C_ON=1'b0;
    defparam sRead_data_RNI74VQ_LC_15_18_6.SEQ_MODE=4'b0000;
    defparam sRead_data_RNI74VQ_LC_15_18_6.LUT_INIT=16'b1111111111011101;
    LogicCell40 sRead_data_RNI74VQ_LC_15_18_6 (
            .in0(N__33982),
            .in1(N__39548),
            .in2(_gnd_net_),
            .in3(N__39566),
            .lcout(spi_data_miso_0_sqmuxa_2_i_o2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterRAM_RNISREI1_7_LC_15_18_7.C_ON=1'b0;
    defparam sCounterRAM_RNISREI1_7_LC_15_18_7.SEQ_MODE=4'b0000;
    defparam sCounterRAM_RNISREI1_7_LC_15_18_7.LUT_INIT=16'b1111111011111111;
    LogicCell40 sCounterRAM_RNISREI1_7_LC_15_18_7 (
            .in0(N__39530),
            .in1(N__39047),
            .in2(N__39479),
            .in3(N__39584),
            .lcout(spi_data_miso_0_sqmuxa_2_i_o2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_1_3_LC_15_20_4.C_ON=1'b0;
    defparam RAM_DATA_1_3_LC_15_20_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_3_LC_15_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_3_LC_15_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33959),
            .lcout(RAM_DATA_1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52311),
            .ce(N__51890),
            .sr(N__51647));
    defparam sDAC_mem_19_4_LC_16_3_0.C_ON=1'b0;
    defparam sDAC_mem_19_4_LC_16_3_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_4_LC_16_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_4_LC_16_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45508),
            .lcout(sDAC_mem_19Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52290),
            .ce(N__34997),
            .sr(N__51806));
    defparam sDAC_mem_19_5_LC_16_3_1.C_ON=1'b0;
    defparam sDAC_mem_19_5_LC_16_3_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_5_LC_16_3_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_5_LC_16_3_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44982),
            .lcout(sDAC_mem_19Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52290),
            .ce(N__34997),
            .sr(N__51806));
    defparam sDAC_mem_19_6_LC_16_3_2.C_ON=1'b0;
    defparam sDAC_mem_19_6_LC_16_3_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_6_LC_16_3_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_6_LC_16_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50484),
            .lcout(sDAC_mem_19Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52290),
            .ce(N__34997),
            .sr(N__51806));
    defparam sDAC_mem_19_7_LC_16_3_3.C_ON=1'b0;
    defparam sDAC_mem_19_7_LC_16_3_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_7_LC_16_3_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_7_LC_16_3_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50054),
            .lcout(sDAC_mem_19Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52290),
            .ce(N__34997),
            .sr(N__51806));
    defparam sDAC_mem_21_0_LC_16_4_0.C_ON=1'b0;
    defparam sDAC_mem_21_0_LC_16_4_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_0_LC_16_4_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_21_0_LC_16_4_0 (
            .in0(N__46385),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_21Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52278),
            .ce(N__34247),
            .sr(N__51797));
    defparam sDAC_mem_21_1_LC_16_4_1.C_ON=1'b0;
    defparam sDAC_mem_21_1_LC_16_4_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_1_LC_16_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_1_LC_16_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51053),
            .lcout(sDAC_mem_21Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52278),
            .ce(N__34247),
            .sr(N__51797));
    defparam sDAC_mem_21_2_LC_16_4_2.C_ON=1'b0;
    defparam sDAC_mem_21_2_LC_16_4_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_2_LC_16_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_2_LC_16_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47348),
            .lcout(sDAC_mem_21Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52278),
            .ce(N__34247),
            .sr(N__51797));
    defparam sDAC_mem_21_3_LC_16_4_3.C_ON=1'b0;
    defparam sDAC_mem_21_3_LC_16_4_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_3_LC_16_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_3_LC_16_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46751),
            .lcout(sDAC_mem_21Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52278),
            .ce(N__34247),
            .sr(N__51797));
    defparam sDAC_mem_21_4_LC_16_4_4.C_ON=1'b0;
    defparam sDAC_mem_21_4_LC_16_4_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_4_LC_16_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_4_LC_16_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45507),
            .lcout(sDAC_mem_21Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52278),
            .ce(N__34247),
            .sr(N__51797));
    defparam sDAC_mem_21_5_LC_16_4_5.C_ON=1'b0;
    defparam sDAC_mem_21_5_LC_16_4_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_5_LC_16_4_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_21_5_LC_16_4_5 (
            .in0(N__44981),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_21Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52278),
            .ce(N__34247),
            .sr(N__51797));
    defparam sDAC_mem_21_6_LC_16_4_6.C_ON=1'b0;
    defparam sDAC_mem_21_6_LC_16_4_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_6_LC_16_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_6_LC_16_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50483),
            .lcout(sDAC_mem_21Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52278),
            .ce(N__34247),
            .sr(N__51797));
    defparam sDAC_mem_21_7_LC_16_4_7.C_ON=1'b0;
    defparam sDAC_mem_21_7_LC_16_4_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_7_LC_16_4_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_7_LC_16_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50053),
            .lcout(sDAC_mem_21Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52278),
            .ce(N__34247),
            .sr(N__51797));
    defparam sDAC_mem_3_4_LC_16_5_0.C_ON=1'b0;
    defparam sDAC_mem_3_4_LC_16_5_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_4_LC_16_5_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_3_4_LC_16_5_0 (
            .in0(N__45349),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_3Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52268),
            .ce(N__44237),
            .sr(N__51783));
    defparam sDAC_data_RNO_27_7_LC_16_5_1.C_ON=1'b0;
    defparam sDAC_data_RNO_27_7_LC_16_5_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_7_LC_16_5_1.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_27_7_LC_16_5_1 (
            .in0(N__42557),
            .in1(N__34235),
            .in2(N__42264),
            .in3(N__34223),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_7_LC_16_5_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_7_LC_16_5_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_7_LC_16_5_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_7_LC_16_5_2 (
            .in0(N__42095),
            .in1(N__34211),
            .in2(N__34196),
            .in3(N__34193),
            .lcout(sDAC_data_RNO_15Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_7_LC_16_5_3.C_ON=1'b0;
    defparam sDAC_data_RNO_16_7_LC_16_5_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_7_LC_16_5_3.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_16_7_LC_16_5_3 (
            .in0(N__42558),
            .in1(N__34181),
            .in2(N__42265),
            .in3(N__34169),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_7_LC_16_5_4.C_ON=1'b0;
    defparam sDAC_data_RNO_7_7_LC_16_5_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_7_LC_16_5_4.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_7_7_LC_16_5_4 (
            .in0(N__36800),
            .in1(N__42259),
            .in2(N__34157),
            .in3(N__39680),
            .lcout(),
            .ltout(sDAC_data_RNO_7Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_7_LC_16_5_5.C_ON=1'b0;
    defparam sDAC_data_RNO_2_7_LC_16_5_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_7_LC_16_5_5.LUT_INIT=16'b0111010101100100;
    LogicCell40 sDAC_data_RNO_2_7_LC_16_5_5 (
            .in0(N__34154),
            .in1(N__38131),
            .in2(N__34145),
            .in3(N__34121),
            .lcout(sDAC_data_RNO_2Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_7_LC_16_5_6.C_ON=1'b0;
    defparam sDAC_data_RNO_8_7_LC_16_5_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_7_LC_16_5_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_8_7_LC_16_5_6 (
            .in0(N__42096),
            .in1(N__34136),
            .in2(_gnd_net_),
            .in3(N__34097),
            .lcout(sDAC_data_RNO_8Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_7_LC_16_5_7.C_ON=1'b0;
    defparam sDAC_data_RNO_17_7_LC_16_5_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_7_LC_16_5_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_7_LC_16_5_7 (
            .in0(N__42556),
            .in1(N__34115),
            .in2(_gnd_net_),
            .in3(N__34106),
            .lcout(sDAC_data_RNO_17Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_3_6_LC_16_6_0.C_ON=1'b0;
    defparam sDAC_mem_3_6_LC_16_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_6_LC_16_6_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_3_6_LC_16_6_0 (
            .in0(N__50430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_3Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52257),
            .ce(N__44244),
            .sr(N__51771));
    defparam sDAC_data_RNO_27_9_LC_16_6_1.C_ON=1'b0;
    defparam sDAC_data_RNO_27_9_LC_16_6_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_9_LC_16_6_1.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_27_9_LC_16_6_1 (
            .in0(N__42551),
            .in1(N__34376),
            .in2(N__42239),
            .in3(N__34364),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_9_LC_16_6_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_9_LC_16_6_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_9_LC_16_6_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_9_LC_16_6_2 (
            .in0(N__42165),
            .in1(N__34355),
            .in2(N__34346),
            .in3(N__34343),
            .lcout(sDAC_data_RNO_15Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_9_LC_16_6_3.C_ON=1'b0;
    defparam sDAC_data_RNO_17_9_LC_16_6_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_9_LC_16_6_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_9_LC_16_6_3 (
            .in0(N__42552),
            .in1(N__34331),
            .in2(_gnd_net_),
            .in3(N__34316),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_9_LC_16_6_4.C_ON=1'b0;
    defparam sDAC_data_RNO_8_9_LC_16_6_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_9_LC_16_6_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_8_9_LC_16_6_4 (
            .in0(_gnd_net_),
            .in1(N__42157),
            .in2(N__34301),
            .in3(N__34298),
            .lcout(sDAC_data_RNO_8Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_9_LC_16_6_5.C_ON=1'b0;
    defparam sDAC_data_RNO_16_9_LC_16_6_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_9_LC_16_6_5.LUT_INIT=16'b0001110000011111;
    LogicCell40 sDAC_data_RNO_16_9_LC_16_6_5 (
            .in0(N__34289),
            .in1(N__42166),
            .in2(N__42575),
            .in3(N__34277),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_9_LC_16_6_6.C_ON=1'b0;
    defparam sDAC_data_RNO_7_9_LC_16_6_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_9_LC_16_6_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_7_9_LC_16_6_6 (
            .in0(N__42167),
            .in1(N__39842),
            .in2(N__34265),
            .in3(N__37040),
            .lcout(),
            .ltout(sDAC_data_RNO_7Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_9_LC_16_6_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_9_LC_16_6_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_9_LC_16_6_7.LUT_INIT=16'b0111001101100010;
    LogicCell40 sDAC_data_RNO_2_9_LC_16_6_7 (
            .in0(N__38031),
            .in1(N__36983),
            .in2(N__34262),
            .in3(N__34259),
            .lcout(sDAC_data_RNO_2Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_32_6_LC_16_7_0.C_ON=1'b0;
    defparam sDAC_mem_32_6_LC_16_7_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_6_LC_16_7_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_32_6_LC_16_7_0 (
            .in0(N__50486),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_32Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52247),
            .ce(N__41265),
            .sr(N__51758));
    defparam sDAC_data_RNO_26_9_LC_16_7_1.C_ON=1'b0;
    defparam sDAC_data_RNO_26_9_LC_16_7_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_9_LC_16_7_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_26_9_LC_16_7_1 (
            .in0(N__42430),
            .in1(N__44324),
            .in2(_gnd_net_),
            .in3(N__44423),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_9_LC_16_7_2.C_ON=1'b0;
    defparam sDAC_data_RNO_14_9_LC_16_7_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_9_LC_16_7_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 sDAC_data_RNO_14_9_LC_16_7_2 (
            .in0(N__42111),
            .in1(_gnd_net_),
            .in2(N__34469),
            .in3(N__34466),
            .lcout(sDAC_data_RNO_14Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_20_3_LC_16_7_3.C_ON=1'b0;
    defparam sDAC_data_RNO_20_3_LC_16_7_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_3_LC_16_7_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_20_3_LC_16_7_3 (
            .in0(N__34454),
            .in1(N__42105),
            .in2(_gnd_net_),
            .in3(N__36449),
            .lcout(sDAC_data_RNO_20Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_20_4_LC_16_7_4.C_ON=1'b0;
    defparam sDAC_data_RNO_20_4_LC_16_7_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_4_LC_16_7_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_20_4_LC_16_7_4 (
            .in0(N__42104),
            .in1(N__34445),
            .in2(_gnd_net_),
            .in3(N__36437),
            .lcout(sDAC_data_RNO_20Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_20_5_LC_16_7_5.C_ON=1'b0;
    defparam sDAC_data_RNO_20_5_LC_16_7_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_5_LC_16_7_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_20_5_LC_16_7_5 (
            .in0(N__34424),
            .in1(N__42109),
            .in2(_gnd_net_),
            .in3(N__36425),
            .lcout(sDAC_data_RNO_20Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_20_6_LC_16_7_6.C_ON=1'b0;
    defparam sDAC_data_RNO_20_6_LC_16_7_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_6_LC_16_7_6.LUT_INIT=16'b1111101000001010;
    LogicCell40 sDAC_data_RNO_20_6_LC_16_7_6 (
            .in0(N__36413),
            .in1(_gnd_net_),
            .in2(N__42214),
            .in3(N__34415),
            .lcout(sDAC_data_RNO_20Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_20_7_LC_16_7_7.C_ON=1'b0;
    defparam sDAC_data_RNO_20_7_LC_16_7_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_7_LC_16_7_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_20_7_LC_16_7_7 (
            .in0(N__34394),
            .in1(N__42110),
            .in2(_gnd_net_),
            .in3(N__36662),
            .lcout(sDAC_data_RNO_20Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_pointer_RNI3NFH_1_LC_16_8_0.C_ON=1'b1;
    defparam sDAC_mem_pointer_RNI3NFH_1_LC_16_8_0.SEQ_MODE=4'b0000;
    defparam sDAC_mem_pointer_RNI3NFH_1_LC_16_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 sDAC_mem_pointer_RNI3NFH_1_LC_16_8_0 (
            .in0(_gnd_net_),
            .in1(N__42168),
            .in2(N__38552),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(sDAC_mem_pointer_0_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_pointer_2_LC_16_8_1.C_ON=1'b1;
    defparam sDAC_mem_pointer_2_LC_16_8_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_2_LC_16_8_1.LUT_INIT=16'b0010001010001000;
    LogicCell40 sDAC_mem_pointer_2_LC_16_8_1 (
            .in0(N__37632),
            .in1(N__38001),
            .in2(_gnd_net_),
            .in3(N__34577),
            .lcout(sDAC_mem_pointerZ0Z_2),
            .ltout(),
            .carryin(sDAC_mem_pointer_0_cry_1),
            .carryout(sDAC_mem_pointer_0_cry_2),
            .clk(N__48462),
            .ce(N__43949),
            .sr(N__51746));
    defparam sDAC_mem_pointer_3_LC_16_8_2.C_ON=1'b1;
    defparam sDAC_mem_pointer_3_LC_16_8_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_3_LC_16_8_2.LUT_INIT=16'b0010001010001000;
    LogicCell40 sDAC_mem_pointer_3_LC_16_8_2 (
            .in0(N__37635),
            .in1(N__37327),
            .in2(_gnd_net_),
            .in3(N__34574),
            .lcout(sDAC_mem_pointerZ0Z_3),
            .ltout(),
            .carryin(sDAC_mem_pointer_0_cry_2),
            .carryout(sDAC_mem_pointer_0_cry_3),
            .clk(N__48462),
            .ce(N__43949),
            .sr(N__51746));
    defparam sDAC_mem_pointer_4_LC_16_8_3.C_ON=1'b1;
    defparam sDAC_mem_pointer_4_LC_16_8_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_4_LC_16_8_3.LUT_INIT=16'b0010001010001000;
    LogicCell40 sDAC_mem_pointer_4_LC_16_8_3 (
            .in0(N__37633),
            .in1(N__37419),
            .in2(_gnd_net_),
            .in3(N__34571),
            .lcout(sDAC_mem_pointerZ0Z_4),
            .ltout(),
            .carryin(sDAC_mem_pointer_0_cry_3),
            .carryout(sDAC_mem_pointer_0_cry_4),
            .clk(N__48462),
            .ce(N__43949),
            .sr(N__51746));
    defparam sDAC_mem_pointer_5_LC_16_8_4.C_ON=1'b0;
    defparam sDAC_mem_pointer_5_LC_16_8_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_5_LC_16_8_4.LUT_INIT=16'b0100010010001000;
    LogicCell40 sDAC_mem_pointer_5_LC_16_8_4 (
            .in0(N__42433),
            .in1(N__37634),
            .in2(_gnd_net_),
            .in3(N__34568),
            .lcout(sDAC_mem_pointerZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48462),
            .ce(N__43949),
            .sr(N__51746));
    defparam sDAC_mem_3_2_LC_16_9_0.C_ON=1'b0;
    defparam sDAC_mem_3_2_LC_16_9_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_2_LC_16_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_3_2_LC_16_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47447),
            .lcout(sDAC_mem_3Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52225),
            .ce(N__44246),
            .sr(N__51731));
    defparam sDAC_data_RNO_27_5_LC_16_9_1.C_ON=1'b0;
    defparam sDAC_data_RNO_27_5_LC_16_9_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_5_LC_16_9_1.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_27_5_LC_16_9_1 (
            .in0(N__42427),
            .in1(N__34565),
            .in2(N__42240),
            .in3(N__34553),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_5_LC_16_9_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_5_LC_16_9_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_5_LC_16_9_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_5_LC_16_9_2 (
            .in0(N__42143),
            .in1(N__34541),
            .in2(N__34523),
            .in3(N__34520),
            .lcout(sDAC_data_RNO_15Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_5_LC_16_9_3.C_ON=1'b0;
    defparam sDAC_data_RNO_17_5_LC_16_9_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_5_LC_16_9_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_5_LC_16_9_3 (
            .in0(N__42428),
            .in1(N__34514),
            .in2(_gnd_net_),
            .in3(N__34502),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_5_LC_16_9_4.C_ON=1'b0;
    defparam sDAC_data_RNO_8_5_LC_16_9_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_5_LC_16_9_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_8_5_LC_16_9_4 (
            .in0(_gnd_net_),
            .in1(N__42161),
            .in2(N__34487),
            .in3(N__34484),
            .lcout(sDAC_data_RNO_8Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_5_LC_16_9_5.C_ON=1'b0;
    defparam sDAC_data_RNO_16_5_LC_16_9_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_5_LC_16_9_5.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_16_5_LC_16_9_5 (
            .in0(N__42429),
            .in1(N__34757),
            .in2(N__42241),
            .in3(N__34742),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_5_LC_16_9_6.C_ON=1'b0;
    defparam sDAC_data_RNO_7_5_LC_16_9_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_5_LC_16_9_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_7_5_LC_16_9_6 (
            .in0(N__42144),
            .in1(N__39884),
            .in2(N__34727),
            .in3(N__36821),
            .lcout(),
            .ltout(sDAC_data_RNO_7Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_5_LC_16_9_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_5_LC_16_9_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_5_LC_16_9_7.LUT_INIT=16'b0111001101100010;
    LogicCell40 sDAC_data_RNO_2_5_LC_16_9_7 (
            .in0(N__37997),
            .in1(N__34724),
            .in2(N__34715),
            .in3(N__34712),
            .lcout(sDAC_data_RNO_2Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_3_0_LC_16_10_0.C_ON=1'b0;
    defparam sDAC_mem_3_0_LC_16_10_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_0_LC_16_10_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_3_0_LC_16_10_0 (
            .in0(N__46314),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52219),
            .ce(N__44245),
            .sr(N__51719));
    defparam sDAC_data_RNO_27_3_LC_16_10_1.C_ON=1'b0;
    defparam sDAC_data_RNO_27_3_LC_16_10_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_3_LC_16_10_1.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_27_3_LC_16_10_1 (
            .in0(N__42522),
            .in1(N__34706),
            .in2(N__42174),
            .in3(N__34694),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_3_LC_16_10_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_3_LC_16_10_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_3_LC_16_10_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_3_LC_16_10_2 (
            .in0(N__41983),
            .in1(N__34682),
            .in2(N__34664),
            .in3(N__34661),
            .lcout(sDAC_data_RNO_15Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_3_LC_16_10_3.C_ON=1'b0;
    defparam sDAC_data_RNO_17_3_LC_16_10_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_3_LC_16_10_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_3_LC_16_10_3 (
            .in0(N__42523),
            .in1(N__34655),
            .in2(_gnd_net_),
            .in3(N__34637),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_3_LC_16_10_4.C_ON=1'b0;
    defparam sDAC_data_RNO_8_3_LC_16_10_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_3_LC_16_10_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_8_3_LC_16_10_4 (
            .in0(_gnd_net_),
            .in1(N__42006),
            .in2(N__34622),
            .in3(N__34619),
            .lcout(sDAC_data_RNO_8Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_3_LC_16_10_5.C_ON=1'b0;
    defparam sDAC_data_RNO_16_3_LC_16_10_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_3_LC_16_10_5.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_16_3_LC_16_10_5 (
            .in0(N__42524),
            .in1(N__34607),
            .in2(N__42175),
            .in3(N__34592),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_3_LC_16_10_6.C_ON=1'b0;
    defparam sDAC_data_RNO_7_3_LC_16_10_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_3_LC_16_10_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_7_3_LC_16_10_6 (
            .in0(N__41984),
            .in1(N__39908),
            .in2(N__34898),
            .in3(N__36845),
            .lcout(),
            .ltout(sDAC_data_RNO_7Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_3_LC_16_10_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_3_LC_16_10_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_3_LC_16_10_7.LUT_INIT=16'b0111001101100010;
    LogicCell40 sDAC_data_RNO_2_3_LC_16_10_7 (
            .in0(N__38097),
            .in1(N__34895),
            .in2(N__34883),
            .in3(N__34880),
            .lcout(sDAC_data_RNO_2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_8_3_LC_16_11_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_8_3_LC_16_11_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_8_3_LC_16_11_0.LUT_INIT=16'b0001000100000000;
    LogicCell40 sAddress_RNI9IH12_8_3_LC_16_11_0 (
            .in0(N__40428),
            .in1(N__34874),
            .in2(_gnd_net_),
            .in3(N__40028),
            .lcout(sDAC_mem_19_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_19_0_LC_16_11_1.C_ON=1'b0;
    defparam sDAC_mem_19_0_LC_16_11_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_0_LC_16_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_0_LC_16_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46315),
            .lcout(sDAC_mem_19Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52212),
            .ce(N__34990),
            .sr(N__51708));
    defparam sDAC_data_RNO_29_3_LC_16_11_2.C_ON=1'b0;
    defparam sDAC_data_RNO_29_3_LC_16_11_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_3_LC_16_11_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_29_3_LC_16_11_2 (
            .in0(N__41885),
            .in1(N__34829),
            .in2(_gnd_net_),
            .in3(N__34823),
            .lcout(sDAC_data_RNO_29Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_19_1_LC_16_11_3.C_ON=1'b0;
    defparam sDAC_mem_19_1_LC_16_11_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_1_LC_16_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_1_LC_16_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50985),
            .lcout(sDAC_mem_19Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52212),
            .ce(N__34990),
            .sr(N__51708));
    defparam sDAC_data_RNO_29_4_LC_16_11_4.C_ON=1'b0;
    defparam sDAC_data_RNO_29_4_LC_16_11_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_4_LC_16_11_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_29_4_LC_16_11_4 (
            .in0(N__41884),
            .in1(N__34808),
            .in2(_gnd_net_),
            .in3(N__34802),
            .lcout(sDAC_data_RNO_29Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_19_2_LC_16_11_5.C_ON=1'b0;
    defparam sDAC_mem_19_2_LC_16_11_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_2_LC_16_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_2_LC_16_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47496),
            .lcout(sDAC_mem_19Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52212),
            .ce(N__34990),
            .sr(N__51708));
    defparam sDAC_data_RNO_29_5_LC_16_11_6.C_ON=1'b0;
    defparam sDAC_data_RNO_29_5_LC_16_11_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_5_LC_16_11_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_29_5_LC_16_11_6 (
            .in0(N__41886),
            .in1(N__34775),
            .in2(_gnd_net_),
            .in3(N__34769),
            .lcout(sDAC_data_RNO_29Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_19_3_LC_16_11_7.C_ON=1'b0;
    defparam sDAC_mem_19_3_LC_16_11_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_3_LC_16_11_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_19_3_LC_16_11_7 (
            .in0(N__46854),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_19Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52212),
            .ce(N__34990),
            .sr(N__51708));
    defparam sDAC_data_RNO_15_10_LC_16_12_0.C_ON=1'b0;
    defparam sDAC_data_RNO_15_10_LC_16_12_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_10_LC_16_12_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_15_10_LC_16_12_0 (
            .in0(N__34976),
            .in1(N__44261),
            .in2(N__42170),
            .in3(N__34964),
            .lcout(),
            .ltout(sDAC_data_RNO_15Z0Z_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_10_LC_16_12_1.C_ON=1'b0;
    defparam sDAC_data_RNO_6_10_LC_16_12_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_10_LC_16_12_1.LUT_INIT=16'b0010011000110111;
    LogicCell40 sDAC_data_RNO_6_10_LC_16_12_1 (
            .in0(N__38231),
            .in1(N__38526),
            .in2(N__34958),
            .in3(N__34904),
            .lcout(),
            .ltout(sDAC_data_2_14_ns_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_10_LC_16_12_2.C_ON=1'b0;
    defparam sDAC_data_RNO_1_10_LC_16_12_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_10_LC_16_12_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_1_10_LC_16_12_2 (
            .in0(N__38030),
            .in1(N__34955),
            .in2(N__34946),
            .in3(N__34916),
            .lcout(sDAC_data_RNO_1Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_26_10_LC_16_12_3.C_ON=1'b0;
    defparam sDAC_data_RNO_26_10_LC_16_12_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_10_LC_16_12_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_26_10_LC_16_12_3 (
            .in0(N__44414),
            .in1(N__42513),
            .in2(_gnd_net_),
            .in3(N__44543),
            .lcout(sDAC_data_RNO_26Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_12_10_LC_16_12_4.C_ON=1'b0;
    defparam sDAC_data_RNO_12_10_LC_16_12_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_10_LC_16_12_4.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_12_10_LC_16_12_4 (
            .in0(N__42514),
            .in1(N__34937),
            .in2(N__42169),
            .in3(N__36461),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_10_LC_16_12_5.C_ON=1'b0;
    defparam sDAC_data_RNO_4_10_LC_16_12_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_10_LC_16_12_5.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_10_LC_16_12_5 (
            .in0(N__41982),
            .in1(N__41087),
            .in2(N__34919),
            .in3(N__44447),
            .lcout(sDAC_data_RNO_4Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_10_LC_16_12_6.C_ON=1'b0;
    defparam sDAC_data_RNO_14_10_LC_16_12_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_10_LC_16_12_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_14_10_LC_16_12_6 (
            .in0(N__41975),
            .in1(N__39623),
            .in2(_gnd_net_),
            .in3(N__34910),
            .lcout(sDAC_data_RNO_14Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_button_debounce_counter_cry_1_c_LC_16_13_0.C_ON=1'b1;
    defparam un1_button_debounce_counter_cry_1_c_LC_16_13_0.SEQ_MODE=4'b0000;
    defparam un1_button_debounce_counter_cry_1_c_LC_16_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_button_debounce_counter_cry_1_c_LC_16_13_0 (
            .in0(_gnd_net_),
            .in1(N__45772),
            .in2(N__45751),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(un1_button_debounce_counter_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam button_debounce_counter_2_LC_16_13_1.C_ON=1'b1;
    defparam button_debounce_counter_2_LC_16_13_1.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_2_LC_16_13_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_2_LC_16_13_1 (
            .in0(N__49428),
            .in1(N__35101),
            .in2(_gnd_net_),
            .in3(N__35090),
            .lcout(button_debounce_counterZ0Z_2),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_1),
            .carryout(un1_button_debounce_counter_cry_2),
            .clk(N__48476),
            .ce(),
            .sr(N__45714));
    defparam button_debounce_counter_3_LC_16_13_2.C_ON=1'b1;
    defparam button_debounce_counter_3_LC_16_13_2.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_3_LC_16_13_2.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_3_LC_16_13_2 (
            .in0(N__49191),
            .in1(N__35086),
            .in2(_gnd_net_),
            .in3(N__35075),
            .lcout(button_debounce_counterZ0Z_3),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_2),
            .carryout(un1_button_debounce_counter_cry_3),
            .clk(N__48476),
            .ce(),
            .sr(N__45714));
    defparam button_debounce_counter_4_LC_16_13_3.C_ON=1'b1;
    defparam button_debounce_counter_4_LC_16_13_3.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_4_LC_16_13_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_4_LC_16_13_3 (
            .in0(N__49429),
            .in1(N__35071),
            .in2(_gnd_net_),
            .in3(N__35060),
            .lcout(button_debounce_counterZ0Z_4),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_3),
            .carryout(un1_button_debounce_counter_cry_4),
            .clk(N__48476),
            .ce(),
            .sr(N__45714));
    defparam button_debounce_counter_5_LC_16_13_4.C_ON=1'b1;
    defparam button_debounce_counter_5_LC_16_13_4.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_5_LC_16_13_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_5_LC_16_13_4 (
            .in0(N__49192),
            .in1(N__35053),
            .in2(_gnd_net_),
            .in3(N__35042),
            .lcout(button_debounce_counterZ0Z_5),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_4),
            .carryout(un1_button_debounce_counter_cry_5),
            .clk(N__48476),
            .ce(),
            .sr(N__45714));
    defparam button_debounce_counter_6_LC_16_13_5.C_ON=1'b1;
    defparam button_debounce_counter_6_LC_16_13_5.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_6_LC_16_13_5.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_6_LC_16_13_5 (
            .in0(N__49430),
            .in1(N__35035),
            .in2(_gnd_net_),
            .in3(N__35024),
            .lcout(button_debounce_counterZ0Z_6),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_5),
            .carryout(un1_button_debounce_counter_cry_6),
            .clk(N__48476),
            .ce(),
            .sr(N__45714));
    defparam button_debounce_counter_7_LC_16_13_6.C_ON=1'b1;
    defparam button_debounce_counter_7_LC_16_13_6.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_7_LC_16_13_6.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_7_LC_16_13_6 (
            .in0(N__49193),
            .in1(N__38815),
            .in2(_gnd_net_),
            .in3(N__35021),
            .lcout(button_debounce_counterZ0Z_7),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_6),
            .carryout(un1_button_debounce_counter_cry_7),
            .clk(N__48476),
            .ce(),
            .sr(N__45714));
    defparam button_debounce_counter_8_LC_16_13_7.C_ON=1'b1;
    defparam button_debounce_counter_8_LC_16_13_7.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_8_LC_16_13_7.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_8_LC_16_13_7 (
            .in0(N__49431),
            .in1(N__38779),
            .in2(_gnd_net_),
            .in3(N__35018),
            .lcout(button_debounce_counterZ0Z_8),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_7),
            .carryout(un1_button_debounce_counter_cry_8),
            .clk(N__48476),
            .ce(),
            .sr(N__45714));
    defparam button_debounce_counter_9_LC_16_14_0.C_ON=1'b1;
    defparam button_debounce_counter_9_LC_16_14_0.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_9_LC_16_14_0.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_9_LC_16_14_0 (
            .in0(N__49295),
            .in1(N__38830),
            .in2(_gnd_net_),
            .in3(N__35015),
            .lcout(button_debounce_counterZ0Z_9),
            .ltout(),
            .carryin(bfn_16_14_0_),
            .carryout(un1_button_debounce_counter_cry_9),
            .clk(N__48480),
            .ce(),
            .sr(N__45715));
    defparam button_debounce_counter_10_LC_16_14_1.C_ON=1'b1;
    defparam button_debounce_counter_10_LC_16_14_1.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_10_LC_16_14_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_10_LC_16_14_1 (
            .in0(N__49288),
            .in1(N__38794),
            .in2(_gnd_net_),
            .in3(N__35195),
            .lcout(button_debounce_counterZ0Z_10),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_9),
            .carryout(un1_button_debounce_counter_cry_10),
            .clk(N__48480),
            .ce(),
            .sr(N__45715));
    defparam button_debounce_counter_11_LC_16_14_2.C_ON=1'b1;
    defparam button_debounce_counter_11_LC_16_14_2.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_11_LC_16_14_2.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_11_LC_16_14_2 (
            .in0(N__49292),
            .in1(N__38857),
            .in2(_gnd_net_),
            .in3(N__35192),
            .lcout(button_debounce_counterZ0Z_11),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_10),
            .carryout(un1_button_debounce_counter_cry_11),
            .clk(N__48480),
            .ce(),
            .sr(N__45715));
    defparam button_debounce_counter_12_LC_16_14_3.C_ON=1'b1;
    defparam button_debounce_counter_12_LC_16_14_3.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_12_LC_16_14_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_12_LC_16_14_3 (
            .in0(N__49289),
            .in1(N__38890),
            .in2(_gnd_net_),
            .in3(N__35189),
            .lcout(button_debounce_counterZ0Z_12),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_11),
            .carryout(un1_button_debounce_counter_cry_12),
            .clk(N__48480),
            .ce(),
            .sr(N__45715));
    defparam button_debounce_counter_13_LC_16_14_4.C_ON=1'b1;
    defparam button_debounce_counter_13_LC_16_14_4.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_13_LC_16_14_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_13_LC_16_14_4 (
            .in0(N__49293),
            .in1(N__38905),
            .in2(_gnd_net_),
            .in3(N__35186),
            .lcout(button_debounce_counterZ0Z_13),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_12),
            .carryout(un1_button_debounce_counter_cry_13),
            .clk(N__48480),
            .ce(),
            .sr(N__45715));
    defparam button_debounce_counter_14_LC_16_14_5.C_ON=1'b1;
    defparam button_debounce_counter_14_LC_16_14_5.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_14_LC_16_14_5.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_14_LC_16_14_5 (
            .in0(N__49290),
            .in1(N__38872),
            .in2(_gnd_net_),
            .in3(N__35183),
            .lcout(button_debounce_counterZ0Z_14),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_13),
            .carryout(un1_button_debounce_counter_cry_14),
            .clk(N__48480),
            .ce(),
            .sr(N__45715));
    defparam button_debounce_counter_15_LC_16_14_6.C_ON=1'b1;
    defparam button_debounce_counter_15_LC_16_14_6.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_15_LC_16_14_6.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_15_LC_16_14_6 (
            .in0(N__49294),
            .in1(N__35179),
            .in2(_gnd_net_),
            .in3(N__35165),
            .lcout(button_debounce_counterZ0Z_15),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_14),
            .carryout(un1_button_debounce_counter_cry_15),
            .clk(N__48480),
            .ce(),
            .sr(N__45715));
    defparam button_debounce_counter_16_LC_16_14_7.C_ON=1'b1;
    defparam button_debounce_counter_16_LC_16_14_7.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_16_LC_16_14_7.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_16_LC_16_14_7 (
            .in0(N__49291),
            .in1(N__35158),
            .in2(_gnd_net_),
            .in3(N__35144),
            .lcout(button_debounce_counterZ0Z_16),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_15),
            .carryout(un1_button_debounce_counter_cry_16),
            .clk(N__48480),
            .ce(),
            .sr(N__45715));
    defparam button_debounce_counter_17_LC_16_15_0.C_ON=1'b1;
    defparam button_debounce_counter_17_LC_16_15_0.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_17_LC_16_15_0.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_17_LC_16_15_0 (
            .in0(N__49302),
            .in1(N__35140),
            .in2(_gnd_net_),
            .in3(N__35126),
            .lcout(button_debounce_counterZ0Z_17),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(un1_button_debounce_counter_cry_17),
            .clk(N__48483),
            .ce(),
            .sr(N__45716));
    defparam button_debounce_counter_18_LC_16_15_1.C_ON=1'b1;
    defparam button_debounce_counter_18_LC_16_15_1.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_18_LC_16_15_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_18_LC_16_15_1 (
            .in0(N__49305),
            .in1(N__35123),
            .in2(_gnd_net_),
            .in3(N__35111),
            .lcout(button_debounce_counterZ0Z_18),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_17),
            .carryout(un1_button_debounce_counter_cry_18),
            .clk(N__48483),
            .ce(),
            .sr(N__45716));
    defparam button_debounce_counter_19_LC_16_15_2.C_ON=1'b1;
    defparam button_debounce_counter_19_LC_16_15_2.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_19_LC_16_15_2.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_19_LC_16_15_2 (
            .in0(N__49303),
            .in1(N__35360),
            .in2(_gnd_net_),
            .in3(N__35348),
            .lcout(button_debounce_counterZ0Z_19),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_18),
            .carryout(un1_button_debounce_counter_cry_19),
            .clk(N__48483),
            .ce(),
            .sr(N__45716));
    defparam button_debounce_counter_20_LC_16_15_3.C_ON=1'b1;
    defparam button_debounce_counter_20_LC_16_15_3.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_20_LC_16_15_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_20_LC_16_15_3 (
            .in0(N__49306),
            .in1(N__35345),
            .in2(_gnd_net_),
            .in3(N__35333),
            .lcout(button_debounce_counterZ0Z_20),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_19),
            .carryout(un1_button_debounce_counter_cry_20),
            .clk(N__48483),
            .ce(),
            .sr(N__45716));
    defparam button_debounce_counter_21_LC_16_15_4.C_ON=1'b1;
    defparam button_debounce_counter_21_LC_16_15_4.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_21_LC_16_15_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_21_LC_16_15_4 (
            .in0(N__49304),
            .in1(N__35329),
            .in2(_gnd_net_),
            .in3(N__35315),
            .lcout(button_debounce_counterZ0Z_21),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_20),
            .carryout(un1_button_debounce_counter_cry_21),
            .clk(N__48483),
            .ce(),
            .sr(N__45716));
    defparam button_debounce_counter_22_LC_16_15_5.C_ON=1'b1;
    defparam button_debounce_counter_22_LC_16_15_5.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_22_LC_16_15_5.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_22_LC_16_15_5 (
            .in0(N__49307),
            .in1(N__35305),
            .in2(_gnd_net_),
            .in3(N__35291),
            .lcout(button_debounce_counterZ0Z_22),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_21),
            .carryout(un1_button_debounce_counter_cry_22),
            .clk(N__48483),
            .ce(),
            .sr(N__45716));
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_0_LC_16_15_6.C_ON=1'b1;
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_0_LC_16_15_6.SEQ_MODE=4'b0000;
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_0_LC_16_15_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_button_debounce_counter_cry_22_c_THRU_CRY_0_LC_16_15_6 (
            .in0(_gnd_net_),
            .in1(N__52510),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_22),
            .carryout(un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_1_LC_16_15_7.C_ON=1'b1;
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_1_LC_16_15_7.SEQ_MODE=4'b0000;
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_1_LC_16_15_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_button_debounce_counter_cry_22_c_THRU_CRY_1_LC_16_15_7 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__52586),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO),
            .carryout(un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam button_debounce_counter_esr_23_LC_16_16_0.C_ON=1'b0;
    defparam button_debounce_counter_esr_23_LC_16_16_0.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_esr_23_LC_16_16_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 button_debounce_counter_esr_23_LC_16_16_0 (
            .in0(_gnd_net_),
            .in1(N__35284),
            .in2(_gnd_net_),
            .in3(N__35288),
            .lcout(button_debounce_counterZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48486),
            .ce(N__35270),
            .sr(N__45717));
    defparam sRAM_ADD_5_LC_16_17_0.C_ON=1'b0;
    defparam sRAM_ADD_5_LC_16_17_0.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_5_LC_16_17_0.LUT_INIT=16'b1110110001001100;
    LogicCell40 sRAM_ADD_5_LC_16_17_0 (
            .in0(N__43344),
            .in1(N__35255),
            .in2(N__43491),
            .in3(N__35237),
            .lcout(RAM_ADD_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52269),
            .ce(N__43218),
            .sr(_gnd_net_));
    defparam sRAM_ADD_0_LC_16_17_1.C_ON=1'b0;
    defparam sRAM_ADD_0_LC_16_17_1.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_0_LC_16_17_1.LUT_INIT=16'b1110001010101010;
    LogicCell40 sRAM_ADD_0_LC_16_17_1 (
            .in0(N__35909),
            .in1(N__43450),
            .in2(N__35891),
            .in3(N__43337),
            .lcout(RAM_ADD_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52269),
            .ce(N__43218),
            .sr(_gnd_net_));
    defparam sRAM_ADD_10_LC_16_17_2.C_ON=1'b0;
    defparam sRAM_ADD_10_LC_16_17_2.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_10_LC_16_17_2.LUT_INIT=16'b1110110001001100;
    LogicCell40 sRAM_ADD_10_LC_16_17_2 (
            .in0(N__43338),
            .in1(N__35846),
            .in2(N__43488),
            .in3(N__35828),
            .lcout(RAM_ADD_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52269),
            .ce(N__43218),
            .sr(_gnd_net_));
    defparam sRAM_ADD_11_LC_16_17_3.C_ON=1'b0;
    defparam sRAM_ADD_11_LC_16_17_3.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_11_LC_16_17_3.LUT_INIT=16'b1110001010101010;
    LogicCell40 sRAM_ADD_11_LC_16_17_3 (
            .in0(N__35774),
            .in1(N__43454),
            .in2(N__35756),
            .in3(N__43339),
            .lcout(RAM_ADD_c_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52269),
            .ce(N__43218),
            .sr(_gnd_net_));
    defparam sRAM_ADD_12_LC_16_17_4.C_ON=1'b0;
    defparam sRAM_ADD_12_LC_16_17_4.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_12_LC_16_17_4.LUT_INIT=16'b1101111110000000;
    LogicCell40 sRAM_ADD_12_LC_16_17_4 (
            .in0(N__43340),
            .in1(N__35705),
            .in2(N__43489),
            .in3(N__35678),
            .lcout(RAM_ADD_c_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52269),
            .ce(N__43218),
            .sr(_gnd_net_));
    defparam sRAM_ADD_13_LC_16_17_5.C_ON=1'b0;
    defparam sRAM_ADD_13_LC_16_17_5.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_13_LC_16_17_5.LUT_INIT=16'b1110001010101010;
    LogicCell40 sRAM_ADD_13_LC_16_17_5 (
            .in0(N__35639),
            .in1(N__43458),
            .in2(N__35621),
            .in3(N__43341),
            .lcout(RAM_ADD_c_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52269),
            .ce(N__43218),
            .sr(_gnd_net_));
    defparam sRAM_ADD_14_LC_16_17_6.C_ON=1'b0;
    defparam sRAM_ADD_14_LC_16_17_6.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_14_LC_16_17_6.LUT_INIT=16'b1101111110000000;
    LogicCell40 sRAM_ADD_14_LC_16_17_6 (
            .in0(N__43342),
            .in1(N__35576),
            .in2(N__43490),
            .in3(N__35549),
            .lcout(RAM_ADD_c_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52269),
            .ce(N__43218),
            .sr(_gnd_net_));
    defparam sRAM_ADD_15_LC_16_17_7.C_ON=1'b0;
    defparam sRAM_ADD_15_LC_16_17_7.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_15_LC_16_17_7.LUT_INIT=16'b1110001010101010;
    LogicCell40 sRAM_ADD_15_LC_16_17_7 (
            .in0(N__35504),
            .in1(N__43462),
            .in2(N__35486),
            .in3(N__43343),
            .lcout(RAM_ADD_c_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52269),
            .ce(N__43218),
            .sr(_gnd_net_));
    defparam sRAM_ADD_16_LC_16_18_0.C_ON=1'b0;
    defparam sRAM_ADD_16_LC_16_18_0.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_16_LC_16_18_0.LUT_INIT=16'b1110001010101010;
    LogicCell40 sRAM_ADD_16_LC_16_18_0 (
            .in0(N__35432),
            .in1(N__43492),
            .in2(N__35414),
            .in3(N__43348),
            .lcout(RAM_ADD_c_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52279),
            .ce(N__43226),
            .sr(_gnd_net_));
    defparam sRAM_ADD_17_LC_16_18_1.C_ON=1'b0;
    defparam sRAM_ADD_17_LC_16_18_1.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_17_LC_16_18_1.LUT_INIT=16'b1101100011110000;
    LogicCell40 sRAM_ADD_17_LC_16_18_1 (
            .in0(N__43349),
            .in1(N__36404),
            .in2(N__36377),
            .in3(N__43496),
            .lcout(RAM_ADD_c_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52279),
            .ce(N__43226),
            .sr(_gnd_net_));
    defparam sRAM_ADD_18_LC_16_18_2.C_ON=1'b0;
    defparam sRAM_ADD_18_LC_16_18_2.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_18_LC_16_18_2.LUT_INIT=16'b1011100011110000;
    LogicCell40 sRAM_ADD_18_LC_16_18_2 (
            .in0(N__36338),
            .in1(N__43493),
            .in2(N__36311),
            .in3(N__43350),
            .lcout(RAM_ADD_c_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52279),
            .ce(N__43226),
            .sr(_gnd_net_));
    defparam sRAM_ADD_9_LC_16_18_3.C_ON=1'b0;
    defparam sRAM_ADD_9_LC_16_18_3.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_9_LC_16_18_3.LUT_INIT=16'b1101100011110000;
    LogicCell40 sRAM_ADD_9_LC_16_18_3 (
            .in0(N__43355),
            .in1(N__36266),
            .in2(N__36239),
            .in3(N__43499),
            .lcout(RAM_ADD_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52279),
            .ce(N__43226),
            .sr(_gnd_net_));
    defparam sRAM_ADD_7_LC_16_18_4.C_ON=1'b0;
    defparam sRAM_ADD_7_LC_16_18_4.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_7_LC_16_18_4.LUT_INIT=16'b1011100011110000;
    LogicCell40 sRAM_ADD_7_LC_16_18_4 (
            .in0(N__36197),
            .in1(N__43495),
            .in2(N__36170),
            .in3(N__43354),
            .lcout(RAM_ADD_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52279),
            .ce(N__43226),
            .sr(_gnd_net_));
    defparam sRAM_ADD_2_LC_16_18_5.C_ON=1'b0;
    defparam sRAM_ADD_2_LC_16_18_5.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_2_LC_16_18_5.LUT_INIT=16'b1110010011001100;
    LogicCell40 sRAM_ADD_2_LC_16_18_5 (
            .in0(N__43352),
            .in1(N__36134),
            .in2(N__36119),
            .in3(N__43497),
            .lcout(RAM_ADD_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52279),
            .ce(N__43226),
            .sr(_gnd_net_));
    defparam sRAM_ADD_1_LC_16_18_6.C_ON=1'b0;
    defparam sRAM_ADD_1_LC_16_18_6.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_1_LC_16_18_6.LUT_INIT=16'b1011100011110000;
    LogicCell40 sRAM_ADD_1_LC_16_18_6 (
            .in0(N__36074),
            .in1(N__43494),
            .in2(N__36047),
            .in3(N__43351),
            .lcout(RAM_ADD_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52279),
            .ce(N__43226),
            .sr(_gnd_net_));
    defparam sRAM_ADD_6_LC_16_18_7.C_ON=1'b0;
    defparam sRAM_ADD_6_LC_16_18_7.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_6_LC_16_18_7.LUT_INIT=16'b1101100011110000;
    LogicCell40 sRAM_ADD_6_LC_16_18_7 (
            .in0(N__43353),
            .in1(N__36017),
            .in2(N__35990),
            .in3(N__43498),
            .lcout(RAM_ADD_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52279),
            .ce(N__43226),
            .sr(_gnd_net_));
    defparam RAM_DATA_1_4_LC_16_20_0.C_ON=1'b0;
    defparam RAM_DATA_1_4_LC_16_20_0.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_4_LC_16_20_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 RAM_DATA_1_4_LC_16_20_0 (
            .in0(N__35951),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RAM_DATA_1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52301),
            .ce(N__51895),
            .sr(N__51650));
    defparam sDAC_mem_pointer_6_LC_17_1_0.C_ON=1'b0;
    defparam sDAC_mem_pointer_6_LC_17_1_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_6_LC_17_1_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_pointer_6_LC_17_1_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_mem_pointerZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48447),
            .ce(N__43957),
            .sr(N__51823));
    defparam sDAC_mem_pointer_7_LC_17_1_1.C_ON=1'b0;
    defparam sDAC_mem_pointer_7_LC_17_1_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_7_LC_17_1_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_pointer_7_LC_17_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_mem_pointerZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48447),
            .ce(N__43957),
            .sr(N__51823));
    defparam sDAC_mem_4_2_LC_17_3_0.C_ON=1'b0;
    defparam sDAC_mem_4_2_LC_17_3_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_2_LC_17_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_2_LC_17_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47438),
            .lcout(sDAC_mem_4Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52281),
            .ce(N__42626),
            .sr(N__51813));
    defparam sDAC_mem_4_5_LC_17_3_1.C_ON=1'b0;
    defparam sDAC_mem_4_5_LC_17_3_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_5_LC_17_3_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_5_LC_17_3_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45104),
            .lcout(sDAC_mem_4Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52281),
            .ce(N__42626),
            .sr(N__51813));
    defparam sDAC_mem_4_7_LC_17_3_2.C_ON=1'b0;
    defparam sDAC_mem_4_7_LC_17_3_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_7_LC_17_3_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_7_LC_17_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50055),
            .lcout(sDAC_mem_4Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52281),
            .ce(N__42626),
            .sr(N__51813));
    defparam sDAC_mem_20_0_LC_17_4_0.C_ON=1'b0;
    defparam sDAC_mem_20_0_LC_17_4_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_0_LC_17_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_0_LC_17_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46386),
            .lcout(sDAC_mem_20Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52270),
            .ce(N__36638),
            .sr(N__51807));
    defparam sDAC_mem_20_1_LC_17_4_1.C_ON=1'b0;
    defparam sDAC_mem_20_1_LC_17_4_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_1_LC_17_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_1_LC_17_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51054),
            .lcout(sDAC_mem_20Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52270),
            .ce(N__36638),
            .sr(N__51807));
    defparam sDAC_mem_20_2_LC_17_4_2.C_ON=1'b0;
    defparam sDAC_mem_20_2_LC_17_4_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_2_LC_17_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_2_LC_17_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47437),
            .lcout(sDAC_mem_20Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52270),
            .ce(N__36638),
            .sr(N__51807));
    defparam sDAC_mem_20_3_LC_17_4_3.C_ON=1'b0;
    defparam sDAC_mem_20_3_LC_17_4_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_3_LC_17_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_3_LC_17_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46752),
            .lcout(sDAC_mem_20Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52270),
            .ce(N__36638),
            .sr(N__51807));
    defparam sDAC_mem_20_4_LC_17_4_4.C_ON=1'b0;
    defparam sDAC_mem_20_4_LC_17_4_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_4_LC_17_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_4_LC_17_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45558),
            .lcout(sDAC_mem_20Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52270),
            .ce(N__36638),
            .sr(N__51807));
    defparam sDAC_mem_20_7_LC_17_4_5.C_ON=1'b0;
    defparam sDAC_mem_20_7_LC_17_4_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_7_LC_17_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_7_LC_17_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49865),
            .lcout(sDAC_mem_20Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52270),
            .ce(N__36638),
            .sr(N__51807));
    defparam sDAC_mem_6_0_LC_17_5_0.C_ON=1'b0;
    defparam sDAC_mem_6_0_LC_17_5_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_0_LC_17_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_0_LC_17_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46388),
            .lcout(sDAC_mem_6Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52258),
            .ce(N__36554),
            .sr(N__51798));
    defparam sDAC_mem_6_1_LC_17_5_1.C_ON=1'b0;
    defparam sDAC_mem_6_1_LC_17_5_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_1_LC_17_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_1_LC_17_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51052),
            .lcout(sDAC_mem_6Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52258),
            .ce(N__36554),
            .sr(N__51798));
    defparam sDAC_mem_6_4_LC_17_5_2.C_ON=1'b0;
    defparam sDAC_mem_6_4_LC_17_5_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_4_LC_17_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_4_LC_17_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45350),
            .lcout(sDAC_mem_6Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52258),
            .ce(N__36554),
            .sr(N__51798));
    defparam sDAC_mem_6_7_LC_17_5_3.C_ON=1'b0;
    defparam sDAC_mem_6_7_LC_17_5_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_7_LC_17_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_7_LC_17_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49847),
            .lcout(sDAC_mem_6Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52258),
            .ce(N__36554),
            .sr(N__51798));
    defparam sDAC_mem_23_0_LC_17_6_0.C_ON=1'b0;
    defparam sDAC_mem_23_0_LC_17_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_0_LC_17_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_0_LC_17_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46387),
            .lcout(sDAC_mem_23Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52248),
            .ce(N__36701),
            .sr(N__51784));
    defparam sDAC_mem_23_1_LC_17_6_1.C_ON=1'b0;
    defparam sDAC_mem_23_1_LC_17_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_1_LC_17_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_1_LC_17_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51055),
            .lcout(sDAC_mem_23Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52248),
            .ce(N__36701),
            .sr(N__51784));
    defparam sDAC_mem_23_2_LC_17_6_2.C_ON=1'b0;
    defparam sDAC_mem_23_2_LC_17_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_2_LC_17_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_2_LC_17_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47446),
            .lcout(sDAC_mem_23Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52248),
            .ce(N__36701),
            .sr(N__51784));
    defparam sDAC_mem_23_3_LC_17_6_3.C_ON=1'b0;
    defparam sDAC_mem_23_3_LC_17_6_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_3_LC_17_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_3_LC_17_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46858),
            .lcout(sDAC_mem_23Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52248),
            .ce(N__36701),
            .sr(N__51784));
    defparam sDAC_mem_23_4_LC_17_6_4.C_ON=1'b0;
    defparam sDAC_mem_23_4_LC_17_6_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_4_LC_17_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_4_LC_17_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45559),
            .lcout(sDAC_mem_23Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52248),
            .ce(N__36701),
            .sr(N__51784));
    defparam sDAC_mem_23_5_LC_17_6_5.C_ON=1'b0;
    defparam sDAC_mem_23_5_LC_17_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_5_LC_17_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_5_LC_17_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45100),
            .lcout(sDAC_mem_23Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52248),
            .ce(N__36701),
            .sr(N__51784));
    defparam sDAC_mem_23_6_LC_17_6_6.C_ON=1'b0;
    defparam sDAC_mem_23_6_LC_17_6_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_6_LC_17_6_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_23_6_LC_17_6_6 (
            .in0(N__50485),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_23Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52248),
            .ce(N__36701),
            .sr(N__51784));
    defparam sDAC_mem_23_7_LC_17_6_7.C_ON=1'b0;
    defparam sDAC_mem_23_7_LC_17_6_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_7_LC_17_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_7_LC_17_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49866),
            .lcout(sDAC_mem_23Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52248),
            .ce(N__36701),
            .sr(N__51784));
    defparam sDAC_mem_32_3_LC_17_7_0.C_ON=1'b0;
    defparam sDAC_mem_32_3_LC_17_7_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_3_LC_17_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_3_LC_17_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46920),
            .lcout(sDAC_mem_32Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52236),
            .ce(N__41258),
            .sr(N__51772));
    defparam sDAC_data_RNO_26_6_LC_17_7_1.C_ON=1'b0;
    defparam sDAC_data_RNO_26_6_LC_17_7_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_6_LC_17_7_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_26_6_LC_17_7_1 (
            .in0(N__42422),
            .in1(N__44360),
            .in2(_gnd_net_),
            .in3(N__44102),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_6_LC_17_7_2.C_ON=1'b0;
    defparam sDAC_data_RNO_14_6_LC_17_7_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_6_LC_17_7_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 sDAC_data_RNO_14_6_LC_17_7_2 (
            .in0(_gnd_net_),
            .in1(N__42189),
            .in2(N__36683),
            .in3(N__36680),
            .lcout(sDAC_data_RNO_14Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_26_7_LC_17_7_3.C_ON=1'b0;
    defparam sDAC_data_RNO_26_7_LC_17_7_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_7_LC_17_7_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_26_7_LC_17_7_3 (
            .in0(N__42423),
            .in1(N__44093),
            .in2(_gnd_net_),
            .in3(N__44348),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_7_LC_17_7_4.C_ON=1'b0;
    defparam sDAC_data_RNO_14_7_LC_17_7_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_7_LC_17_7_4.LUT_INIT=16'b1111001111000000;
    LogicCell40 sDAC_data_RNO_14_7_LC_17_7_4 (
            .in0(_gnd_net_),
            .in1(N__42190),
            .in2(N__36884),
            .in3(N__36869),
            .lcout(sDAC_data_RNO_14Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_32_4_LC_17_7_5.C_ON=1'b0;
    defparam sDAC_mem_32_4_LC_17_7_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_4_LC_17_7_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_32_4_LC_17_7_5 (
            .in0(N__45592),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_32Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52236),
            .ce(N__41258),
            .sr(N__51772));
    defparam sDAC_data_RNO_26_8_LC_17_7_6.C_ON=1'b0;
    defparam sDAC_data_RNO_26_8_LC_17_7_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_8_LC_17_7_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_26_8_LC_17_7_6 (
            .in0(N__42431),
            .in1(N__44336),
            .in2(_gnd_net_),
            .in3(N__44084),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_8_LC_17_7_7.C_ON=1'b0;
    defparam sDAC_data_RNO_14_8_LC_17_7_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_8_LC_17_7_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 sDAC_data_RNO_14_8_LC_17_7_7 (
            .in0(N__42191),
            .in1(_gnd_net_),
            .in2(N__36863),
            .in3(N__39632),
            .lcout(sDAC_data_RNO_14Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_9_0_LC_17_8_0.C_ON=1'b0;
    defparam sDAC_mem_9_0_LC_17_8_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_0_LC_17_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_9_0_LC_17_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46352),
            .lcout(sDAC_mem_9Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52226),
            .ce(N__39818),
            .sr(N__51759));
    defparam sDAC_mem_9_1_LC_17_8_1.C_ON=1'b0;
    defparam sDAC_mem_9_1_LC_17_8_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_1_LC_17_8_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_9_1_LC_17_8_1 (
            .in0(N__51070),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_9Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52226),
            .ce(N__39818),
            .sr(N__51759));
    defparam sDAC_mem_9_2_LC_17_8_2.C_ON=1'b0;
    defparam sDAC_mem_9_2_LC_17_8_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_2_LC_17_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_9_2_LC_17_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47439),
            .lcout(sDAC_mem_9Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52226),
            .ce(N__39818),
            .sr(N__51759));
    defparam sDAC_mem_9_3_LC_17_8_3.C_ON=1'b0;
    defparam sDAC_mem_9_3_LC_17_8_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_3_LC_17_8_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_9_3_LC_17_8_3 (
            .in0(N__46859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_9Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52226),
            .ce(N__39818),
            .sr(N__51759));
    defparam sDAC_mem_9_4_LC_17_8_4.C_ON=1'b0;
    defparam sDAC_mem_9_4_LC_17_8_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_4_LC_17_8_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_9_4_LC_17_8_4 (
            .in0(N__45560),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_9Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52226),
            .ce(N__39818),
            .sr(N__51759));
    defparam sDAC_mem_9_5_LC_17_8_5.C_ON=1'b0;
    defparam sDAC_mem_9_5_LC_17_8_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_5_LC_17_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_9_5_LC_17_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45103),
            .lcout(sDAC_mem_9Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52226),
            .ce(N__39818),
            .sr(N__51759));
    defparam sDAC_mem_9_6_LC_17_8_6.C_ON=1'b0;
    defparam sDAC_mem_9_6_LC_17_8_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_6_LC_17_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_9_6_LC_17_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50487),
            .lcout(sDAC_mem_9Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52226),
            .ce(N__39818),
            .sr(N__51759));
    defparam sDAC_mem_9_7_LC_17_8_7.C_ON=1'b0;
    defparam sDAC_mem_9_7_LC_17_8_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_7_LC_17_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_9_7_LC_17_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49867),
            .lcout(sDAC_mem_9Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52226),
            .ce(N__39818),
            .sr(N__51759));
    defparam sDAC_data_RNO_19_9_LC_17_9_0.C_ON=1'b0;
    defparam sDAC_data_RNO_19_9_LC_17_9_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_9_LC_17_9_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_9_LC_17_9_0 (
            .in0(N__41841),
            .in1(N__37016),
            .in2(_gnd_net_),
            .in3(N__37007),
            .lcout(sDAC_data_RNO_19Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_9_LC_17_9_1.C_ON=1'b0;
    defparam sDAC_data_RNO_18_9_LC_17_9_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_9_LC_17_9_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_9_LC_17_9_1 (
            .in0(N__42142),
            .in1(N__44609),
            .in2(_gnd_net_),
            .in3(N__36971),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_9_LC_17_9_2.C_ON=1'b0;
    defparam sDAC_data_RNO_9_9_LC_17_9_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_9_LC_17_9_2.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_9_9_LC_17_9_2 (
            .in0(N__38096),
            .in1(N__38460),
            .in2(N__36992),
            .in3(N__36989),
            .lcout(sDAC_data_2_24_ns_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_12_6_LC_17_9_3.C_ON=1'b0;
    defparam sDAC_mem_12_6_LC_17_9_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_6_LC_17_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_6_LC_17_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50488),
            .lcout(sDAC_mem_12Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52220),
            .ce(N__36964),
            .sr(N__51747));
    defparam sDAC_mem_pointer_RNIAIV21_3_LC_17_9_4.C_ON=1'b0;
    defparam sDAC_mem_pointer_RNIAIV21_3_LC_17_9_4.SEQ_MODE=4'b0000;
    defparam sDAC_mem_pointer_RNIAIV21_3_LC_17_9_4.LUT_INIT=16'b1110101000000000;
    LogicCell40 sDAC_mem_pointer_RNIAIV21_3_LC_17_9_4 (
            .in0(N__38095),
            .in1(N__38459),
            .in2(N__42074),
            .in3(N__37305),
            .lcout(),
            .ltout(op_le_op_le_un15_sdacdynlt4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_pointer_RNI4LV52_4_LC_17_9_5.C_ON=1'b0;
    defparam sDAC_mem_pointer_RNI4LV52_4_LC_17_9_5.SEQ_MODE=4'b0000;
    defparam sDAC_mem_pointer_RNI4LV52_4_LC_17_9_5.LUT_INIT=16'b0011011100000000;
    LogicCell40 sDAC_mem_pointer_RNI4LV52_4_LC_17_9_5 (
            .in0(N__37390),
            .in1(N__42411),
            .in2(N__36902),
            .in3(N__37172),
            .lcout(un17_sdacdyn_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_pointer_RNIF3GH_6_LC_17_9_6.C_ON=1'b0;
    defparam sDAC_mem_pointer_RNIF3GH_6_LC_17_9_6.SEQ_MODE=4'b0000;
    defparam sDAC_mem_pointer_RNIF3GH_6_LC_17_9_6.LUT_INIT=16'b0000000000110011;
    LogicCell40 sDAC_mem_pointer_RNIF3GH_6_LC_17_9_6 (
            .in0(_gnd_net_),
            .in1(N__37196),
            .in2(_gnd_net_),
            .in3(N__37181),
            .lcout(un17_sdacdyn_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_26_3_LC_17_9_7.C_ON=1'b0;
    defparam sDAC_data_RNO_26_3_LC_17_9_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_3_LC_17_9_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_26_3_LC_17_9_7 (
            .in0(N__42421),
            .in1(N__44390),
            .in2(_gnd_net_),
            .in3(N__44135),
            .lcout(sDAC_data_RNO_26Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_5_LC_17_10_0.C_ON=1'b0;
    defparam sDAC_data_RNO_1_5_LC_17_10_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_5_LC_17_10_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_1_5_LC_17_10_0 (
            .in0(N__37166),
            .in1(N__41375),
            .in2(N__38196),
            .in3(N__37100),
            .lcout(),
            .ltout(sDAC_data_RNO_1Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_5_LC_17_10_1.C_ON=1'b0;
    defparam sDAC_data_RNO_0_5_LC_17_10_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_5_LC_17_10_1.LUT_INIT=16'b0101000011101110;
    LogicCell40 sDAC_data_RNO_0_5_LC_17_10_1 (
            .in0(N__37442),
            .in1(N__37154),
            .in2(N__37148),
            .in3(N__37046),
            .lcout(),
            .ltout(sDAC_data_2_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_5_LC_17_10_2.C_ON=1'b0;
    defparam sDAC_data_5_LC_17_10_2.SEQ_MODE=4'b1010;
    defparam sDAC_data_5_LC_17_10_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 sDAC_data_5_LC_17_10_2 (
            .in0(_gnd_net_),
            .in1(N__37145),
            .in2(N__37130),
            .in3(N__37631),
            .lcout(sDAC_dataZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48470),
            .ce(N__43947),
            .sr(N__51732));
    defparam sDAC_data_RNO_6_5_LC_17_10_3.C_ON=1'b0;
    defparam sDAC_data_RNO_6_5_LC_17_10_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_5_LC_17_10_3.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_6_5_LC_17_10_3 (
            .in0(N__38530),
            .in1(N__37106),
            .in2(N__38253),
            .in3(N__41288),
            .lcout(sDAC_data_2_14_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_5_LC_17_10_4.C_ON=1'b0;
    defparam sDAC_data_RNO_22_5_LC_17_10_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_5_LC_17_10_4.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_22_5_LC_17_10_4 (
            .in0(N__38506),
            .in1(N__37094),
            .in2(N__38195),
            .in3(N__37088),
            .lcout(),
            .ltout(sDAC_data_2_32_ns_1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_5_LC_17_10_5.C_ON=1'b0;
    defparam sDAC_data_RNO_10_5_LC_17_10_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_5_LC_17_10_5.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_10_5_LC_17_10_5 (
            .in0(N__37073),
            .in1(N__38091),
            .in2(N__37064),
            .in3(N__37061),
            .lcout(),
            .ltout(sDAC_data_RNO_10Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_5_LC_17_10_6.C_ON=1'b0;
    defparam sDAC_data_RNO_3_5_LC_17_10_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_5_LC_17_10_6.LUT_INIT=16'b0001010110011101;
    LogicCell40 sDAC_data_RNO_3_5_LC_17_10_6 (
            .in0(N__37334),
            .in1(N__37441),
            .in2(N__37049),
            .in3(N__37205),
            .lcout(sDAC_data_2_41_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_3_LC_17_11_0.C_ON=1'b0;
    defparam sDAC_data_RNO_1_3_LC_17_11_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_3_LC_17_11_0.LUT_INIT=16'b1100000010111011;
    LogicCell40 sDAC_data_RNO_1_3_LC_17_11_0 (
            .in0(N__37676),
            .in1(N__38177),
            .in2(N__41189),
            .in3(N__37244),
            .lcout(),
            .ltout(sDAC_data_RNO_1Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_3_LC_17_11_1.C_ON=1'b0;
    defparam sDAC_data_RNO_0_3_LC_17_11_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_3_LC_17_11_1.LUT_INIT=16'b0011000011101110;
    LogicCell40 sDAC_data_RNO_0_3_LC_17_11_1 (
            .in0(N__37664),
            .in1(N__37455),
            .in2(N__37658),
            .in3(N__37256),
            .lcout(),
            .ltout(sDAC_data_2_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_3_LC_17_11_2.C_ON=1'b0;
    defparam sDAC_data_3_LC_17_11_2.SEQ_MODE=4'b1010;
    defparam sDAC_data_3_LC_17_11_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 sDAC_data_3_LC_17_11_2 (
            .in0(N__37655),
            .in1(_gnd_net_),
            .in2(N__37640),
            .in3(N__37629),
            .lcout(sDAC_dataZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48473),
            .ce(N__43948),
            .sr(N__51720));
    defparam sDAC_data_RNO_10_3_LC_17_11_3.C_ON=1'b0;
    defparam sDAC_data_RNO_10_3_LC_17_11_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_3_LC_17_11_3.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_10_3_LC_17_11_3 (
            .in0(N__37511),
            .in1(N__37499),
            .in2(N__38232),
            .in3(N__37220),
            .lcout(),
            .ltout(sDAC_data_RNO_10Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_3_LC_17_11_4.C_ON=1'b0;
    defparam sDAC_data_RNO_3_3_LC_17_11_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_3_LC_17_11_4.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_3_3_LC_17_11_4 (
            .in0(N__37454),
            .in1(N__37335),
            .in2(N__37271),
            .in3(N__37268),
            .lcout(sDAC_data_2_41_ns_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_3_LC_17_11_5.C_ON=1'b0;
    defparam sDAC_data_RNO_6_3_LC_17_11_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_3_LC_17_11_5.LUT_INIT=16'b0101000101011011;
    LogicCell40 sDAC_data_RNO_6_3_LC_17_11_5 (
            .in0(N__38507),
            .in1(N__41054),
            .in2(N__38233),
            .in3(N__37250),
            .lcout(sDAC_data_2_14_ns_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_3_LC_17_11_6.C_ON=1'b0;
    defparam sDAC_data_RNO_22_3_LC_17_11_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_3_LC_17_11_6.LUT_INIT=16'b0000110100111101;
    LogicCell40 sDAC_data_RNO_22_3_LC_17_11_6 (
            .in0(N__37238),
            .in1(N__38170),
            .in2(N__38531),
            .in3(N__37226),
            .lcout(sDAC_data_2_32_ns_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_5_LC_17_12_0.C_ON=1'b0;
    defparam sDAC_data_RNO_11_5_LC_17_12_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_5_LC_17_12_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_11_5_LC_17_12_0 (
            .in0(N__37712),
            .in1(N__38579),
            .in2(N__38251),
            .in3(N__37214),
            .lcout(sDAC_data_RNO_11Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_5_LC_17_12_1.C_ON=1'b0;
    defparam sDAC_data_RNO_23_5_LC_17_12_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_5_LC_17_12_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_5_LC_17_12_1 (
            .in0(N__42036),
            .in1(N__38597),
            .in2(_gnd_net_),
            .in3(N__37814),
            .lcout(sDAC_data_RNO_23Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_30_6_LC_17_12_2.C_ON=1'b0;
    defparam sDAC_data_RNO_30_6_LC_17_12_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_6_LC_17_12_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 sDAC_data_RNO_30_6_LC_17_12_2 (
            .in0(N__38573),
            .in1(N__41345),
            .in2(_gnd_net_),
            .in3(N__42038),
            .lcout(),
            .ltout(sDAC_data_RNO_30Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_25_6_LC_17_12_3.C_ON=1'b0;
    defparam sDAC_data_RNO_25_6_LC_17_12_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_6_LC_17_12_3.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_25_6_LC_17_12_3 (
            .in0(N__38190),
            .in1(N__38511),
            .in2(N__38306),
            .in3(N__37682),
            .lcout(),
            .ltout(sDAC_data_2_39_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_6_LC_17_12_4.C_ON=1'b0;
    defparam sDAC_data_RNO_11_6_LC_17_12_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_6_LC_17_12_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_11_6_LC_17_12_4 (
            .in0(N__38194),
            .in1(N__37856),
            .in2(N__37844),
            .in3(N__37841),
            .lcout(sDAC_data_RNO_11Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_28_2_LC_17_12_5.C_ON=1'b0;
    defparam sDAC_mem_28_2_LC_17_12_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_2_LC_17_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_2_LC_17_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47492),
            .lcout(sDAC_mem_28Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52213),
            .ce(N__37806),
            .sr(N__51709));
    defparam sDAC_data_RNO_24_5_LC_17_12_6.C_ON=1'b0;
    defparam sDAC_data_RNO_24_5_LC_17_12_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_5_LC_17_12_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 sDAC_data_RNO_24_5_LC_17_12_6 (
            .in0(N__37739),
            .in1(N__37724),
            .in2(_gnd_net_),
            .in3(N__42037),
            .lcout(sDAC_data_RNO_24Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_31_6_LC_17_12_7.C_ON=1'b0;
    defparam sDAC_data_RNO_31_6_LC_17_12_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_6_LC_17_12_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_31_6_LC_17_12_7 (
            .in0(N__42035),
            .in1(N__37706),
            .in2(_gnd_net_),
            .in3(N__37694),
            .lcout(sDAC_data_RNO_31Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_c_LC_17_13_0 .C_ON=1'b1;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_c_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_c_LC_17_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_c_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__42787),
            .in2(N__42772),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_LUT4_0_LC_17_13_1 .C_ON=1'b1;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_LUT4_0_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_LUT4_0_LC_17_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_LUT4_0_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__42729),
            .in2(_gnd_net_),
            .in3(N__38672),
            .lcout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_LUT4_0_LC_17_13_2 .C_ON=1'b1;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_LUT4_0_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_LUT4_0_LC_17_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_LUT4_0_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__42678),
            .in2(_gnd_net_),
            .in3(N__38669),
            .lcout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_3_LC_17_13_3 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_3_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_3_LC_17_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_3_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(N__48303),
            .in2(_gnd_net_),
            .in3(N__38666),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3 ),
            .clk(N__48263),
            .ce(),
            .sr(N__51700));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_4_LC_17_13_4 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_4_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_4_LC_17_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_4_LC_17_13_4  (
            .in0(_gnd_net_),
            .in1(N__48324),
            .in2(_gnd_net_),
            .in3(N__38663),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4 ),
            .clk(N__48263),
            .ce(),
            .sr(N__51700));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_5_LC_17_13_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_5_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_5_LC_17_13_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_5_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(N__38653),
            .in2(_gnd_net_),
            .in3(N__38660),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48263),
            .ce(),
            .sr(N__51700));
    defparam sDAC_mem_17_0_LC_17_14_0.C_ON=1'b0;
    defparam sDAC_mem_17_0_LC_17_14_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_0_LC_17_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_0_LC_17_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46293),
            .lcout(sDAC_mem_17Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52227),
            .ce(N__39920),
            .sr(N__51691));
    defparam sDAC_mem_17_1_LC_17_14_1.C_ON=1'b0;
    defparam sDAC_mem_17_1_LC_17_14_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_1_LC_17_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_1_LC_17_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50880),
            .lcout(sDAC_mem_17Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52227),
            .ce(N__39920),
            .sr(N__51691));
    defparam sDAC_mem_17_2_LC_17_14_2.C_ON=1'b0;
    defparam sDAC_mem_17_2_LC_17_14_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_2_LC_17_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_2_LC_17_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47511),
            .lcout(sDAC_mem_17Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52227),
            .ce(N__39920),
            .sr(N__51691));
    defparam sDAC_mem_17_3_LC_17_14_3.C_ON=1'b0;
    defparam sDAC_mem_17_3_LC_17_14_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_3_LC_17_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_3_LC_17_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46907),
            .lcout(sDAC_mem_17Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52227),
            .ce(N__39920),
            .sr(N__51691));
    defparam sDAC_mem_17_4_LC_17_14_4.C_ON=1'b0;
    defparam sDAC_mem_17_4_LC_17_14_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_4_LC_17_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_4_LC_17_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45611),
            .lcout(sDAC_mem_17Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52227),
            .ce(N__39920),
            .sr(N__51691));
    defparam sDAC_mem_17_5_LC_17_14_5.C_ON=1'b0;
    defparam sDAC_mem_17_5_LC_17_14_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_5_LC_17_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_5_LC_17_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45107),
            .lcout(sDAC_mem_17Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52227),
            .ce(N__39920),
            .sr(N__51691));
    defparam sDAC_mem_17_6_LC_17_14_6.C_ON=1'b0;
    defparam sDAC_mem_17_6_LC_17_14_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_6_LC_17_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_6_LC_17_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50527),
            .lcout(sDAC_mem_17Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52227),
            .ce(N__39920),
            .sr(N__51691));
    defparam sDAC_mem_17_7_LC_17_14_7.C_ON=1'b0;
    defparam sDAC_mem_17_7_LC_17_14_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_7_LC_17_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_7_LC_17_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49874),
            .lcout(sDAC_mem_17Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52227),
            .ce(N__39920),
            .sr(N__51691));
    defparam spi_data_miso_6_LC_17_15_6.C_ON=1'b0;
    defparam spi_data_miso_6_LC_17_15_6.SEQ_MODE=4'b1010;
    defparam spi_data_miso_6_LC_17_15_6.LUT_INIT=16'b0000000011100010;
    LogicCell40 spi_data_miso_6_LC_17_15_6 (
            .in0(N__38951),
            .in1(N__43767),
            .in2(N__38930),
            .in3(N__48946),
            .lcout(spi_data_misoZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52237),
            .ce(N__43687),
            .sr(N__51685));
    defparam sbuttonModeStatus_RNO_6_LC_17_16_0.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_6_LC_17_16_0.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_6_LC_17_16_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_6_LC_17_16_0 (
            .in0(N__38906),
            .in1(N__38891),
            .in2(N__38876),
            .in3(N__38858),
            .lcout(sbuttonModeStatus_0_sqmuxa_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_7_LC_17_16_1.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_7_LC_17_16_1.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_7_LC_17_16_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_7_LC_17_16_1 (
            .in0(N__38834),
            .in1(N__38816),
            .in2(N__38801),
            .in3(N__38780),
            .lcout(sbuttonModeStatus_0_sqmuxa_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam spi_data_miso_0_LC_17_16_2.C_ON=1'b0;
    defparam spi_data_miso_0_LC_17_16_2.SEQ_MODE=4'b1010;
    defparam spi_data_miso_0_LC_17_16_2.LUT_INIT=16'b1110111011111100;
    LogicCell40 spi_data_miso_0_LC_17_16_2 (
            .in0(N__38756),
            .in1(N__48902),
            .in2(N__38738),
            .in3(N__43768),
            .lcout(spi_data_misoZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52249),
            .ce(N__43686),
            .sr(N__51680));
    defparam spi_data_miso_4_LC_17_16_6.C_ON=1'b0;
    defparam spi_data_miso_4_LC_17_16_6.SEQ_MODE=4'b1011;
    defparam spi_data_miso_4_LC_17_16_6.LUT_INIT=16'b0011000000100010;
    LogicCell40 spi_data_miso_4_LC_17_16_6 (
            .in0(N__38714),
            .in1(N__48903),
            .in2(N__38693),
            .in3(N__43769),
            .lcout(spi_data_misoZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52249),
            .ce(N__43686),
            .sr(N__51680));
    defparam reset_rpi_ibuf_RNI8S8K1_LC_17_17_0.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNI8S8K1_LC_17_17_0.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNI8S8K1_LC_17_17_0.LUT_INIT=16'b0100000011100000;
    LogicCell40 reset_rpi_ibuf_RNI8S8K1_LC_17_17_0 (
            .in0(N__48899),
            .in1(N__39129),
            .in2(N__49433),
            .in3(N__49479),
            .lcout(N_67_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_23_c_RNITTS3_LC_17_17_1.C_ON=1'b0;
    defparam un4_sacqtime_cry_23_c_RNITTS3_LC_17_17_1.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_23_c_RNITTS3_LC_17_17_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 un4_sacqtime_cry_23_c_RNITTS3_LC_17_17_1 (
            .in0(_gnd_net_),
            .in1(N__43445),
            .in2(_gnd_net_),
            .in3(N__43334),
            .lcout(un4_sacqtime_cry_23_c_RNITTSZ0Z3),
            .ltout(un4_sacqtime_cry_23_c_RNITTSZ0Z3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sSPI_MSB0LSB1_RNILL2C1_LC_17_17_2.C_ON=1'b0;
    defparam sSPI_MSB0LSB1_RNILL2C1_LC_17_17_2.SEQ_MODE=4'b0000;
    defparam sSPI_MSB0LSB1_RNILL2C1_LC_17_17_2.LUT_INIT=16'b1100111011001100;
    LogicCell40 sSPI_MSB0LSB1_RNILL2C1_LC_17_17_2 (
            .in0(N__39165),
            .in1(N__39248),
            .in2(N__39194),
            .in3(N__39127),
            .lcout(N_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sSPI_MSB0LSB1_RNIOT3R1_LC_17_17_3.C_ON=1'b0;
    defparam sSPI_MSB0LSB1_RNIOT3R1_LC_17_17_3.SEQ_MODE=4'b0000;
    defparam sSPI_MSB0LSB1_RNIOT3R1_LC_17_17_3.LUT_INIT=16'b0011001100001010;
    LogicCell40 sSPI_MSB0LSB1_RNIOT3R1_LC_17_17_3 (
            .in0(N__39128),
            .in1(N__49484),
            .in2(N__39173),
            .in3(N__48897),
            .lcout(N_70_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sSPI_MSB0LSB1_RNIGRPG4_LC_17_17_4.C_ON=1'b0;
    defparam sSPI_MSB0LSB1_RNIGRPG4_LC_17_17_4.SEQ_MODE=4'b0000;
    defparam sSPI_MSB0LSB1_RNIGRPG4_LC_17_17_4.LUT_INIT=16'b1111101110111011;
    LogicCell40 sSPI_MSB0LSB1_RNIGRPG4_LC_17_17_4 (
            .in0(N__48898),
            .in1(N__43736),
            .in2(N__39172),
            .in3(N__39130),
            .lcout(sSPI_MSB0LSB1_RNIGRPGZ0Z4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_11_15_LC_17_17_6.C_ON=1'b0;
    defparam RAM_DATA_cl_11_15_LC_17_17_6.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_11_15_LC_17_17_6.LUT_INIT=16'b1000000010100000;
    LogicCell40 RAM_DATA_cl_11_15_LC_17_17_6 (
            .in0(N__48900),
            .in1(N__39082),
            .in2(N__49432),
            .in3(N__49483),
            .lcout(RAM_DATA_cl_11Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52259),
            .ce(),
            .sr(N__51672));
    defparam RAM_DATA_cl_12_15_LC_17_17_7.C_ON=1'b0;
    defparam RAM_DATA_cl_12_15_LC_17_17_7.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_12_15_LC_17_17_7.LUT_INIT=16'b1000110000000000;
    LogicCell40 RAM_DATA_cl_12_15_LC_17_17_7 (
            .in0(N__39058),
            .in1(N__49386),
            .in2(N__49495),
            .in3(N__48901),
            .lcout(RAM_DATA_cl_12Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52259),
            .ce(),
            .sr(N__51672));
    defparam sCounterRAM_0_LC_17_18_0.C_ON=1'b1;
    defparam sCounterRAM_0_LC_17_18_0.SEQ_MODE=4'b1010;
    defparam sCounterRAM_0_LC_17_18_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_0_LC_17_18_0 (
            .in0(N__39509),
            .in1(N__39046),
            .in2(_gnd_net_),
            .in3(N__39032),
            .lcout(sCounterRAMZ0Z_0),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(sCounterRAM_cry_0),
            .clk(N__52271),
            .ce(),
            .sr(N__51664));
    defparam sCounterRAM_1_LC_17_18_1.C_ON=1'b1;
    defparam sCounterRAM_1_LC_17_18_1.SEQ_MODE=4'b1010;
    defparam sCounterRAM_1_LC_17_18_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_1_LC_17_18_1 (
            .in0(N__39505),
            .in1(N__39025),
            .in2(_gnd_net_),
            .in3(N__39011),
            .lcout(sCounterRAMZ0Z_1),
            .ltout(),
            .carryin(sCounterRAM_cry_0),
            .carryout(sCounterRAM_cry_1),
            .clk(N__52271),
            .ce(),
            .sr(N__51664));
    defparam sCounterRAM_2_LC_17_18_2.C_ON=1'b1;
    defparam sCounterRAM_2_LC_17_18_2.SEQ_MODE=4'b1010;
    defparam sCounterRAM_2_LC_17_18_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_2_LC_17_18_2 (
            .in0(N__39510),
            .in1(N__39601),
            .in2(_gnd_net_),
            .in3(N__39587),
            .lcout(sCounterRAMZ0Z_2),
            .ltout(),
            .carryin(sCounterRAM_cry_1),
            .carryout(sCounterRAM_cry_2),
            .clk(N__52271),
            .ce(),
            .sr(N__51664));
    defparam sCounterRAM_3_LC_17_18_3.C_ON=1'b1;
    defparam sCounterRAM_3_LC_17_18_3.SEQ_MODE=4'b1010;
    defparam sCounterRAM_3_LC_17_18_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_3_LC_17_18_3 (
            .in0(N__39506),
            .in1(N__39583),
            .in2(_gnd_net_),
            .in3(N__39569),
            .lcout(sCounterRAMZ0Z_3),
            .ltout(),
            .carryin(sCounterRAM_cry_2),
            .carryout(sCounterRAM_cry_3),
            .clk(N__52271),
            .ce(),
            .sr(N__51664));
    defparam sCounterRAM_4_LC_17_18_4.C_ON=1'b1;
    defparam sCounterRAM_4_LC_17_18_4.SEQ_MODE=4'b1010;
    defparam sCounterRAM_4_LC_17_18_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_4_LC_17_18_4 (
            .in0(N__39511),
            .in1(N__39565),
            .in2(_gnd_net_),
            .in3(N__39551),
            .lcout(sCounterRAMZ0Z_4),
            .ltout(),
            .carryin(sCounterRAM_cry_3),
            .carryout(sCounterRAM_cry_4),
            .clk(N__52271),
            .ce(),
            .sr(N__51664));
    defparam sCounterRAM_5_LC_17_18_5.C_ON=1'b1;
    defparam sCounterRAM_5_LC_17_18_5.SEQ_MODE=4'b1010;
    defparam sCounterRAM_5_LC_17_18_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_5_LC_17_18_5 (
            .in0(N__39507),
            .in1(N__39547),
            .in2(_gnd_net_),
            .in3(N__39533),
            .lcout(sCounterRAMZ0Z_5),
            .ltout(),
            .carryin(sCounterRAM_cry_4),
            .carryout(sCounterRAM_cry_5),
            .clk(N__52271),
            .ce(),
            .sr(N__51664));
    defparam sCounterRAM_6_LC_17_18_6.C_ON=1'b1;
    defparam sCounterRAM_6_LC_17_18_6.SEQ_MODE=4'b1010;
    defparam sCounterRAM_6_LC_17_18_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_6_LC_17_18_6 (
            .in0(N__39512),
            .in1(N__39529),
            .in2(_gnd_net_),
            .in3(N__39515),
            .lcout(sCounterRAMZ0Z_6),
            .ltout(),
            .carryin(sCounterRAM_cry_5),
            .carryout(sCounterRAM_cry_6),
            .clk(N__52271),
            .ce(),
            .sr(N__51664));
    defparam sCounterRAM_7_LC_17_18_7.C_ON=1'b0;
    defparam sCounterRAM_7_LC_17_18_7.SEQ_MODE=4'b1010;
    defparam sCounterRAM_7_LC_17_18_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_7_LC_17_18_7 (
            .in0(N__39508),
            .in1(N__39475),
            .in2(_gnd_net_),
            .in3(N__39482),
            .lcout(sCounterRAMZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52271),
            .ce(),
            .sr(N__51664));
    defparam RAM_DATA_cl_6_15_LC_17_19_0.C_ON=1'b0;
    defparam RAM_DATA_cl_6_15_LC_17_19_0.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_6_15_LC_17_19_0.LUT_INIT=16'b1000000010001000;
    LogicCell40 RAM_DATA_cl_6_15_LC_17_19_0 (
            .in0(N__48948),
            .in1(N__49413),
            .in2(N__39445),
            .in3(N__49536),
            .lcout(RAM_DATA_cl_6Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52280),
            .ce(),
            .sr(N__51659));
    defparam RAM_DATA_cl_7_15_LC_17_19_1.C_ON=1'b0;
    defparam RAM_DATA_cl_7_15_LC_17_19_1.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_7_15_LC_17_19_1.LUT_INIT=16'b1011000000000000;
    LogicCell40 RAM_DATA_cl_7_15_LC_17_19_1 (
            .in0(N__39421),
            .in1(N__49531),
            .in2(N__49440),
            .in3(N__48949),
            .lcout(RAM_DATA_cl_7Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52280),
            .ce(),
            .sr(N__51659));
    defparam RAM_DATA_cl_8_15_LC_17_19_2.C_ON=1'b0;
    defparam RAM_DATA_cl_8_15_LC_17_19_2.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_8_15_LC_17_19_2.LUT_INIT=16'b1000000010001000;
    LogicCell40 RAM_DATA_cl_8_15_LC_17_19_2 (
            .in0(N__48950),
            .in1(N__49417),
            .in2(N__39772),
            .in3(N__49537),
            .lcout(RAM_DATA_cl_8Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52280),
            .ce(),
            .sr(N__51659));
    defparam RAM_DATA_cl_9_15_LC_17_19_4.C_ON=1'b0;
    defparam RAM_DATA_cl_9_15_LC_17_19_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_9_15_LC_17_19_4.LUT_INIT=16'b1000000010001000;
    LogicCell40 RAM_DATA_cl_9_15_LC_17_19_4 (
            .in0(N__48951),
            .in1(N__49418),
            .in2(N__39742),
            .in3(N__49538),
            .lcout(RAM_DATA_cl_9Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52280),
            .ce(),
            .sr(N__51659));
    defparam RAM_DATA_cl_15_LC_17_19_5.C_ON=1'b0;
    defparam RAM_DATA_cl_15_LC_17_19_5.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_15_LC_17_19_5.LUT_INIT=16'b1011000000000000;
    LogicCell40 RAM_DATA_cl_15_LC_17_19_5 (
            .in0(N__39712),
            .in1(N__49530),
            .in2(N__49439),
            .in3(N__48947),
            .lcout(RAM_DATA_clZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52280),
            .ce(),
            .sr(N__51659));
    defparam RAM_DATA_1_7_LC_17_20_4.C_ON=1'b0;
    defparam RAM_DATA_1_7_LC_17_20_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_7_LC_17_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_7_LC_17_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(RAM_DATA_1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52291),
            .ce(N__51896),
            .sr(N__51653));
    defparam sDAC_mem_41_4_LC_18_4_3.C_ON=1'b0;
    defparam sDAC_mem_41_4_LC_18_4_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_4_LC_18_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_4_LC_18_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45600),
            .lcout(sDAC_mem_41Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52260),
            .ce(N__39806),
            .sr(N__51814));
    defparam sDAC_data_RNO_12_6_LC_18_5_6.C_ON=1'b0;
    defparam sDAC_data_RNO_12_6_LC_18_5_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_6_LC_18_5_6.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_12_6_LC_18_5_6 (
            .in0(N__42550),
            .in1(N__39668),
            .in2(N__42263),
            .in3(N__39656),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_6_LC_18_5_7.C_ON=1'b0;
    defparam sDAC_data_RNO_4_6_LC_18_5_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_6_LC_18_5_7.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_6_LC_18_5_7 (
            .in0(N__42094),
            .in1(N__41132),
            .in2(N__39644),
            .in3(N__44495),
            .lcout(sDAC_data_RNO_4Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_32_5_LC_18_6_0.C_ON=1'b0;
    defparam sDAC_mem_32_5_LC_18_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_5_LC_18_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_5_LC_18_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45101),
            .lcout(sDAC_mem_32Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52238),
            .ce(N__41275),
            .sr(N__51799));
    defparam sDAC_mem_32_7_LC_18_6_1.C_ON=1'b0;
    defparam sDAC_mem_32_7_LC_18_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_7_LC_18_6_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_32_7_LC_18_6_1 (
            .in0(N__50032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_32Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52238),
            .ce(N__41275),
            .sr(N__51799));
    defparam sDAC_mem_41_0_LC_18_7_0.C_ON=1'b0;
    defparam sDAC_mem_41_0_LC_18_7_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_0_LC_18_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_0_LC_18_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46389),
            .lcout(sDAC_mem_41Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52228),
            .ce(N__39802),
            .sr(N__51785));
    defparam sDAC_mem_41_1_LC_18_7_1.C_ON=1'b0;
    defparam sDAC_mem_41_1_LC_18_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_1_LC_18_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_1_LC_18_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51050),
            .lcout(sDAC_mem_41Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52228),
            .ce(N__39802),
            .sr(N__51785));
    defparam sDAC_mem_41_2_LC_18_7_2.C_ON=1'b0;
    defparam sDAC_mem_41_2_LC_18_7_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_2_LC_18_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_2_LC_18_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47481),
            .lcout(sDAC_mem_41Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52228),
            .ce(N__39802),
            .sr(N__51785));
    defparam sDAC_mem_41_3_LC_18_7_3.C_ON=1'b0;
    defparam sDAC_mem_41_3_LC_18_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_3_LC_18_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_3_LC_18_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46921),
            .lcout(sDAC_mem_41Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52228),
            .ce(N__39802),
            .sr(N__51785));
    defparam sDAC_mem_41_5_LC_18_7_5.C_ON=1'b0;
    defparam sDAC_mem_41_5_LC_18_7_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_5_LC_18_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_5_LC_18_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45102),
            .lcout(sDAC_mem_41Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52228),
            .ce(N__39802),
            .sr(N__51785));
    defparam sDAC_mem_41_6_LC_18_7_6.C_ON=1'b0;
    defparam sDAC_mem_41_6_LC_18_7_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_6_LC_18_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_6_LC_18_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50379),
            .lcout(sDAC_mem_41Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52228),
            .ce(N__39802),
            .sr(N__51785));
    defparam sDAC_mem_41_7_LC_18_7_7.C_ON=1'b0;
    defparam sDAC_mem_41_7_LC_18_7_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_7_LC_18_7_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_41_7_LC_18_7_7 (
            .in0(N__50034),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_41Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52228),
            .ce(N__39802),
            .sr(N__51785));
    defparam sAddress_RNI9IH12_9_5_LC_18_8_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_9_5_LC_18_8_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_9_5_LC_18_8_0.LUT_INIT=16'b0000100000000000;
    LogicCell40 sAddress_RNI9IH12_9_5_LC_18_8_0 (
            .in0(N__40799),
            .in1(N__41026),
            .in2(N__41000),
            .in3(N__40418),
            .lcout(sDAC_mem_9_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_1_5_LC_18_8_1.C_ON=1'b0;
    defparam sAddress_RNI9IH12_1_5_LC_18_8_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_1_5_LC_18_8_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 sAddress_RNI9IH12_1_5_LC_18_8_1 (
            .in0(N__40417),
            .in1(N__40978),
            .in2(N__41027),
            .in3(N__40797),
            .lcout(sDAC_mem_41_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI6VH7_6_1_LC_18_8_2.C_ON=1'b0;
    defparam sAddress_RNI6VH7_6_1_LC_18_8_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI6VH7_6_1_LC_18_8_2.LUT_INIT=16'b0000000000010001;
    LogicCell40 sAddress_RNI6VH7_6_1_LC_18_8_2 (
            .in0(N__40652),
            .in1(N__40546),
            .in2(_gnd_net_),
            .in3(N__40197),
            .lcout(sAddress_RNI6VH7_6Z0Z_1),
            .ltout(sAddress_RNI6VH7_6Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_1_3_LC_18_8_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_1_3_LC_18_8_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_1_3_LC_18_8_3.LUT_INIT=16'b1100000000000000;
    LogicCell40 sAddress_RNI9IH12_1_3_LC_18_8_3 (
            .in0(_gnd_net_),
            .in1(N__40416),
            .in2(N__41015),
            .in3(N__40027),
            .lcout(sDAC_mem_25_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_4_5_LC_18_8_4.C_ON=1'b0;
    defparam sAddress_RNI9IH12_4_5_LC_18_8_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_4_5_LC_18_8_4.LUT_INIT=16'b0000101000000000;
    LogicCell40 sAddress_RNI9IH12_4_5_LC_18_8_4 (
            .in0(N__40798),
            .in1(_gnd_net_),
            .in2(N__40999),
            .in3(N__40053),
            .lcout(sDAC_mem_1_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_0_5_LC_18_8_5.C_ON=1'b0;
    defparam sAddress_RNI9IH12_0_5_LC_18_8_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_0_5_LC_18_8_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 sAddress_RNI9IH12_0_5_LC_18_8_5 (
            .in0(N__40052),
            .in1(N__40985),
            .in2(_gnd_net_),
            .in3(N__40800),
            .lcout(sDAC_mem_33_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIAM2A_1_1_LC_18_8_6.C_ON=1'b0;
    defparam sAddress_RNIAM2A_1_1_LC_18_8_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNIAM2A_1_1_LC_18_8_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 sAddress_RNIAM2A_1_1_LC_18_8_6 (
            .in0(N__40651),
            .in1(N__40547),
            .in2(N__40429),
            .in3(N__40196),
            .lcout(sAddress_RNIAM2A_1Z0Z_1),
            .ltout(sAddress_RNIAM2A_1Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_0_1_LC_18_8_7.C_ON=1'b0;
    defparam sAddress_RNI9IH12_0_1_LC_18_8_7.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_0_1_LC_18_8_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 sAddress_RNI9IH12_0_1_LC_18_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40031),
            .in3(N__40026),
            .lcout(sDAC_mem_17_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_37_0_LC_18_9_0.C_ON=1'b0;
    defparam sDAC_mem_37_0_LC_18_9_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_0_LC_18_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_0_LC_18_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46374),
            .lcout(sDAC_mem_37Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52214),
            .ce(N__41075),
            .sr(N__51760));
    defparam sDAC_mem_37_1_LC_18_9_1.C_ON=1'b0;
    defparam sDAC_mem_37_1_LC_18_9_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_1_LC_18_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_1_LC_18_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51042),
            .lcout(sDAC_mem_37Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52214),
            .ce(N__41075),
            .sr(N__51760));
    defparam sDAC_mem_37_2_LC_18_9_2.C_ON=1'b0;
    defparam sDAC_mem_37_2_LC_18_9_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_2_LC_18_9_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_37_2_LC_18_9_2 (
            .in0(N__47484),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_37Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52214),
            .ce(N__41075),
            .sr(N__51760));
    defparam sDAC_mem_37_3_LC_18_9_3.C_ON=1'b0;
    defparam sDAC_mem_37_3_LC_18_9_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_3_LC_18_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_3_LC_18_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46855),
            .lcout(sDAC_mem_37Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52214),
            .ce(N__41075),
            .sr(N__51760));
    defparam sDAC_mem_37_4_LC_18_9_4.C_ON=1'b0;
    defparam sDAC_mem_37_4_LC_18_9_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_4_LC_18_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_4_LC_18_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45593),
            .lcout(sDAC_mem_37Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52214),
            .ce(N__41075),
            .sr(N__51760));
    defparam sDAC_mem_37_5_LC_18_9_5.C_ON=1'b0;
    defparam sDAC_mem_37_5_LC_18_9_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_5_LC_18_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_5_LC_18_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45106),
            .lcout(sDAC_mem_37Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52214),
            .ce(N__41075),
            .sr(N__51760));
    defparam sDAC_mem_37_6_LC_18_9_6.C_ON=1'b0;
    defparam sDAC_mem_37_6_LC_18_9_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_6_LC_18_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_6_LC_18_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50380),
            .lcout(sDAC_mem_37Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52214),
            .ce(N__41075),
            .sr(N__51760));
    defparam sDAC_mem_37_7_LC_18_9_7.C_ON=1'b0;
    defparam sDAC_mem_37_7_LC_18_9_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_7_LC_18_9_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_37_7_LC_18_9_7 (
            .in0(N__50037),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_37Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52214),
            .ce(N__41075),
            .sr(N__51760));
    defparam sDAC_data_RNO_14_3_LC_18_10_0.C_ON=1'b0;
    defparam sDAC_data_RNO_14_3_LC_18_10_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_3_LC_18_10_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_14_3_LC_18_10_0 (
            .in0(N__42188),
            .in1(N__41033),
            .in2(_gnd_net_),
            .in3(N__41060),
            .lcout(sDAC_data_RNO_14Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_26_4_LC_18_10_1.C_ON=1'b0;
    defparam sDAC_data_RNO_26_4_LC_18_10_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_4_LC_18_10_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_26_4_LC_18_10_1 (
            .in0(N__42526),
            .in1(N__44378),
            .in2(_gnd_net_),
            .in3(N__44123),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_4_LC_18_10_2.C_ON=1'b0;
    defparam sDAC_data_RNO_14_4_LC_18_10_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_4_LC_18_10_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 sDAC_data_RNO_14_4_LC_18_10_2 (
            .in0(_gnd_net_),
            .in1(N__42001),
            .in2(N__41048),
            .in3(N__41297),
            .lcout(sDAC_data_RNO_14Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_32_0_LC_18_10_3.C_ON=1'b0;
    defparam sDAC_mem_32_0_LC_18_10_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_0_LC_18_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_0_LC_18_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46344),
            .lcout(sDAC_mem_32Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52208),
            .ce(N__41276),
            .sr(N__51748));
    defparam sDAC_mem_32_1_LC_18_10_4.C_ON=1'b0;
    defparam sDAC_mem_32_1_LC_18_10_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_1_LC_18_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_1_LC_18_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51063),
            .lcout(sDAC_mem_32Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52208),
            .ce(N__41276),
            .sr(N__51748));
    defparam sDAC_data_RNO_26_5_LC_18_10_5.C_ON=1'b0;
    defparam sDAC_data_RNO_26_5_LC_18_10_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_5_LC_18_10_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_26_5_LC_18_10_5 (
            .in0(N__42527),
            .in1(N__44369),
            .in2(_gnd_net_),
            .in3(N__44111),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_5_LC_18_10_6.C_ON=1'b0;
    defparam sDAC_data_RNO_14_5_LC_18_10_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_5_LC_18_10_6.LUT_INIT=16'b1111001111000000;
    LogicCell40 sDAC_data_RNO_14_5_LC_18_10_6 (
            .in0(_gnd_net_),
            .in1(N__42002),
            .in2(N__41291),
            .in3(N__41282),
            .lcout(sDAC_data_RNO_14Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_32_2_LC_18_10_7.C_ON=1'b0;
    defparam sDAC_mem_32_2_LC_18_10_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_2_LC_18_10_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_32_2_LC_18_10_7 (
            .in0(N__47497),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_32Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52208),
            .ce(N__41276),
            .sr(N__51748));
    defparam sDAC_data_RNO_12_3_LC_18_11_0.C_ON=1'b0;
    defparam sDAC_data_RNO_12_3_LC_18_11_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_3_LC_18_11_0.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_12_3_LC_18_11_0 (
            .in0(N__42528),
            .in1(N__41213),
            .in2(N__42244),
            .in3(N__41177),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_3_LC_18_11_1.C_ON=1'b0;
    defparam sDAC_data_RNO_4_3_LC_18_11_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_3_LC_18_11_1.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_3_LC_18_11_1 (
            .in0(N__42033),
            .in1(N__41201),
            .in2(N__41192),
            .in3(N__44522),
            .lcout(sDAC_data_RNO_4Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_4_0_LC_18_11_2.C_ON=1'b0;
    defparam sDAC_mem_4_0_LC_18_11_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_0_LC_18_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_0_LC_18_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46384),
            .lcout(sDAC_mem_4Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52205),
            .ce(N__42641),
            .sr(N__51733));
    defparam sDAC_data_RNO_12_4_LC_18_11_3.C_ON=1'b0;
    defparam sDAC_data_RNO_12_4_LC_18_11_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_4_LC_18_11_3.LUT_INIT=16'b0101010100100111;
    LogicCell40 sDAC_data_RNO_12_4_LC_18_11_3 (
            .in0(N__42566),
            .in1(N__41171),
            .in2(N__42650),
            .in3(N__42181),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_4_LC_18_11_4.C_ON=1'b0;
    defparam sDAC_data_RNO_4_4_LC_18_11_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_4_LC_18_11_4.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_4_4_LC_18_11_4 (
            .in0(N__44513),
            .in1(N__42032),
            .in2(N__41156),
            .in3(N__41153),
            .lcout(sDAC_data_RNO_4Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_4_1_LC_18_11_5.C_ON=1'b0;
    defparam sDAC_mem_4_1_LC_18_11_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_1_LC_18_11_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_4_1_LC_18_11_5 (
            .in0(N__51077),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_4Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52205),
            .ce(N__42641),
            .sr(N__51733));
    defparam sDAC_data_RNO_12_5_LC_18_11_6.C_ON=1'b0;
    defparam sDAC_data_RNO_12_5_LC_18_11_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_5_LC_18_11_6.LUT_INIT=16'b0101001001010111;
    LogicCell40 sDAC_data_RNO_12_5_LC_18_11_6 (
            .in0(N__42529),
            .in1(N__42293),
            .in2(N__42245),
            .in3(N__42278),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_5_LC_18_11_7.C_ON=1'b0;
    defparam sDAC_data_RNO_4_5_LC_18_11_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_5_LC_18_11_7.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_5_LC_18_11_7 (
            .in0(N__42034),
            .in1(N__41387),
            .in2(N__41378),
            .in3(N__44504),
            .lcout(sDAC_data_RNO_4Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_25_5_LC_18_12_1.C_ON=1'b0;
    defparam sDAC_mem_25_5_LC_18_12_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_5_LC_18_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_5_LC_18_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45115),
            .lcout(sDAC_mem_25Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52209),
            .ce(N__50593),
            .sr(N__51721));
    defparam sDAC_mem_25_2_LC_18_12_2.C_ON=1'b0;
    defparam sDAC_mem_25_2_LC_18_12_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_2_LC_18_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_2_LC_18_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47507),
            .lcout(sDAC_mem_25Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52209),
            .ce(N__50593),
            .sr(N__51721));
    defparam sDAC_mem_25_3_LC_18_12_3.C_ON=1'b0;
    defparam sDAC_mem_25_3_LC_18_12_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_3_LC_18_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_3_LC_18_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46923),
            .lcout(sDAC_mem_25Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52209),
            .ce(N__50593),
            .sr(N__51721));
    defparam sDAC_mem_25_4_LC_18_12_4.C_ON=1'b0;
    defparam sDAC_mem_25_4_LC_18_12_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_4_LC_18_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_4_LC_18_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45607),
            .lcout(sDAC_mem_25Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52209),
            .ce(N__50593),
            .sr(N__51721));
    defparam sDAC_mem_25_0_LC_18_12_5.C_ON=1'b0;
    defparam sDAC_mem_25_0_LC_18_12_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_0_LC_18_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_0_LC_18_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46317),
            .lcout(sDAC_mem_25Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52209),
            .ce(N__50593),
            .sr(N__51721));
    defparam sDAC_mem_25_6_LC_18_12_6.C_ON=1'b0;
    defparam sDAC_mem_25_6_LC_18_12_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_6_LC_18_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_6_LC_18_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50381),
            .lcout(sDAC_mem_25Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52209),
            .ce(N__50593),
            .sr(N__51721));
    defparam sDAC_mem_25_7_LC_18_12_7.C_ON=1'b0;
    defparam sDAC_mem_25_7_LC_18_12_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_7_LC_18_12_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_25_7_LC_18_12_7 (
            .in0(N__50063),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_25Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52209),
            .ce(N__50593),
            .sr(N__51721));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_0_LC_18_13_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_0_LC_18_13_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_0_LC_18_13_0 .LUT_INIT=16'b0000101110110000;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_0_LC_18_13_0  (
            .in0(N__51213),
            .in1(N__42706),
            .in2(N__42791),
            .in3(N__42768),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48264),
            .ce(),
            .sr(N__51710));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_1_LC_18_13_1 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_1_LC_18_13_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_1_LC_18_13_1 .LUT_INIT=16'b0011110000010100;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_1_LC_18_13_1  (
            .in0(N__42705),
            .in1(N__42746),
            .in2(N__42736),
            .in3(N__51214),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48264),
            .ce(),
            .sr(N__51710));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_2_LC_18_13_2 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_2_LC_18_13_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_2_LC_18_13_2 .LUT_INIT=16'b0010001110001100;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_2_LC_18_13_2  (
            .in0(N__51215),
            .in1(N__42679),
            .in2(N__42710),
            .in3(N__42689),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48264),
            .ce(),
            .sr(N__51710));
    defparam \spi_slave_inst.txdata_reg_i_RNI3KQC_1_LC_18_13_3 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_RNI3KQC_1_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.txdata_reg_i_RNI3KQC_1_LC_18_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi_slave_inst.txdata_reg_i_RNI3KQC_1_LC_18_13_3  (
            .in0(N__47519),
            .in1(N__45782),
            .in2(_gnd_net_),
            .in3(N__48729),
            .lcout(\spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.txdata_reg_i_RNI5MQC_2_LC_18_13_4 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_RNI5MQC_2_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.txdata_reg_i_RNI5MQC_2_LC_18_13_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi_slave_inst.txdata_reg_i_RNI5MQC_2_LC_18_13_4  (
            .in0(N__48730),
            .in1(N__45674),
            .in2(_gnd_net_),
            .in3(N__45797),
            .lcout(\spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.txdata_reg_i_RNI7OQC_3_LC_18_13_5 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_RNI7OQC_3_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.txdata_reg_i_RNI7OQC_3_LC_18_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi_slave_inst.txdata_reg_i_RNI7OQC_3_LC_18_13_5  (
            .in0(N__45686),
            .in1(N__50558),
            .in2(_gnd_net_),
            .in3(N__48731),
            .lcout(\spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.data_in_reg_i_0_LC_18_14_0 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_0_LC_18_14_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_0_LC_18_14_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.data_in_reg_i_0_LC_18_14_0  (
            .in0(N__42659),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52221),
            .ce(N__42830),
            .sr(N__51701));
    defparam \spi_slave_inst.data_in_reg_i_1_LC_18_14_1 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_1_LC_18_14_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_1_LC_18_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_1_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43700),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52221),
            .ce(N__42830),
            .sr(N__51701));
    defparam \spi_slave_inst.data_in_reg_i_2_LC_18_14_2 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_2_LC_18_14_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_2_LC_18_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_2_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42854),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52221),
            .ce(N__42830),
            .sr(N__51701));
    defparam \spi_slave_inst.data_in_reg_i_3_LC_18_14_3 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_3_LC_18_14_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_3_LC_18_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_3_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42896),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52221),
            .ce(N__42830),
            .sr(N__51701));
    defparam \spi_slave_inst.data_in_reg_i_4_LC_18_14_4 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_4_LC_18_14_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_4_LC_18_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_4_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42845),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52221),
            .ce(N__42830),
            .sr(N__51701));
    defparam \spi_slave_inst.data_in_reg_i_5_LC_18_14_5 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_5_LC_18_14_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_5_LC_18_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_5_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42989),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52221),
            .ce(N__42830),
            .sr(N__51701));
    defparam \spi_slave_inst.data_in_reg_i_6_LC_18_14_6 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_6_LC_18_14_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_6_LC_18_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_6_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42836),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52221),
            .ce(N__42830),
            .sr(N__51701));
    defparam \spi_slave_inst.data_in_reg_i_7_LC_18_14_7 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_7_LC_18_14_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_7_LC_18_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_7_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42944),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52221),
            .ce(N__42830),
            .sr(N__51701));
    defparam sCounterADC_0_LC_18_15_0.C_ON=1'b1;
    defparam sCounterADC_0_LC_18_15_0.SEQ_MODE=4'b1010;
    defparam sCounterADC_0_LC_18_15_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_0_LC_18_15_0 (
            .in0(N__46960),
            .in1(N__46409),
            .in2(_gnd_net_),
            .in3(N__42812),
            .lcout(sCounterADCZ0Z_0),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(sCounterADC_cry_0),
            .clk(N__52229),
            .ce(N__48960),
            .sr(N__51692));
    defparam sCounterADC_1_LC_18_15_1.C_ON=1'b1;
    defparam sCounterADC_1_LC_18_15_1.SEQ_MODE=4'b1010;
    defparam sCounterADC_1_LC_18_15_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_1_LC_18_15_1 (
            .in0(N__46956),
            .in1(N__46421),
            .in2(_gnd_net_),
            .in3(N__42809),
            .lcout(sCounterADCZ0Z_1),
            .ltout(),
            .carryin(sCounterADC_cry_0),
            .carryout(sCounterADC_cry_1),
            .clk(N__52229),
            .ce(N__48960),
            .sr(N__51692));
    defparam sCounterADC_2_LC_18_15_2.C_ON=1'b1;
    defparam sCounterADC_2_LC_18_15_2.SEQ_MODE=4'b1010;
    defparam sCounterADC_2_LC_18_15_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_2_LC_18_15_2 (
            .in0(N__46961),
            .in1(N__47018),
            .in2(_gnd_net_),
            .in3(N__42806),
            .lcout(sCounterADCZ0Z_2),
            .ltout(),
            .carryin(sCounterADC_cry_1),
            .carryout(sCounterADC_cry_2),
            .clk(N__52229),
            .ce(N__48960),
            .sr(N__51692));
    defparam sCounterADC_3_LC_18_15_3.C_ON=1'b1;
    defparam sCounterADC_3_LC_18_15_3.SEQ_MODE=4'b1010;
    defparam sCounterADC_3_LC_18_15_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_3_LC_18_15_3 (
            .in0(N__46957),
            .in1(N__47000),
            .in2(_gnd_net_),
            .in3(N__43082),
            .lcout(sCounterADCZ0Z_3),
            .ltout(),
            .carryin(sCounterADC_cry_2),
            .carryout(sCounterADC_cry_3),
            .clk(N__52229),
            .ce(N__48960),
            .sr(N__51692));
    defparam sCounterADC_4_LC_18_15_4.C_ON=1'b1;
    defparam sCounterADC_4_LC_18_15_4.SEQ_MODE=4'b1010;
    defparam sCounterADC_4_LC_18_15_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_4_LC_18_15_4 (
            .in0(N__46962),
            .in1(N__43069),
            .in2(_gnd_net_),
            .in3(N__43055),
            .lcout(sCounterADCZ0Z_4),
            .ltout(),
            .carryin(sCounterADC_cry_3),
            .carryout(sCounterADC_cry_4),
            .clk(N__52229),
            .ce(N__48960),
            .sr(N__51692));
    defparam sCounterADC_5_LC_18_15_5.C_ON=1'b1;
    defparam sCounterADC_5_LC_18_15_5.SEQ_MODE=4'b1010;
    defparam sCounterADC_5_LC_18_15_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_5_LC_18_15_5 (
            .in0(N__46958),
            .in1(N__43042),
            .in2(_gnd_net_),
            .in3(N__43028),
            .lcout(sCounterADCZ0Z_5),
            .ltout(),
            .carryin(sCounterADC_cry_4),
            .carryout(sCounterADC_cry_5),
            .clk(N__52229),
            .ce(N__48960),
            .sr(N__51692));
    defparam sCounterADC_6_LC_18_15_6.C_ON=1'b1;
    defparam sCounterADC_6_LC_18_15_6.SEQ_MODE=4'b1010;
    defparam sCounterADC_6_LC_18_15_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_6_LC_18_15_6 (
            .in0(N__46963),
            .in1(N__45844),
            .in2(_gnd_net_),
            .in3(N__43025),
            .lcout(sCounterADCZ0Z_6),
            .ltout(),
            .carryin(sCounterADC_cry_5),
            .carryout(sCounterADC_cry_6),
            .clk(N__52229),
            .ce(N__48960),
            .sr(N__51692));
    defparam sCounterADC_7_LC_18_15_7.C_ON=1'b0;
    defparam sCounterADC_7_LC_18_15_7.SEQ_MODE=4'b1010;
    defparam sCounterADC_7_LC_18_15_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_7_LC_18_15_7 (
            .in0(N__46959),
            .in1(N__45857),
            .in2(_gnd_net_),
            .in3(N__43022),
            .lcout(sCounterADCZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52229),
            .ce(N__48960),
            .sr(N__51692));
    defparam spi_data_miso_5_LC_18_16_0.C_ON=1'b0;
    defparam spi_data_miso_5_LC_18_16_0.SEQ_MODE=4'b1011;
    defparam spi_data_miso_5_LC_18_16_0.LUT_INIT=16'b0000000010101100;
    LogicCell40 spi_data_miso_5_LC_18_16_0 (
            .in0(N__43019),
            .in1(N__43001),
            .in2(N__43772),
            .in3(N__48910),
            .lcout(spi_data_misoZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52239),
            .ce(N__43691),
            .sr(N__51686));
    defparam spi_data_miso_7_LC_18_16_1.C_ON=1'b0;
    defparam spi_data_miso_7_LC_18_16_1.SEQ_MODE=4'b1010;
    defparam spi_data_miso_7_LC_18_16_1.LUT_INIT=16'b1111101011101110;
    LogicCell40 spi_data_miso_7_LC_18_16_1 (
            .in0(N__48911),
            .in1(N__42980),
            .in2(N__42968),
            .in3(N__43766),
            .lcout(spi_data_misoZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52239),
            .ce(N__43691),
            .sr(N__51686));
    defparam spi_data_miso_3_LC_18_16_3.C_ON=1'b0;
    defparam spi_data_miso_3_LC_18_16_3.SEQ_MODE=4'b1010;
    defparam spi_data_miso_3_LC_18_16_3.LUT_INIT=16'b0100010001010000;
    LogicCell40 spi_data_miso_3_LC_18_16_3 (
            .in0(N__48909),
            .in1(N__42935),
            .in2(N__42917),
            .in3(N__43765),
            .lcout(spi_data_misoZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52239),
            .ce(N__43691),
            .sr(N__51686));
    defparam spi_data_miso_2_LC_18_16_4.C_ON=1'b0;
    defparam spi_data_miso_2_LC_18_16_4.SEQ_MODE=4'b1011;
    defparam spi_data_miso_2_LC_18_16_4.LUT_INIT=16'b0000000011001010;
    LogicCell40 spi_data_miso_2_LC_18_16_4 (
            .in0(N__42887),
            .in1(N__42872),
            .in2(N__43771),
            .in3(N__48908),
            .lcout(spi_data_misoZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52239),
            .ce(N__43691),
            .sr(N__51686));
    defparam spi_data_miso_1_LC_18_16_6.C_ON=1'b0;
    defparam spi_data_miso_1_LC_18_16_6.SEQ_MODE=4'b1011;
    defparam spi_data_miso_1_LC_18_16_6.LUT_INIT=16'b0000000010101100;
    LogicCell40 spi_data_miso_1_LC_18_16_6 (
            .in0(N__43808),
            .in1(N__43787),
            .in2(N__43770),
            .in3(N__48907),
            .lcout(spi_data_misoZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52239),
            .ce(N__43691),
            .sr(N__51686));
    defparam sRAM_ADD_8_LC_18_17_0.C_ON=1'b0;
    defparam sRAM_ADD_8_LC_18_17_0.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_8_LC_18_17_0.LUT_INIT=16'b1101100011110000;
    LogicCell40 sRAM_ADD_8_LC_18_17_0 (
            .in0(N__43347),
            .in1(N__43661),
            .in2(N__43634),
            .in3(N__43468),
            .lcout(RAM_ADD_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52250),
            .ce(N__43225),
            .sr(_gnd_net_));
    defparam sRAM_ADD_4_LC_18_17_6.C_ON=1'b0;
    defparam sRAM_ADD_4_LC_18_17_6.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_4_LC_18_17_6.LUT_INIT=16'b1101100011110000;
    LogicCell40 sRAM_ADD_4_LC_18_17_6 (
            .in0(N__43346),
            .in1(N__43589),
            .in2(N__43562),
            .in3(N__43467),
            .lcout(RAM_ADD_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52250),
            .ce(N__43225),
            .sr(_gnd_net_));
    defparam sRAM_ADD_3_LC_18_17_7.C_ON=1'b0;
    defparam sRAM_ADD_3_LC_18_17_7.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_3_LC_18_17_7.LUT_INIT=16'b1011100011110000;
    LogicCell40 sRAM_ADD_3_LC_18_17_7 (
            .in0(N__43520),
            .in1(N__43466),
            .in2(N__43376),
            .in3(N__43345),
            .lcout(RAM_ADD_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52250),
            .ce(N__43225),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_13_15_LC_18_18_0.C_ON=1'b0;
    defparam RAM_DATA_cl_13_15_LC_18_18_0.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_13_15_LC_18_18_0.LUT_INIT=16'b1011000000000000;
    LogicCell40 RAM_DATA_cl_13_15_LC_18_18_0 (
            .in0(N__43183),
            .in1(N__49527),
            .in2(N__49436),
            .in3(N__48930),
            .lcout(RAM_DATA_cl_13Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52261),
            .ce(),
            .sr(N__51673));
    defparam RAM_DATA_cl_14_15_LC_18_18_1.C_ON=1'b0;
    defparam RAM_DATA_cl_14_15_LC_18_18_1.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_14_15_LC_18_18_1.LUT_INIT=16'b1000000010001000;
    LogicCell40 RAM_DATA_cl_14_15_LC_18_18_1 (
            .in0(N__48931),
            .in1(N__49400),
            .in2(N__43159),
            .in3(N__49532),
            .lcout(RAM_DATA_cl_14Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52261),
            .ce(),
            .sr(N__51673));
    defparam RAM_DATA_cl_15_15_LC_18_18_2.C_ON=1'b0;
    defparam RAM_DATA_cl_15_15_LC_18_18_2.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_15_15_LC_18_18_2.LUT_INIT=16'b1011000000000000;
    LogicCell40 RAM_DATA_cl_15_15_LC_18_18_2 (
            .in0(N__43126),
            .in1(N__49528),
            .in2(N__49437),
            .in3(N__48932),
            .lcout(RAM_DATA_cl_15Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52261),
            .ce(),
            .sr(N__51673));
    defparam RAM_DATA_cl_1_15_LC_18_18_3.C_ON=1'b0;
    defparam RAM_DATA_cl_1_15_LC_18_18_3.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_1_15_LC_18_18_3.LUT_INIT=16'b1000000010001000;
    LogicCell40 RAM_DATA_cl_1_15_LC_18_18_3 (
            .in0(N__48933),
            .in1(N__49404),
            .in2(N__43099),
            .in3(N__49533),
            .lcout(RAM_DATA_cl_1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52261),
            .ce(),
            .sr(N__51673));
    defparam RAM_DATA_cl_10_15_LC_18_18_4.C_ON=1'b0;
    defparam RAM_DATA_cl_10_15_LC_18_18_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_10_15_LC_18_18_4.LUT_INIT=16'b1011000000000000;
    LogicCell40 RAM_DATA_cl_10_15_LC_18_18_4 (
            .in0(N__44056),
            .in1(N__49526),
            .in2(N__49435),
            .in3(N__48929),
            .lcout(RAM_DATA_cl_10Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52261),
            .ce(),
            .sr(N__51673));
    defparam RAM_DATA_cl_3_15_LC_18_18_5.C_ON=1'b0;
    defparam RAM_DATA_cl_3_15_LC_18_18_5.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_3_15_LC_18_18_5.LUT_INIT=16'b1000000010001000;
    LogicCell40 RAM_DATA_cl_3_15_LC_18_18_5 (
            .in0(N__48935),
            .in1(N__49406),
            .in2(N__44032),
            .in3(N__49535),
            .lcout(RAM_DATA_cl_3Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52261),
            .ce(),
            .sr(N__51673));
    defparam RAM_DATA_cl_4_15_LC_18_18_6.C_ON=1'b0;
    defparam RAM_DATA_cl_4_15_LC_18_18_6.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_4_15_LC_18_18_6.LUT_INIT=16'b1011000000000000;
    LogicCell40 RAM_DATA_cl_4_15_LC_18_18_6 (
            .in0(N__43999),
            .in1(N__49529),
            .in2(N__49438),
            .in3(N__48936),
            .lcout(RAM_DATA_cl_4Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52261),
            .ce(),
            .sr(N__51673));
    defparam RAM_DATA_cl_2_15_LC_18_18_7.C_ON=1'b0;
    defparam RAM_DATA_cl_2_15_LC_18_18_7.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_2_15_LC_18_18_7.LUT_INIT=16'b1000000010001000;
    LogicCell40 RAM_DATA_cl_2_15_LC_18_18_7 (
            .in0(N__48934),
            .in1(N__49405),
            .in2(N__43975),
            .in3(N__49534),
            .lcout(RAM_DATA_cl_2Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52261),
            .ce(),
            .sr(N__51673));
    defparam sDAC_data_2_LC_19_1_1.C_ON=1'b0;
    defparam sDAC_data_2_LC_19_1_1.SEQ_MODE=4'b1010;
    defparam sDAC_data_2_LC_19_1_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_2_LC_19_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48454),
            .ce(N__43955),
            .sr(N__51826));
    defparam \spi_master_inst.spi_data_path_u1.data_in_2_LC_19_3_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_2_LC_19_3_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_2_LC_19_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_2_LC_19_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43916),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48458),
            .ce(N__43907),
            .sr(N__51824));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_2_LC_19_4_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_2_LC_19_4_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_2_LC_19_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_2_LC_19_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43853),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48460),
            .ce(),
            .sr(N__51820));
    defparam sDAC_mem_7_2_LC_19_5_0.C_ON=1'b0;
    defparam sDAC_mem_7_2_LC_19_5_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_2_LC_19_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_7_2_LC_19_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47329),
            .lcout(sDAC_mem_7Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52240),
            .ce(N__44285),
            .sr(N__51815));
    defparam sDAC_mem_7_3_LC_19_5_1.C_ON=1'b0;
    defparam sDAC_mem_7_3_LC_19_5_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_3_LC_19_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_7_3_LC_19_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46789),
            .lcout(sDAC_mem_7Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52240),
            .ce(N__44285),
            .sr(N__51815));
    defparam sDAC_mem_7_4_LC_19_5_2.C_ON=1'b0;
    defparam sDAC_mem_7_4_LC_19_5_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_4_LC_19_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_7_4_LC_19_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45359),
            .lcout(sDAC_mem_7Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52240),
            .ce(N__44285),
            .sr(N__51815));
    defparam sDAC_mem_7_6_LC_19_5_3.C_ON=1'b0;
    defparam sDAC_mem_7_6_LC_19_5_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_6_LC_19_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_7_6_LC_19_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50374),
            .lcout(sDAC_mem_7Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52240),
            .ce(N__44285),
            .sr(N__51815));
    defparam sDAC_mem_3_7_LC_19_6_0.C_ON=1'b0;
    defparam sDAC_mem_3_7_LC_19_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_7_LC_19_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_3_7_LC_19_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50033),
            .lcout(sDAC_mem_3Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52230),
            .ce(N__44239),
            .sr(N__51808));
    defparam sDAC_mem_1_0_LC_19_7_0.C_ON=1'b0;
    defparam sDAC_mem_1_0_LC_19_7_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_0_LC_19_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_0_LC_19_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46390),
            .lcout(sDAC_mem_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52222),
            .ce(N__44402),
            .sr(N__51800));
    defparam sDAC_mem_1_1_LC_19_7_1.C_ON=1'b0;
    defparam sDAC_mem_1_1_LC_19_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_1_LC_19_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_1_LC_19_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51051),
            .lcout(sDAC_mem_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52222),
            .ce(N__44402),
            .sr(N__51800));
    defparam sDAC_mem_1_2_LC_19_7_2.C_ON=1'b0;
    defparam sDAC_mem_1_2_LC_19_7_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_2_LC_19_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_2_LC_19_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47482),
            .lcout(sDAC_mem_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52222),
            .ce(N__44402),
            .sr(N__51800));
    defparam sDAC_mem_1_3_LC_19_7_3.C_ON=1'b0;
    defparam sDAC_mem_1_3_LC_19_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_3_LC_19_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_3_LC_19_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46922),
            .lcout(sDAC_mem_1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52222),
            .ce(N__44402),
            .sr(N__51800));
    defparam sDAC_mem_1_4_LC_19_7_4.C_ON=1'b0;
    defparam sDAC_mem_1_4_LC_19_7_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_4_LC_19_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_4_LC_19_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45561),
            .lcout(sDAC_mem_1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52222),
            .ce(N__44402),
            .sr(N__51800));
    defparam sDAC_mem_1_5_LC_19_7_5.C_ON=1'b0;
    defparam sDAC_mem_1_5_LC_19_7_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_5_LC_19_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_5_LC_19_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45064),
            .lcout(sDAC_mem_1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52222),
            .ce(N__44402),
            .sr(N__51800));
    defparam sDAC_mem_1_6_LC_19_7_6.C_ON=1'b0;
    defparam sDAC_mem_1_6_LC_19_7_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_6_LC_19_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_6_LC_19_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50464),
            .lcout(sDAC_mem_1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52222),
            .ce(N__44402),
            .sr(N__51800));
    defparam sDAC_mem_1_7_LC_19_7_7.C_ON=1'b0;
    defparam sDAC_mem_1_7_LC_19_7_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_7_LC_19_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_7_LC_19_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50035),
            .lcout(sDAC_mem_1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52222),
            .ce(N__44402),
            .sr(N__51800));
    defparam sDAC_mem_33_0_LC_19_8_0.C_ON=1'b0;
    defparam sDAC_mem_33_0_LC_19_8_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_0_LC_19_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_0_LC_19_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46382),
            .lcout(sDAC_mem_33Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52215),
            .ce(N__44531),
            .sr(N__51786));
    defparam sDAC_mem_33_1_LC_19_8_1.C_ON=1'b0;
    defparam sDAC_mem_33_1_LC_19_8_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_1_LC_19_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_1_LC_19_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51076),
            .lcout(sDAC_mem_33Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52215),
            .ce(N__44531),
            .sr(N__51786));
    defparam sDAC_mem_33_2_LC_19_8_2.C_ON=1'b0;
    defparam sDAC_mem_33_2_LC_19_8_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_2_LC_19_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_2_LC_19_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47483),
            .lcout(sDAC_mem_33Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52215),
            .ce(N__44531),
            .sr(N__51786));
    defparam sDAC_mem_33_3_LC_19_8_3.C_ON=1'b0;
    defparam sDAC_mem_33_3_LC_19_8_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_3_LC_19_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_3_LC_19_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46857),
            .lcout(sDAC_mem_33Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52215),
            .ce(N__44531),
            .sr(N__51786));
    defparam sDAC_mem_33_4_LC_19_8_4.C_ON=1'b0;
    defparam sDAC_mem_33_4_LC_19_8_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_4_LC_19_8_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_33_4_LC_19_8_4 (
            .in0(N__45562),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_33Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52215),
            .ce(N__44531),
            .sr(N__51786));
    defparam sDAC_mem_33_5_LC_19_8_5.C_ON=1'b0;
    defparam sDAC_mem_33_5_LC_19_8_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_5_LC_19_8_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_33_5_LC_19_8_5 (
            .in0(N__45065),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_33Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52215),
            .ce(N__44531),
            .sr(N__51786));
    defparam sDAC_mem_33_6_LC_19_8_6.C_ON=1'b0;
    defparam sDAC_mem_33_6_LC_19_8_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_6_LC_19_8_6.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_33_6_LC_19_8_6 (
            .in0(_gnd_net_),
            .in1(N__50465),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_33Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52215),
            .ce(N__44531),
            .sr(N__51786));
    defparam sDAC_mem_33_7_LC_19_8_7.C_ON=1'b0;
    defparam sDAC_mem_33_7_LC_19_8_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_7_LC_19_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_7_LC_19_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50036),
            .lcout(sDAC_mem_33Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52215),
            .ce(N__44531),
            .sr(N__51786));
    defparam sDAC_mem_5_0_LC_19_9_0.C_ON=1'b0;
    defparam sDAC_mem_5_0_LC_19_9_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_0_LC_19_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_0_LC_19_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46383),
            .lcout(sDAC_mem_5Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52210),
            .ce(N__44435),
            .sr(N__51773));
    defparam sDAC_mem_5_1_LC_19_9_1.C_ON=1'b0;
    defparam sDAC_mem_5_1_LC_19_9_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_1_LC_19_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_1_LC_19_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51043),
            .lcout(sDAC_mem_5Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52210),
            .ce(N__44435),
            .sr(N__51773));
    defparam sDAC_mem_5_2_LC_19_9_2.C_ON=1'b0;
    defparam sDAC_mem_5_2_LC_19_9_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_2_LC_19_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_2_LC_19_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47485),
            .lcout(sDAC_mem_5Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52210),
            .ce(N__44435),
            .sr(N__51773));
    defparam sDAC_mem_5_3_LC_19_9_3.C_ON=1'b0;
    defparam sDAC_mem_5_3_LC_19_9_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_3_LC_19_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_3_LC_19_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46856),
            .lcout(sDAC_mem_5Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52210),
            .ce(N__44435),
            .sr(N__51773));
    defparam sDAC_mem_5_4_LC_19_9_4.C_ON=1'b0;
    defparam sDAC_mem_5_4_LC_19_9_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_4_LC_19_9_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_5_4_LC_19_9_4 (
            .in0(N__45563),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_5Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52210),
            .ce(N__44435),
            .sr(N__51773));
    defparam sDAC_mem_5_5_LC_19_9_5.C_ON=1'b0;
    defparam sDAC_mem_5_5_LC_19_9_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_5_LC_19_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_5_LC_19_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45066),
            .lcout(sDAC_mem_5Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52210),
            .ce(N__44435),
            .sr(N__51773));
    defparam sDAC_mem_5_6_LC_19_9_6.C_ON=1'b0;
    defparam sDAC_mem_5_6_LC_19_9_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_6_LC_19_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_6_LC_19_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50466),
            .lcout(sDAC_mem_5Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52210),
            .ce(N__44435),
            .sr(N__51773));
    defparam sDAC_mem_5_7_LC_19_9_7.C_ON=1'b0;
    defparam sDAC_mem_5_7_LC_19_9_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_7_LC_19_9_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_5_7_LC_19_9_7 (
            .in0(_gnd_net_),
            .in1(N__50061),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_5Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52210),
            .ce(N__44435),
            .sr(N__51773));
    defparam sDAC_mem_13_0_LC_19_10_0.C_ON=1'b0;
    defparam sDAC_mem_13_0_LC_19_10_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_0_LC_19_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_0_LC_19_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46345),
            .lcout(sDAC_mem_13Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52206),
            .ce(N__44585),
            .sr(N__51761));
    defparam sDAC_mem_13_1_LC_19_10_1.C_ON=1'b0;
    defparam sDAC_mem_13_1_LC_19_10_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_1_LC_19_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_1_LC_19_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51064),
            .lcout(sDAC_mem_13Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52206),
            .ce(N__44585),
            .sr(N__51761));
    defparam sDAC_mem_13_2_LC_19_10_2.C_ON=1'b0;
    defparam sDAC_mem_13_2_LC_19_10_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_2_LC_19_10_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_13_2_LC_19_10_2 (
            .in0(N__47498),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_13Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52206),
            .ce(N__44585),
            .sr(N__51761));
    defparam sDAC_mem_13_3_LC_19_10_3.C_ON=1'b0;
    defparam sDAC_mem_13_3_LC_19_10_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_3_LC_19_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_3_LC_19_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46906),
            .lcout(sDAC_mem_13Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52206),
            .ce(N__44585),
            .sr(N__51761));
    defparam sDAC_mem_13_4_LC_19_10_4.C_ON=1'b0;
    defparam sDAC_mem_13_4_LC_19_10_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_4_LC_19_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_4_LC_19_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45602),
            .lcout(sDAC_mem_13Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52206),
            .ce(N__44585),
            .sr(N__51761));
    defparam sDAC_mem_13_5_LC_19_10_5.C_ON=1'b0;
    defparam sDAC_mem_13_5_LC_19_10_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_5_LC_19_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_5_LC_19_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45105),
            .lcout(sDAC_mem_13Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52206),
            .ce(N__44585),
            .sr(N__51761));
    defparam sDAC_mem_13_6_LC_19_10_6.C_ON=1'b0;
    defparam sDAC_mem_13_6_LC_19_10_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_6_LC_19_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_6_LC_19_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50526),
            .lcout(sDAC_mem_13Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52206),
            .ce(N__44585),
            .sr(N__51761));
    defparam sDAC_mem_13_7_LC_19_10_7.C_ON=1'b0;
    defparam sDAC_mem_13_7_LC_19_10_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_7_LC_19_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_7_LC_19_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50062),
            .lcout(sDAC_mem_13Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52206),
            .ce(N__44585),
            .sr(N__51761));
    defparam \spi_slave_inst.tx_ready_i_LC_19_11_3 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_ready_i_LC_19_11_3 .SEQ_MODE=4'b1011;
    defparam \spi_slave_inst.tx_ready_i_LC_19_11_3 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \spi_slave_inst.tx_ready_i_LC_19_11_3  (
            .in0(N__51191),
            .in1(N__44557),
            .in2(N__49390),
            .in3(N__51089),
            .lcout(\spi_slave_inst.tx_ready_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52203),
            .ce(),
            .sr(N__51749));
    defparam \spi_slave_inst.txdata_reg_i_4_LC_19_12_0 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_4_LC_19_12_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_4_LC_19_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_4_LC_19_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45824),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52207),
            .ce(),
            .sr(N__51734));
    defparam \spi_slave_inst.txdata_reg_i_0_LC_19_12_1 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_0_LC_19_12_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_0_LC_19_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_0_LC_19_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45815),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52207),
            .ce(),
            .sr(N__51734));
    defparam \spi_slave_inst.txdata_reg_i_2_LC_19_12_4 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_2_LC_19_12_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_2_LC_19_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_2_LC_19_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45806),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52207),
            .ce(),
            .sr(N__51734));
    defparam \spi_slave_inst.txdata_reg_i_1_LC_19_12_7 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_1_LC_19_12_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_1_LC_19_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_1_LC_19_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45791),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52207),
            .ce(),
            .sr(N__51734));
    defparam button_debounce_counter_1_LC_19_13_0.C_ON=1'b0;
    defparam button_debounce_counter_1_LC_19_13_0.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_1_LC_19_13_0.LUT_INIT=16'b0111011110001000;
    LogicCell40 button_debounce_counter_1_LC_19_13_0 (
            .in0(N__45744),
            .in1(N__49240),
            .in2(_gnd_net_),
            .in3(N__45771),
            .lcout(button_debounce_counterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48487),
            .ce(),
            .sr(N__45718));
    defparam button_debounce_counter_0_LC_19_13_1.C_ON=1'b0;
    defparam button_debounce_counter_0_LC_19_13_1.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_0_LC_19_13_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 button_debounce_counter_0_LC_19_13_1 (
            .in0(_gnd_net_),
            .in1(N__49145),
            .in2(_gnd_net_),
            .in3(N__45743),
            .lcout(button_debounce_counterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48487),
            .ce(),
            .sr(N__45718));
    defparam \spi_slave_inst.txdata_reg_i_3_LC_19_14_5 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_3_LC_19_14_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_3_LC_19_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_3_LC_19_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45692),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52216),
            .ce(),
            .sr(N__51711));
    defparam \spi_slave_inst.txdata_reg_i_6_LC_19_14_6 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_6_LC_19_14_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_6_LC_19_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_6_LC_19_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45680),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52216),
            .ce(),
            .sr(N__51711));
    defparam \spi_slave_inst.txdata_reg_i_5_LC_19_14_7 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_5_LC_19_14_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_5_LC_19_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_5_LC_19_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47525),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52216),
            .ce(),
            .sr(N__51711));
    defparam sEEADC_freq_2_LC_19_16_0.C_ON=1'b0;
    defparam sEEADC_freq_2_LC_19_16_0.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_2_LC_19_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEADC_freq_2_LC_19_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47513),
            .lcout(sEEADC_freqZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52231),
            .ce(N__49576),
            .sr(_gnd_net_));
    defparam sEEADC_freq_RNI4KIA1_2_LC_19_16_1.C_ON=1'b0;
    defparam sEEADC_freq_RNI4KIA1_2_LC_19_16_1.SEQ_MODE=4'b0000;
    defparam sEEADC_freq_RNI4KIA1_2_LC_19_16_1.LUT_INIT=16'b1001000000001001;
    LogicCell40 sEEADC_freq_RNI4KIA1_2_LC_19_16_1 (
            .in0(N__47017),
            .in1(N__47006),
            .in2(N__46430),
            .in3(N__46999),
            .lcout(),
            .ltout(un11_sacqtime_NE_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEADC_freq_RNI01BA5_0_LC_19_16_2.C_ON=1'b0;
    defparam sEEADC_freq_RNI01BA5_0_LC_19_16_2.SEQ_MODE=4'b0000;
    defparam sEEADC_freq_RNI01BA5_0_LC_19_16_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 sEEADC_freq_RNI01BA5_0_LC_19_16_2 (
            .in0(N__46988),
            .in1(N__45830),
            .in2(N__46973),
            .in3(N__46397),
            .lcout(un11_sacqtime_NE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEADC_freq_3_LC_19_16_3.C_ON=1'b0;
    defparam sEEADC_freq_3_LC_19_16_3.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_3_LC_19_16_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEADC_freq_3_LC_19_16_3 (
            .in0(N__46765),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEADC_freqZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52231),
            .ce(N__49576),
            .sr(_gnd_net_));
    defparam sEEADC_freq_RNISBIA1_0_LC_19_16_4.C_ON=1'b0;
    defparam sEEADC_freq_RNISBIA1_0_LC_19_16_4.SEQ_MODE=4'b0000;
    defparam sEEADC_freq_RNISBIA1_0_LC_19_16_4.LUT_INIT=16'b1000001001000001;
    LogicCell40 sEEADC_freq_RNISBIA1_0_LC_19_16_4 (
            .in0(N__45872),
            .in1(N__46420),
            .in2(N__45866),
            .in3(N__46408),
            .lcout(un11_sacqtime_NE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEADC_freq_0_LC_19_16_5.C_ON=1'b0;
    defparam sEEADC_freq_0_LC_19_16_5.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_0_LC_19_16_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEADC_freq_0_LC_19_16_5 (
            .in0(N__46316),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEADC_freqZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52231),
            .ce(N__49576),
            .sr(_gnd_net_));
    defparam sEEADC_freq_1_LC_19_16_6.C_ON=1'b0;
    defparam sEEADC_freq_1_LC_19_16_6.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_1_LC_19_16_6.LUT_INIT=16'b1100110011001100;
    LogicCell40 sEEADC_freq_1_LC_19_16_6 (
            .in0(_gnd_net_),
            .in1(N__51019),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEADC_freqZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52231),
            .ce(N__49576),
            .sr(_gnd_net_));
    defparam sEEADC_freq_RNIK4JA1_6_LC_19_16_7.C_ON=1'b0;
    defparam sEEADC_freq_RNIK4JA1_6_LC_19_16_7.SEQ_MODE=4'b0000;
    defparam sEEADC_freq_RNIK4JA1_6_LC_19_16_7.LUT_INIT=16'b1000010000100001;
    LogicCell40 sEEADC_freq_RNIK4JA1_6_LC_19_16_7 (
            .in0(N__50072),
            .in1(N__45856),
            .in2(N__45845),
            .in3(N__49586),
            .lcout(un11_sacqtime_NE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_1_8_LC_19_17_4.C_ON=1'b0;
    defparam RAM_DATA_1_8_LC_19_17_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_8_LC_19_17_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 RAM_DATA_1_8_LC_19_17_4 (
            .in0(N__47717),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RAM_DATA_1Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52241),
            .ce(N__51882),
            .sr(N__51687));
    defparam RAM_DATA_1_9_LC_19_17_5.C_ON=1'b0;
    defparam RAM_DATA_1_9_LC_19_17_5.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_9_LC_19_17_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_9_LC_19_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47678),
            .lcout(RAM_DATA_1Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52241),
            .ce(N__51882),
            .sr(N__51687));
    defparam RAM_DATA_1_12_LC_19_17_7.C_ON=1'b0;
    defparam RAM_DATA_1_12_LC_19_17_7.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_12_LC_19_17_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_12_LC_19_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47636),
            .lcout(RAM_DATA_1Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52241),
            .ce(N__51882),
            .sr(N__51687));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ00Q2_0_LC_20_3_0 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ00Q2_0_LC_20_3_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ00Q2_0_LC_20_3_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ00Q2_0_LC_20_3_0  (
            .in0(_gnd_net_),
            .in1(N__48052),
            .in2(_gnd_net_),
            .in3(N__47782),
            .lcout(spi_miso_ft_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_8_LC_20_4_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_8_LC_20_4_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_8_LC_20_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_8_LC_20_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47582),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48463),
            .ce(),
            .sr(N__51825));
    defparam sCounterDAC_0_LC_20_4_3.C_ON=1'b0;
    defparam sCounterDAC_0_LC_20_4_3.SEQ_MODE=4'b1010;
    defparam sCounterDAC_0_LC_20_4_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 sCounterDAC_0_LC_20_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48126),
            .lcout(sCounterDACZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48463),
            .ce(),
            .sr(N__51825));
    defparam \spi_slave_inst.spi_cs_LC_20_5_6 .C_ON=1'b0;
    defparam \spi_slave_inst.spi_cs_LC_20_5_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.spi_cs_LC_20_5_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \spi_slave_inst.spi_cs_LC_20_5_6  (
            .in0(N__47928),
            .in1(N__48051),
            .in2(_gnd_net_),
            .in3(N__47887),
            .lcout(\spi_slave_inst.spi_csZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_spi_start_LC_20_6_5.C_ON=1'b0;
    defparam sDAC_spi_start_LC_20_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_spi_start_LC_20_6_5.LUT_INIT=16'b1100100011111000;
    LogicCell40 sDAC_spi_start_LC_20_6_5 (
            .in0(N__48554),
            .in1(N__48539),
            .in2(N__47545),
            .in3(N__48140),
            .lcout(sDAC_spi_startZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48466),
            .ce(),
            .sr(N__51816));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIOASC_5_LC_20_7_0 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIOASC_5_LC_20_7_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIOASC_5_LC_20_7_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNIOASC_5_LC_20_7_0  (
            .in0(N__51263),
            .in1(N__51242),
            .in2(N__48689),
            .in3(N__48772),
            .lcout(),
            .ltout(\spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI1DAJ_1_LC_20_7_1 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI1DAJ_1_LC_20_7_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI1DAJ_1_LC_20_7_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNI1DAJ_1_LC_20_7_1  (
            .in0(_gnd_net_),
            .in1(N__48717),
            .in2(N__48059),
            .in3(N__48753),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_i6 ),
            .ltout(\spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1_1_LC_20_7_2 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1_1_LC_20_7_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1_1_LC_20_7_2 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1_1_LC_20_7_2  (
            .in0(N__48056),
            .in1(N__47929),
            .in2(N__47906),
            .in3(N__47888),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIUCSS_1_LC_20_7_3 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIUCSS_1_LC_20_7_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIUCSS_1_LC_20_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNIUCSS_1_LC_20_7_3  (
            .in0(N__47831),
            .in1(N__47816),
            .in2(_gnd_net_),
            .in3(N__48755),
            .lcout(),
            .ltout(\spi_slave_inst.N_1393_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIA0LM2_0_LC_20_7_4 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIA0LM2_0_LC_20_7_4 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIA0LM2_0_LC_20_7_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNIA0LM2_0_LC_20_7_4  (
            .in0(N__47723),
            .in1(N__51178),
            .in2(N__47801),
            .in3(N__48773),
            .lcout(spi_miso),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.txdata_reg_i_RNI1IQC_0_LC_20_7_5 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_RNI1IQC_0_LC_20_7_5 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.txdata_reg_i_RNI1IQC_0_LC_20_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi_slave_inst.txdata_reg_i_RNI1IQC_0_LC_20_7_5  (
            .in0(N__47765),
            .in1(N__47753),
            .in2(_gnd_net_),
            .in3(N__48718),
            .lcout(),
            .ltout(\spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ8SS_1_LC_20_7_6 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ8SS_1_LC_20_7_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ8SS_1_LC_20_7_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ8SS_1_LC_20_7_6  (
            .in0(N__48754),
            .in1(_gnd_net_),
            .in2(N__47741),
            .in3(N__47738),
            .lcout(\spi_slave_inst.N_1396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_RNI9VC2_3_LC_20_8_0.C_ON=1'b0;
    defparam sCounterDAC_RNI9VC2_3_LC_20_8_0.SEQ_MODE=4'b0000;
    defparam sCounterDAC_RNI9VC2_3_LC_20_8_0.LUT_INIT=16'b0000000011001100;
    LogicCell40 sCounterDAC_RNI9VC2_3_LC_20_8_0 (
            .in0(_gnd_net_),
            .in1(N__48668),
            .in2(_gnd_net_),
            .in3(N__48127),
            .lcout(m15_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_1_LC_20_9_0.C_ON=1'b0;
    defparam sCounterDAC_1_LC_20_9_0.SEQ_MODE=4'b1010;
    defparam sCounterDAC_1_LC_20_9_0.LUT_INIT=16'b1010010101011010;
    LogicCell40 sCounterDAC_1_LC_20_9_0 (
            .in0(N__48131),
            .in1(_gnd_net_),
            .in2(N__48097),
            .in3(_gnd_net_),
            .lcout(sCounterDACZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48477),
            .ce(),
            .sr(N__51787));
    defparam sCounterDAC_RNIHIJ3_1_LC_20_9_1.C_ON=1'b0;
    defparam sCounterDAC_RNIHIJ3_1_LC_20_9_1.SEQ_MODE=4'b0000;
    defparam sCounterDAC_RNIHIJ3_1_LC_20_9_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 sCounterDAC_RNIHIJ3_1_LC_20_9_1 (
            .in0(N__48637),
            .in1(N__48090),
            .in2(_gnd_net_),
            .in3(N__48665),
            .lcout(m8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_RNI4HQ4_9_LC_20_9_2.C_ON=1'b0;
    defparam sCounterDAC_RNI4HQ4_9_LC_20_9_2.SEQ_MODE=4'b0000;
    defparam sCounterDAC_RNI4HQ4_9_LC_20_9_2.LUT_INIT=16'b0000000000000100;
    LogicCell40 sCounterDAC_RNI4HQ4_9_LC_20_9_2 (
            .in0(N__48568),
            .in1(N__48073),
            .in2(N__48509),
            .in3(N__48591),
            .lcout(N_23_mux),
            .ltout(N_23_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_RNIFI77_1_LC_20_9_3.C_ON=1'b0;
    defparam sCounterDAC_RNIFI77_1_LC_20_9_3.SEQ_MODE=4'b0000;
    defparam sCounterDAC_RNIFI77_1_LC_20_9_3.LUT_INIT=16'b0001000000010000;
    LogicCell40 sCounterDAC_RNIFI77_1_LC_20_9_3 (
            .in0(N__48636),
            .in1(N__48089),
            .in2(N__48191),
            .in3(_gnd_net_),
            .lcout(N_25_mux),
            .ltout(N_25_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_RNIBR1C_5_LC_20_9_4.C_ON=1'b0;
    defparam sCounterDAC_RNIBR1C_5_LC_20_9_4.SEQ_MODE=4'b0000;
    defparam sCounterDAC_RNIBR1C_5_LC_20_9_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 sCounterDAC_RNIBR1C_5_LC_20_9_4 (
            .in0(N__48533),
            .in1(N__48611),
            .in2(N__48188),
            .in3(N__48185),
            .lcout(op_eq_scounterdac10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_RNI05RA_5_LC_20_9_5.C_ON=1'b0;
    defparam sCounterDAC_RNI05RA_5_LC_20_9_5.SEQ_MODE=4'b0000;
    defparam sCounterDAC_RNI05RA_5_LC_20_9_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 sCounterDAC_RNI05RA_5_LC_20_9_5 (
            .in0(N__48161),
            .in1(N__48155),
            .in2(N__48619),
            .in3(N__48129),
            .lcout(N_30_mux),
            .ltout(N_30_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_6_LC_20_9_6.C_ON=1'b0;
    defparam sCounterDAC_6_LC_20_9_6.SEQ_MODE=4'b1010;
    defparam sCounterDAC_6_LC_20_9_6.LUT_INIT=16'b0001001101001100;
    LogicCell40 sCounterDAC_6_LC_20_9_6 (
            .in0(N__48534),
            .in1(N__48578),
            .in2(N__48149),
            .in3(N__48592),
            .lcout(sCounterDACZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48477),
            .ce(),
            .sr(N__51787));
    defparam sDAC_spi_start_RNO_0_LC_20_9_7.C_ON=1'b0;
    defparam sDAC_spi_start_RNO_0_LC_20_9_7.SEQ_MODE=4'b0000;
    defparam sDAC_spi_start_RNO_0_LC_20_9_7.LUT_INIT=16'b0000010000000000;
    LogicCell40 sDAC_spi_start_RNO_0_LC_20_9_7 (
            .in0(N__48667),
            .in1(N__48130),
            .in2(N__48620),
            .in3(N__48146),
            .lcout(N_32_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_scounterdac_cry_1_c_LC_20_10_0.C_ON=1'b1;
    defparam un2_scounterdac_cry_1_c_LC_20_10_0.SEQ_MODE=4'b0000;
    defparam un2_scounterdac_cry_1_c_LC_20_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_scounterdac_cry_1_c_LC_20_10_0 (
            .in0(_gnd_net_),
            .in1(N__48128),
            .in2(N__48098),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_20_10_0_),
            .carryout(un2_scounterdac_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_2_LC_20_10_1.C_ON=1'b1;
    defparam sCounterDAC_2_LC_20_10_1.SEQ_MODE=4'b1010;
    defparam sCounterDAC_2_LC_20_10_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 sCounterDAC_2_LC_20_10_1 (
            .in0(_gnd_net_),
            .in1(N__48074),
            .in2(_gnd_net_),
            .in3(N__48062),
            .lcout(sCounterDACZ0Z_2),
            .ltout(),
            .carryin(un2_scounterdac_cry_1),
            .carryout(un2_scounterdac_cry_2),
            .clk(N__48481),
            .ce(),
            .sr(N__51774));
    defparam sCounterDAC_3_LC_20_10_2.C_ON=1'b1;
    defparam sCounterDAC_3_LC_20_10_2.SEQ_MODE=4'b1010;
    defparam sCounterDAC_3_LC_20_10_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 sCounterDAC_3_LC_20_10_2 (
            .in0(_gnd_net_),
            .in1(N__48666),
            .in2(_gnd_net_),
            .in3(N__48641),
            .lcout(sCounterDACZ0Z_3),
            .ltout(),
            .carryin(un2_scounterdac_cry_2),
            .carryout(un2_scounterdac_cry_3),
            .clk(N__48481),
            .ce(),
            .sr(N__51774));
    defparam sCounterDAC_4_LC_20_10_3.C_ON=1'b1;
    defparam sCounterDAC_4_LC_20_10_3.SEQ_MODE=4'b1010;
    defparam sCounterDAC_4_LC_20_10_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 sCounterDAC_4_LC_20_10_3 (
            .in0(_gnd_net_),
            .in1(N__48638),
            .in2(_gnd_net_),
            .in3(N__48623),
            .lcout(sCounterDACZ0Z_4),
            .ltout(),
            .carryin(un2_scounterdac_cry_3),
            .carryout(un2_scounterdac_cry_4),
            .clk(N__48481),
            .ce(),
            .sr(N__51774));
    defparam sCounterDAC_5_LC_20_10_4.C_ON=1'b1;
    defparam sCounterDAC_5_LC_20_10_4.SEQ_MODE=4'b1010;
    defparam sCounterDAC_5_LC_20_10_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 sCounterDAC_5_LC_20_10_4 (
            .in0(_gnd_net_),
            .in1(N__48618),
            .in2(_gnd_net_),
            .in3(N__48596),
            .lcout(sCounterDACZ0Z_5),
            .ltout(),
            .carryin(un2_scounterdac_cry_4),
            .carryout(un2_scounterdac_cry_5),
            .clk(N__48481),
            .ce(),
            .sr(N__51774));
    defparam un2_scounterdac_cry_5_THRU_LUT4_0_LC_20_10_5.C_ON=1'b1;
    defparam un2_scounterdac_cry_5_THRU_LUT4_0_LC_20_10_5.SEQ_MODE=4'b0000;
    defparam un2_scounterdac_cry_5_THRU_LUT4_0_LC_20_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_scounterdac_cry_5_THRU_LUT4_0_LC_20_10_5 (
            .in0(_gnd_net_),
            .in1(N__48593),
            .in2(_gnd_net_),
            .in3(N__48572),
            .lcout(un2_scounterdac_cry_5_THRU_CO),
            .ltout(),
            .carryin(un2_scounterdac_cry_5),
            .carryout(un2_scounterdac_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_7_LC_20_10_6.C_ON=1'b1;
    defparam sCounterDAC_7_LC_20_10_6.SEQ_MODE=4'b1010;
    defparam sCounterDAC_7_LC_20_10_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 sCounterDAC_7_LC_20_10_6 (
            .in0(_gnd_net_),
            .in1(N__48569),
            .in2(_gnd_net_),
            .in3(N__48557),
            .lcout(sCounterDACZ0Z_7),
            .ltout(),
            .carryin(un2_scounterdac_cry_6),
            .carryout(un2_scounterdac_cry_7),
            .clk(N__48481),
            .ce(),
            .sr(N__51774));
    defparam sCounterDAC_8_LC_20_10_7.C_ON=1'b1;
    defparam sCounterDAC_8_LC_20_10_7.SEQ_MODE=4'b1010;
    defparam sCounterDAC_8_LC_20_10_7.LUT_INIT=16'b0011001101000100;
    LogicCell40 sCounterDAC_8_LC_20_10_7 (
            .in0(N__48553),
            .in1(N__48535),
            .in2(_gnd_net_),
            .in3(N__48515),
            .lcout(sCounterDACZ0Z_8),
            .ltout(),
            .carryin(un2_scounterdac_cry_7),
            .carryout(un2_scounterdac_cry_8),
            .clk(N__48481),
            .ce(),
            .sr(N__51774));
    defparam sCounterDAC_9_LC_20_11_0.C_ON=1'b0;
    defparam sCounterDAC_9_LC_20_11_0.SEQ_MODE=4'b1010;
    defparam sCounterDAC_9_LC_20_11_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 sCounterDAC_9_LC_20_11_0 (
            .in0(_gnd_net_),
            .in1(N__48505),
            .in2(_gnd_net_),
            .in3(N__48512),
            .lcout(sCounterDACZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48484),
            .ce(),
            .sr(N__51762));
    defparam \spi_slave_inst.rx_done_pos_sclk_i_LC_20_13_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_pos_sclk_i_LC_20_13_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_done_pos_sclk_i_LC_20_13_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \spi_slave_inst.rx_done_pos_sclk_i_LC_20_13_0  (
            .in0(N__48341),
            .in1(N__48328),
            .in2(_gnd_net_),
            .in3(N__48305),
            .lcout(\spi_slave_inst.rx_done_pos_sclk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__48266),
            .ce(N__48232),
            .sr(N__51735));
    defparam \spi_slave_inst.txdata_reg_i_7_LC_20_15_1 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_7_LC_20_15_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_7_LC_20_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_7_LC_20_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50570),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52217),
            .ce(),
            .sr(N__51712));
    defparam sEEADC_freq_6_LC_20_16_0.C_ON=1'b0;
    defparam sEEADC_freq_6_LC_20_16_0.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_6_LC_20_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEADC_freq_6_LC_20_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50480),
            .lcout(sEEADC_freqZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52223),
            .ce(N__49580),
            .sr(_gnd_net_));
    defparam sEEADC_freq_7_LC_20_16_1.C_ON=1'b0;
    defparam sEEADC_freq_7_LC_20_16_1.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_7_LC_20_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEADC_freq_7_LC_20_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50048),
            .lcout(sEEADC_freqZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52223),
            .ce(N__49580),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_5_15_LC_20_17_3.C_ON=1'b0;
    defparam RAM_DATA_cl_5_15_LC_20_17_3.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_5_15_LC_20_17_3.LUT_INIT=16'b1011000000000000;
    LogicCell40 RAM_DATA_cl_5_15_LC_20_17_3 (
            .in0(N__48802),
            .in1(N__49494),
            .in2(N__49434),
            .in3(N__48956),
            .lcout(RAM_DATA_cl_5Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52232),
            .ce(),
            .sr(N__51693));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_0_LC_22_7_0 .C_ON=1'b1;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_0_LC_22_7_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_0_LC_22_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_0_LC_22_7_0  (
            .in0(N__51143),
            .in1(N__48771),
            .in2(N__48791),
            .in3(N__48790),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0 ),
            .ltout(),
            .carryin(bfn_22_7_0_),
            .carryout(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0 ),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51821));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_1_LC_22_7_1 .C_ON=1'b1;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_1_LC_22_7_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_1_LC_22_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_1_LC_22_7_1  (
            .in0(N__51145),
            .in1(N__48752),
            .in2(_gnd_net_),
            .in3(N__48734),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0 ),
            .carryout(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1 ),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51821));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_2_LC_22_7_2 .C_ON=1'b1;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_2_LC_22_7_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_2_LC_22_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_2_LC_22_7_2  (
            .in0(N__51144),
            .in1(N__48713),
            .in2(_gnd_net_),
            .in3(N__48692),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1 ),
            .carryout(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2 ),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51821));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_3_LC_22_7_3 .C_ON=1'b1;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_3_LC_22_7_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_3_LC_22_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_3_LC_22_7_3  (
            .in0(_gnd_net_),
            .in1(N__48685),
            .in2(_gnd_net_),
            .in3(N__48671),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2 ),
            .carryout(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3 ),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51821));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_4_LC_22_7_4 .C_ON=1'b1;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_4_LC_22_7_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_4_LC_22_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_4_LC_22_7_4  (
            .in0(_gnd_net_),
            .in1(N__51262),
            .in2(_gnd_net_),
            .in3(N__51248),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3 ),
            .carryout(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4 ),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51821));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_5_LC_22_7_5 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_5_LC_22_7_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_5_LC_22_7_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_5_LC_22_7_5  (
            .in0(_gnd_net_),
            .in1(N__51241),
            .in2(_gnd_net_),
            .in3(N__51245),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51821));
    defparam \spi_slave_inst.tx_done_neg_sclk_i_LC_22_7_6 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_done_neg_sclk_i_LC_22_7_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_done_neg_sclk_i_LC_22_7_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \spi_slave_inst.tx_done_neg_sclk_i_LC_22_7_6  (
            .in0(N__51197),
            .in1(N__51124),
            .in2(_gnd_net_),
            .in3(N__51146),
            .lcout(\spi_slave_inst.tx_done_neg_sclk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__51821));
    defparam \spi_slave_inst.tx_done_reg1_i_LC_22_8_5 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_done_reg1_i_LC_22_8_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_done_reg1_i_LC_22_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.tx_done_reg1_i_LC_22_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51125),
            .lcout(\spi_slave_inst.tx_done_reg1_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52204),
            .ce(),
            .sr(N__51817));
    defparam \spi_slave_inst.tx_done_reg2_i_LC_22_9_2 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_done_reg2_i_LC_22_9_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_done_reg2_i_LC_22_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.tx_done_reg2_i_LC_22_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51113),
            .lcout(\spi_slave_inst.tx_done_reg2_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52202),
            .ce(),
            .sr(N__51809));
    defparam \spi_slave_inst.tx_done_reg3_i_LC_22_9_5 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_done_reg3_i_LC_22_9_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_done_reg3_i_LC_22_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.tx_done_reg3_i_LC_22_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51101),
            .lcout(\spi_slave_inst.tx_done_reg3_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52202),
            .ce(),
            .sr(N__51809));
    defparam CONSTANT_ONE_LUT4_LC_22_10_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_22_10_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_22_10_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_22_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_ready_i_RNO_0_LC_22_10_7 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_ready_i_RNO_0_LC_22_10_7 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_ready_i_RNO_0_LC_22_10_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \spi_slave_inst.tx_ready_i_RNO_0_LC_22_10_7  (
            .in0(_gnd_net_),
            .in1(N__51107),
            .in2(_gnd_net_),
            .in3(N__51100),
            .lcout(\spi_slave_inst.un4_tx_done_reg2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_25_1_LC_22_12_0.C_ON=1'b0;
    defparam sDAC_mem_25_1_LC_22_12_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_1_LC_22_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_1_LC_22_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51029),
            .lcout(sDAC_mem_25Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52201),
            .ce(N__50594),
            .sr(N__51775));
    defparam RAM_DATA_1_15_LC_23_17_4.C_ON=1'b0;
    defparam RAM_DATA_1_15_LC_23_17_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_15_LC_23_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_15_LC_23_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52408),
            .lcout(RAM_DATA_1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52211),
            .ce(N__51894),
            .sr(N__51722));
endmodule // MATTY_MAIN_VHDL
