pll256M2_inst: pll256M2
port map(
          REFERENCECLK => ,
          PLLOUTCOREA => ,
          PLLOUTCOREB => ,
          PLLOUTGLOBALA => ,
          PLLOUTGLOBALB => ,
          RESET => 
        );
