-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Oct 7 2018 03:23:07

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MATTY_MAIN_VHDL" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MATTY_MAIN_VHDL
entity MATTY_MAIN_VHDL is
port (
    RAM_DATA : inout std_logic_vector(15 downto 0);
    RAM_ADD : out std_logic_vector(18 downto 0);
    spi_sclk_ft : in std_logic;
    button_trig : in std_logic;
    ADC9 : in std_logic;
    spi_cs_ft : in std_logic;
    poff : out std_logic;
    RAM_nOE : out std_logic;
    ADC0 : in std_logic;
    spi_mosi_flash : out std_logic;
    spi_miso_flash : in std_logic;
    trig_ft : in std_logic;
    spi_miso_rpi : out std_logic;
    RAM_nWE : out std_logic;
    DAC_cs : out std_logic;
    ADC6 : in std_logic;
    spi_select : in std_logic;
    clk : in std_logic;
    ADC4 : in std_logic;
    trig_rpi : in std_logic;
    top_tour2 : in std_logic;
    spi_cs_rpi : in std_logic;
    DAC_sclk : out std_logic;
    ADC_clk : out std_logic;
    ADC3 : in std_logic;
    trig_ext : in std_logic;
    spi_mosi_rpi : in std_logic;
    spi_mosi_ft : in std_logic;
    cs_rpi2flash : in std_logic;
    spi_cs_flash : out std_logic;
    pon : out std_logic;
    RAM_nCE : out std_logic;
    LED3 : out std_logic;
    ADC1 : in std_logic;
    reset_rpi : in std_logic;
    RAM_nLB : out std_logic;
    LED_MODE : out std_logic;
    ADC8 : in std_logic;
    spi_sclk_rpi : in std_logic;
    ADC7 : in std_logic;
    top_tour1 : in std_logic;
    spi_miso_ft : out std_logic;
    button_mode : in std_logic;
    DAC_mosi : out std_logic;
    ADC5 : in std_logic;
    reset_ft : in std_logic;
    LED_ACQ : out std_logic;
    spi_sclk_flash : out std_logic;
    reset_alim : in std_logic;
    RAM_nUB : out std_logic;
    ADC2 : in std_logic);
end MATTY_MAIN_VHDL;

-- Architecture of MATTY_MAIN_VHDL
-- View name is \INTERFACE\
architecture \INTERFACE\ of MATTY_MAIN_VHDL is

signal \N__53520\ : std_logic;
signal \N__53519\ : std_logic;
signal \N__53518\ : std_logic;
signal \N__53511\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53509\ : std_logic;
signal \N__53502\ : std_logic;
signal \N__53501\ : std_logic;
signal \N__53500\ : std_logic;
signal \N__53493\ : std_logic;
signal \N__53492\ : std_logic;
signal \N__53491\ : std_logic;
signal \N__53484\ : std_logic;
signal \N__53483\ : std_logic;
signal \N__53482\ : std_logic;
signal \N__53475\ : std_logic;
signal \N__53474\ : std_logic;
signal \N__53473\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53465\ : std_logic;
signal \N__53464\ : std_logic;
signal \N__53457\ : std_logic;
signal \N__53456\ : std_logic;
signal \N__53455\ : std_logic;
signal \N__53448\ : std_logic;
signal \N__53447\ : std_logic;
signal \N__53446\ : std_logic;
signal \N__53439\ : std_logic;
signal \N__53438\ : std_logic;
signal \N__53437\ : std_logic;
signal \N__53430\ : std_logic;
signal \N__53429\ : std_logic;
signal \N__53428\ : std_logic;
signal \N__53421\ : std_logic;
signal \N__53420\ : std_logic;
signal \N__53419\ : std_logic;
signal \N__53412\ : std_logic;
signal \N__53411\ : std_logic;
signal \N__53410\ : std_logic;
signal \N__53403\ : std_logic;
signal \N__53402\ : std_logic;
signal \N__53401\ : std_logic;
signal \N__53394\ : std_logic;
signal \N__53393\ : std_logic;
signal \N__53392\ : std_logic;
signal \N__53385\ : std_logic;
signal \N__53384\ : std_logic;
signal \N__53383\ : std_logic;
signal \N__53376\ : std_logic;
signal \N__53375\ : std_logic;
signal \N__53374\ : std_logic;
signal \N__53367\ : std_logic;
signal \N__53366\ : std_logic;
signal \N__53365\ : std_logic;
signal \N__53358\ : std_logic;
signal \N__53357\ : std_logic;
signal \N__53356\ : std_logic;
signal \N__53349\ : std_logic;
signal \N__53348\ : std_logic;
signal \N__53347\ : std_logic;
signal \N__53340\ : std_logic;
signal \N__53339\ : std_logic;
signal \N__53338\ : std_logic;
signal \N__53331\ : std_logic;
signal \N__53330\ : std_logic;
signal \N__53329\ : std_logic;
signal \N__53322\ : std_logic;
signal \N__53321\ : std_logic;
signal \N__53320\ : std_logic;
signal \N__53313\ : std_logic;
signal \N__53312\ : std_logic;
signal \N__53311\ : std_logic;
signal \N__53304\ : std_logic;
signal \N__53303\ : std_logic;
signal \N__53302\ : std_logic;
signal \N__53295\ : std_logic;
signal \N__53294\ : std_logic;
signal \N__53293\ : std_logic;
signal \N__53286\ : std_logic;
signal \N__53285\ : std_logic;
signal \N__53284\ : std_logic;
signal \N__53277\ : std_logic;
signal \N__53276\ : std_logic;
signal \N__53275\ : std_logic;
signal \N__53268\ : std_logic;
signal \N__53267\ : std_logic;
signal \N__53266\ : std_logic;
signal \N__53259\ : std_logic;
signal \N__53258\ : std_logic;
signal \N__53257\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53249\ : std_logic;
signal \N__53248\ : std_logic;
signal \N__53241\ : std_logic;
signal \N__53240\ : std_logic;
signal \N__53239\ : std_logic;
signal \N__53232\ : std_logic;
signal \N__53231\ : std_logic;
signal \N__53230\ : std_logic;
signal \N__53223\ : std_logic;
signal \N__53222\ : std_logic;
signal \N__53221\ : std_logic;
signal \N__53214\ : std_logic;
signal \N__53213\ : std_logic;
signal \N__53212\ : std_logic;
signal \N__53205\ : std_logic;
signal \N__53204\ : std_logic;
signal \N__53203\ : std_logic;
signal \N__53196\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53194\ : std_logic;
signal \N__53187\ : std_logic;
signal \N__53186\ : std_logic;
signal \N__53185\ : std_logic;
signal \N__53178\ : std_logic;
signal \N__53177\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53169\ : std_logic;
signal \N__53168\ : std_logic;
signal \N__53167\ : std_logic;
signal \N__53160\ : std_logic;
signal \N__53159\ : std_logic;
signal \N__53158\ : std_logic;
signal \N__53151\ : std_logic;
signal \N__53150\ : std_logic;
signal \N__53149\ : std_logic;
signal \N__53142\ : std_logic;
signal \N__53141\ : std_logic;
signal \N__53140\ : std_logic;
signal \N__53133\ : std_logic;
signal \N__53132\ : std_logic;
signal \N__53131\ : std_logic;
signal \N__53124\ : std_logic;
signal \N__53123\ : std_logic;
signal \N__53122\ : std_logic;
signal \N__53115\ : std_logic;
signal \N__53114\ : std_logic;
signal \N__53113\ : std_logic;
signal \N__53106\ : std_logic;
signal \N__53105\ : std_logic;
signal \N__53104\ : std_logic;
signal \N__53097\ : std_logic;
signal \N__53096\ : std_logic;
signal \N__53095\ : std_logic;
signal \N__53088\ : std_logic;
signal \N__53087\ : std_logic;
signal \N__53086\ : std_logic;
signal \N__53079\ : std_logic;
signal \N__53078\ : std_logic;
signal \N__53077\ : std_logic;
signal \N__53070\ : std_logic;
signal \N__53069\ : std_logic;
signal \N__53068\ : std_logic;
signal \N__53061\ : std_logic;
signal \N__53060\ : std_logic;
signal \N__53059\ : std_logic;
signal \N__53052\ : std_logic;
signal \N__53051\ : std_logic;
signal \N__53050\ : std_logic;
signal \N__53043\ : std_logic;
signal \N__53042\ : std_logic;
signal \N__53041\ : std_logic;
signal \N__53034\ : std_logic;
signal \N__53033\ : std_logic;
signal \N__53032\ : std_logic;
signal \N__53025\ : std_logic;
signal \N__53024\ : std_logic;
signal \N__53023\ : std_logic;
signal \N__53016\ : std_logic;
signal \N__53015\ : std_logic;
signal \N__53014\ : std_logic;
signal \N__53007\ : std_logic;
signal \N__53006\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__52998\ : std_logic;
signal \N__52997\ : std_logic;
signal \N__52996\ : std_logic;
signal \N__52989\ : std_logic;
signal \N__52988\ : std_logic;
signal \N__52987\ : std_logic;
signal \N__52980\ : std_logic;
signal \N__52979\ : std_logic;
signal \N__52978\ : std_logic;
signal \N__52971\ : std_logic;
signal \N__52970\ : std_logic;
signal \N__52969\ : std_logic;
signal \N__52962\ : std_logic;
signal \N__52961\ : std_logic;
signal \N__52960\ : std_logic;
signal \N__52953\ : std_logic;
signal \N__52952\ : std_logic;
signal \N__52951\ : std_logic;
signal \N__52944\ : std_logic;
signal \N__52943\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52935\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52933\ : std_logic;
signal \N__52926\ : std_logic;
signal \N__52925\ : std_logic;
signal \N__52924\ : std_logic;
signal \N__52917\ : std_logic;
signal \N__52916\ : std_logic;
signal \N__52915\ : std_logic;
signal \N__52908\ : std_logic;
signal \N__52907\ : std_logic;
signal \N__52906\ : std_logic;
signal \N__52899\ : std_logic;
signal \N__52898\ : std_logic;
signal \N__52897\ : std_logic;
signal \N__52890\ : std_logic;
signal \N__52889\ : std_logic;
signal \N__52888\ : std_logic;
signal \N__52881\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52879\ : std_logic;
signal \N__52872\ : std_logic;
signal \N__52871\ : std_logic;
signal \N__52870\ : std_logic;
signal \N__52863\ : std_logic;
signal \N__52862\ : std_logic;
signal \N__52861\ : std_logic;
signal \N__52854\ : std_logic;
signal \N__52853\ : std_logic;
signal \N__52852\ : std_logic;
signal \N__52845\ : std_logic;
signal \N__52844\ : std_logic;
signal \N__52843\ : std_logic;
signal \N__52836\ : std_logic;
signal \N__52835\ : std_logic;
signal \N__52834\ : std_logic;
signal \N__52827\ : std_logic;
signal \N__52826\ : std_logic;
signal \N__52825\ : std_logic;
signal \N__52818\ : std_logic;
signal \N__52817\ : std_logic;
signal \N__52816\ : std_logic;
signal \N__52809\ : std_logic;
signal \N__52808\ : std_logic;
signal \N__52807\ : std_logic;
signal \N__52790\ : std_logic;
signal \N__52789\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52787\ : std_logic;
signal \N__52786\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52784\ : std_logic;
signal \N__52783\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52781\ : std_logic;
signal \N__52780\ : std_logic;
signal \N__52779\ : std_logic;
signal \N__52770\ : std_logic;
signal \N__52769\ : std_logic;
signal \N__52768\ : std_logic;
signal \N__52767\ : std_logic;
signal \N__52766\ : std_logic;
signal \N__52765\ : std_logic;
signal \N__52764\ : std_logic;
signal \N__52763\ : std_logic;
signal \N__52760\ : std_logic;
signal \N__52759\ : std_logic;
signal \N__52756\ : std_logic;
signal \N__52755\ : std_logic;
signal \N__52752\ : std_logic;
signal \N__52751\ : std_logic;
signal \N__52748\ : std_logic;
signal \N__52747\ : std_logic;
signal \N__52746\ : std_logic;
signal \N__52745\ : std_logic;
signal \N__52744\ : std_logic;
signal \N__52743\ : std_logic;
signal \N__52742\ : std_logic;
signal \N__52739\ : std_logic;
signal \N__52738\ : std_logic;
signal \N__52731\ : std_logic;
signal \N__52728\ : std_logic;
signal \N__52721\ : std_logic;
signal \N__52712\ : std_logic;
signal \N__52711\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52709\ : std_logic;
signal \N__52708\ : std_logic;
signal \N__52707\ : std_logic;
signal \N__52706\ : std_logic;
signal \N__52705\ : std_logic;
signal \N__52688\ : std_logic;
signal \N__52685\ : std_logic;
signal \N__52684\ : std_logic;
signal \N__52681\ : std_logic;
signal \N__52680\ : std_logic;
signal \N__52677\ : std_logic;
signal \N__52676\ : std_logic;
signal \N__52673\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52671\ : std_logic;
signal \N__52670\ : std_logic;
signal \N__52669\ : std_logic;
signal \N__52668\ : std_logic;
signal \N__52661\ : std_logic;
signal \N__52658\ : std_logic;
signal \N__52651\ : std_logic;
signal \N__52650\ : std_logic;
signal \N__52649\ : std_logic;
signal \N__52646\ : std_logic;
signal \N__52643\ : std_logic;
signal \N__52640\ : std_logic;
signal \N__52639\ : std_logic;
signal \N__52636\ : std_logic;
signal \N__52633\ : std_logic;
signal \N__52630\ : std_logic;
signal \N__52627\ : std_logic;
signal \N__52626\ : std_logic;
signal \N__52625\ : std_logic;
signal \N__52624\ : std_logic;
signal \N__52623\ : std_logic;
signal \N__52620\ : std_logic;
signal \N__52603\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52599\ : std_logic;
signal \N__52598\ : std_logic;
signal \N__52595\ : std_logic;
signal \N__52594\ : std_logic;
signal \N__52591\ : std_logic;
signal \N__52590\ : std_logic;
signal \N__52587\ : std_logic;
signal \N__52586\ : std_logic;
signal \N__52579\ : std_logic;
signal \N__52574\ : std_logic;
signal \N__52573\ : std_logic;
signal \N__52572\ : std_logic;
signal \N__52571\ : std_logic;
signal \N__52570\ : std_logic;
signal \N__52563\ : std_logic;
signal \N__52552\ : std_logic;
signal \N__52549\ : std_logic;
signal \N__52548\ : std_logic;
signal \N__52545\ : std_logic;
signal \N__52544\ : std_logic;
signal \N__52541\ : std_logic;
signal \N__52540\ : std_logic;
signal \N__52537\ : std_logic;
signal \N__52536\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52514\ : std_logic;
signal \N__52511\ : std_logic;
signal \N__52510\ : std_logic;
signal \N__52507\ : std_logic;
signal \N__52504\ : std_logic;
signal \N__52503\ : std_logic;
signal \N__52500\ : std_logic;
signal \N__52499\ : std_logic;
signal \N__52496\ : std_logic;
signal \N__52495\ : std_logic;
signal \N__52492\ : std_logic;
signal \N__52491\ : std_logic;
signal \N__52488\ : std_logic;
signal \N__52485\ : std_logic;
signal \N__52482\ : std_logic;
signal \N__52465\ : std_logic;
signal \N__52460\ : std_logic;
signal \N__52455\ : std_logic;
signal \N__52450\ : std_logic;
signal \N__52433\ : std_logic;
signal \N__52428\ : std_logic;
signal \N__52425\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52417\ : std_logic;
signal \N__52414\ : std_logic;
signal \N__52409\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52405\ : std_logic;
signal \N__52402\ : std_logic;
signal \N__52399\ : std_logic;
signal \N__52396\ : std_logic;
signal \N__52393\ : std_logic;
signal \N__52390\ : std_logic;
signal \N__52385\ : std_logic;
signal \N__52380\ : std_logic;
signal \N__52377\ : std_logic;
signal \N__52372\ : std_logic;
signal \N__52367\ : std_logic;
signal \N__52364\ : std_logic;
signal \N__52361\ : std_logic;
signal \N__52358\ : std_logic;
signal \N__52355\ : std_logic;
signal \N__52352\ : std_logic;
signal \N__52349\ : std_logic;
signal \N__52348\ : std_logic;
signal \N__52347\ : std_logic;
signal \N__52346\ : std_logic;
signal \N__52345\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52343\ : std_logic;
signal \N__52342\ : std_logic;
signal \N__52341\ : std_logic;
signal \N__52340\ : std_logic;
signal \N__52339\ : std_logic;
signal \N__52338\ : std_logic;
signal \N__52337\ : std_logic;
signal \N__52336\ : std_logic;
signal \N__52335\ : std_logic;
signal \N__52334\ : std_logic;
signal \N__52333\ : std_logic;
signal \N__52332\ : std_logic;
signal \N__52331\ : std_logic;
signal \N__52330\ : std_logic;
signal \N__52329\ : std_logic;
signal \N__52328\ : std_logic;
signal \N__52327\ : std_logic;
signal \N__52326\ : std_logic;
signal \N__52325\ : std_logic;
signal \N__52324\ : std_logic;
signal \N__52323\ : std_logic;
signal \N__52322\ : std_logic;
signal \N__52321\ : std_logic;
signal \N__52320\ : std_logic;
signal \N__52319\ : std_logic;
signal \N__52318\ : std_logic;
signal \N__52317\ : std_logic;
signal \N__52316\ : std_logic;
signal \N__52315\ : std_logic;
signal \N__52314\ : std_logic;
signal \N__52313\ : std_logic;
signal \N__52312\ : std_logic;
signal \N__52311\ : std_logic;
signal \N__52310\ : std_logic;
signal \N__52309\ : std_logic;
signal \N__52308\ : std_logic;
signal \N__52307\ : std_logic;
signal \N__52306\ : std_logic;
signal \N__52305\ : std_logic;
signal \N__52304\ : std_logic;
signal \N__52303\ : std_logic;
signal \N__52302\ : std_logic;
signal \N__52301\ : std_logic;
signal \N__52300\ : std_logic;
signal \N__52299\ : std_logic;
signal \N__52298\ : std_logic;
signal \N__52297\ : std_logic;
signal \N__52296\ : std_logic;
signal \N__52295\ : std_logic;
signal \N__52294\ : std_logic;
signal \N__52293\ : std_logic;
signal \N__52292\ : std_logic;
signal \N__52291\ : std_logic;
signal \N__52290\ : std_logic;
signal \N__52289\ : std_logic;
signal \N__52288\ : std_logic;
signal \N__52287\ : std_logic;
signal \N__52286\ : std_logic;
signal \N__52285\ : std_logic;
signal \N__52284\ : std_logic;
signal \N__52283\ : std_logic;
signal \N__52282\ : std_logic;
signal \N__52281\ : std_logic;
signal \N__52280\ : std_logic;
signal \N__52279\ : std_logic;
signal \N__52278\ : std_logic;
signal \N__52277\ : std_logic;
signal \N__52276\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52274\ : std_logic;
signal \N__52273\ : std_logic;
signal \N__52272\ : std_logic;
signal \N__52271\ : std_logic;
signal \N__52270\ : std_logic;
signal \N__52269\ : std_logic;
signal \N__52268\ : std_logic;
signal \N__52267\ : std_logic;
signal \N__52266\ : std_logic;
signal \N__52265\ : std_logic;
signal \N__52264\ : std_logic;
signal \N__52263\ : std_logic;
signal \N__52262\ : std_logic;
signal \N__52261\ : std_logic;
signal \N__52260\ : std_logic;
signal \N__52259\ : std_logic;
signal \N__52258\ : std_logic;
signal \N__52257\ : std_logic;
signal \N__52256\ : std_logic;
signal \N__52255\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52253\ : std_logic;
signal \N__52252\ : std_logic;
signal \N__52251\ : std_logic;
signal \N__52250\ : std_logic;
signal \N__52249\ : std_logic;
signal \N__52248\ : std_logic;
signal \N__52247\ : std_logic;
signal \N__52246\ : std_logic;
signal \N__52245\ : std_logic;
signal \N__52244\ : std_logic;
signal \N__52243\ : std_logic;
signal \N__52242\ : std_logic;
signal \N__52241\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52239\ : std_logic;
signal \N__52238\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52236\ : std_logic;
signal \N__52235\ : std_logic;
signal \N__52234\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52232\ : std_logic;
signal \N__52231\ : std_logic;
signal \N__52230\ : std_logic;
signal \N__52229\ : std_logic;
signal \N__52228\ : std_logic;
signal \N__52227\ : std_logic;
signal \N__52226\ : std_logic;
signal \N__52225\ : std_logic;
signal \N__52224\ : std_logic;
signal \N__52223\ : std_logic;
signal \N__52222\ : std_logic;
signal \N__52221\ : std_logic;
signal \N__52220\ : std_logic;
signal \N__52219\ : std_logic;
signal \N__52218\ : std_logic;
signal \N__52217\ : std_logic;
signal \N__52216\ : std_logic;
signal \N__52215\ : std_logic;
signal \N__52214\ : std_logic;
signal \N__52213\ : std_logic;
signal \N__52212\ : std_logic;
signal \N__52211\ : std_logic;
signal \N__52210\ : std_logic;
signal \N__52209\ : std_logic;
signal \N__52208\ : std_logic;
signal \N__52207\ : std_logic;
signal \N__52206\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52204\ : std_logic;
signal \N__52203\ : std_logic;
signal \N__52202\ : std_logic;
signal \N__52201\ : std_logic;
signal \N__51902\ : std_logic;
signal \N__51899\ : std_logic;
signal \N__51896\ : std_logic;
signal \N__51895\ : std_logic;
signal \N__51894\ : std_logic;
signal \N__51891\ : std_logic;
signal \N__51890\ : std_logic;
signal \N__51889\ : std_logic;
signal \N__51886\ : std_logic;
signal \N__51883\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51879\ : std_logic;
signal \N__51876\ : std_logic;
signal \N__51873\ : std_logic;
signal \N__51872\ : std_logic;
signal \N__51869\ : std_logic;
signal \N__51866\ : std_logic;
signal \N__51863\ : std_logic;
signal \N__51858\ : std_logic;
signal \N__51855\ : std_logic;
signal \N__51852\ : std_logic;
signal \N__51849\ : std_logic;
signal \N__51844\ : std_logic;
signal \N__51841\ : std_logic;
signal \N__51836\ : std_logic;
signal \N__51827\ : std_logic;
signal \N__51826\ : std_logic;
signal \N__51825\ : std_logic;
signal \N__51824\ : std_logic;
signal \N__51823\ : std_logic;
signal \N__51822\ : std_logic;
signal \N__51821\ : std_logic;
signal \N__51820\ : std_logic;
signal \N__51819\ : std_logic;
signal \N__51818\ : std_logic;
signal \N__51817\ : std_logic;
signal \N__51816\ : std_logic;
signal \N__51815\ : std_logic;
signal \N__51814\ : std_logic;
signal \N__51813\ : std_logic;
signal \N__51812\ : std_logic;
signal \N__51811\ : std_logic;
signal \N__51810\ : std_logic;
signal \N__51809\ : std_logic;
signal \N__51808\ : std_logic;
signal \N__51807\ : std_logic;
signal \N__51806\ : std_logic;
signal \N__51805\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51803\ : std_logic;
signal \N__51802\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51799\ : std_logic;
signal \N__51798\ : std_logic;
signal \N__51797\ : std_logic;
signal \N__51796\ : std_logic;
signal \N__51795\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51793\ : std_logic;
signal \N__51792\ : std_logic;
signal \N__51791\ : std_logic;
signal \N__51790\ : std_logic;
signal \N__51789\ : std_logic;
signal \N__51788\ : std_logic;
signal \N__51787\ : std_logic;
signal \N__51786\ : std_logic;
signal \N__51785\ : std_logic;
signal \N__51784\ : std_logic;
signal \N__51783\ : std_logic;
signal \N__51782\ : std_logic;
signal \N__51781\ : std_logic;
signal \N__51780\ : std_logic;
signal \N__51779\ : std_logic;
signal \N__51778\ : std_logic;
signal \N__51777\ : std_logic;
signal \N__51776\ : std_logic;
signal \N__51775\ : std_logic;
signal \N__51774\ : std_logic;
signal \N__51773\ : std_logic;
signal \N__51772\ : std_logic;
signal \N__51771\ : std_logic;
signal \N__51770\ : std_logic;
signal \N__51769\ : std_logic;
signal \N__51768\ : std_logic;
signal \N__51767\ : std_logic;
signal \N__51766\ : std_logic;
signal \N__51765\ : std_logic;
signal \N__51764\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51761\ : std_logic;
signal \N__51760\ : std_logic;
signal \N__51759\ : std_logic;
signal \N__51758\ : std_logic;
signal \N__51757\ : std_logic;
signal \N__51756\ : std_logic;
signal \N__51755\ : std_logic;
signal \N__51754\ : std_logic;
signal \N__51753\ : std_logic;
signal \N__51752\ : std_logic;
signal \N__51751\ : std_logic;
signal \N__51750\ : std_logic;
signal \N__51749\ : std_logic;
signal \N__51748\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51746\ : std_logic;
signal \N__51745\ : std_logic;
signal \N__51744\ : std_logic;
signal \N__51743\ : std_logic;
signal \N__51742\ : std_logic;
signal \N__51741\ : std_logic;
signal \N__51740\ : std_logic;
signal \N__51739\ : std_logic;
signal \N__51738\ : std_logic;
signal \N__51737\ : std_logic;
signal \N__51736\ : std_logic;
signal \N__51735\ : std_logic;
signal \N__51734\ : std_logic;
signal \N__51733\ : std_logic;
signal \N__51732\ : std_logic;
signal \N__51731\ : std_logic;
signal \N__51730\ : std_logic;
signal \N__51729\ : std_logic;
signal \N__51728\ : std_logic;
signal \N__51727\ : std_logic;
signal \N__51726\ : std_logic;
signal \N__51725\ : std_logic;
signal \N__51724\ : std_logic;
signal \N__51723\ : std_logic;
signal \N__51722\ : std_logic;
signal \N__51721\ : std_logic;
signal \N__51720\ : std_logic;
signal \N__51719\ : std_logic;
signal \N__51718\ : std_logic;
signal \N__51717\ : std_logic;
signal \N__51716\ : std_logic;
signal \N__51715\ : std_logic;
signal \N__51714\ : std_logic;
signal \N__51713\ : std_logic;
signal \N__51712\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51710\ : std_logic;
signal \N__51709\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51707\ : std_logic;
signal \N__51706\ : std_logic;
signal \N__51705\ : std_logic;
signal \N__51704\ : std_logic;
signal \N__51703\ : std_logic;
signal \N__51702\ : std_logic;
signal \N__51701\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51699\ : std_logic;
signal \N__51698\ : std_logic;
signal \N__51697\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51695\ : std_logic;
signal \N__51694\ : std_logic;
signal \N__51693\ : std_logic;
signal \N__51692\ : std_logic;
signal \N__51691\ : std_logic;
signal \N__51690\ : std_logic;
signal \N__51689\ : std_logic;
signal \N__51688\ : std_logic;
signal \N__51687\ : std_logic;
signal \N__51686\ : std_logic;
signal \N__51685\ : std_logic;
signal \N__51684\ : std_logic;
signal \N__51683\ : std_logic;
signal \N__51682\ : std_logic;
signal \N__51681\ : std_logic;
signal \N__51680\ : std_logic;
signal \N__51679\ : std_logic;
signal \N__51678\ : std_logic;
signal \N__51677\ : std_logic;
signal \N__51676\ : std_logic;
signal \N__51675\ : std_logic;
signal \N__51674\ : std_logic;
signal \N__51673\ : std_logic;
signal \N__51672\ : std_logic;
signal \N__51671\ : std_logic;
signal \N__51670\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51668\ : std_logic;
signal \N__51667\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51665\ : std_logic;
signal \N__51664\ : std_logic;
signal \N__51663\ : std_logic;
signal \N__51662\ : std_logic;
signal \N__51661\ : std_logic;
signal \N__51660\ : std_logic;
signal \N__51659\ : std_logic;
signal \N__51658\ : std_logic;
signal \N__51657\ : std_logic;
signal \N__51656\ : std_logic;
signal \N__51655\ : std_logic;
signal \N__51654\ : std_logic;
signal \N__51653\ : std_logic;
signal \N__51652\ : std_logic;
signal \N__51651\ : std_logic;
signal \N__51650\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51648\ : std_logic;
signal \N__51647\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51644\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51269\ : std_logic;
signal \N__51266\ : std_logic;
signal \N__51263\ : std_logic;
signal \N__51262\ : std_logic;
signal \N__51259\ : std_logic;
signal \N__51256\ : std_logic;
signal \N__51253\ : std_logic;
signal \N__51248\ : std_logic;
signal \N__51245\ : std_logic;
signal \N__51242\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51238\ : std_logic;
signal \N__51235\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51227\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51223\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51217\ : std_logic;
signal \N__51216\ : std_logic;
signal \N__51215\ : std_logic;
signal \N__51214\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51208\ : std_logic;
signal \N__51205\ : std_logic;
signal \N__51198\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51192\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51188\ : std_logic;
signal \N__51185\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51179\ : std_logic;
signal \N__51178\ : std_logic;
signal \N__51175\ : std_logic;
signal \N__51172\ : std_logic;
signal \N__51169\ : std_logic;
signal \N__51166\ : std_logic;
signal \N__51163\ : std_logic;
signal \N__51158\ : std_logic;
signal \N__51151\ : std_logic;
signal \N__51146\ : std_logic;
signal \N__51145\ : std_logic;
signal \N__51144\ : std_logic;
signal \N__51143\ : std_logic;
signal \N__51138\ : std_logic;
signal \N__51133\ : std_logic;
signal \N__51128\ : std_logic;
signal \N__51125\ : std_logic;
signal \N__51124\ : std_logic;
signal \N__51121\ : std_logic;
signal \N__51118\ : std_logic;
signal \N__51113\ : std_logic;
signal \N__51110\ : std_logic;
signal \N__51107\ : std_logic;
signal \N__51104\ : std_logic;
signal \N__51101\ : std_logic;
signal \N__51100\ : std_logic;
signal \N__51097\ : std_logic;
signal \N__51094\ : std_logic;
signal \N__51089\ : std_logic;
signal \N__51086\ : std_logic;
signal \N__51083\ : std_logic;
signal \N__51080\ : std_logic;
signal \N__51077\ : std_logic;
signal \N__51076\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51074\ : std_logic;
signal \N__51071\ : std_logic;
signal \N__51070\ : std_logic;
signal \N__51069\ : std_logic;
signal \N__51068\ : std_logic;
signal \N__51065\ : std_logic;
signal \N__51064\ : std_logic;
signal \N__51063\ : std_logic;
signal \N__51062\ : std_logic;
signal \N__51059\ : std_logic;
signal \N__51056\ : std_logic;
signal \N__51055\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51053\ : std_logic;
signal \N__51052\ : std_logic;
signal \N__51051\ : std_logic;
signal \N__51050\ : std_logic;
signal \N__51047\ : std_logic;
signal \N__51044\ : std_logic;
signal \N__51043\ : std_logic;
signal \N__51042\ : std_logic;
signal \N__51041\ : std_logic;
signal \N__51040\ : std_logic;
signal \N__51039\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51037\ : std_logic;
signal \N__51034\ : std_logic;
signal \N__51031\ : std_logic;
signal \N__51030\ : std_logic;
signal \N__51029\ : std_logic;
signal \N__51026\ : std_logic;
signal \N__51023\ : std_logic;
signal \N__51020\ : std_logic;
signal \N__51019\ : std_logic;
signal \N__51018\ : std_logic;
signal \N__51017\ : std_logic;
signal \N__51014\ : std_logic;
signal \N__51009\ : std_logic;
signal \N__51006\ : std_logic;
signal \N__51003\ : std_logic;
signal \N__51000\ : std_logic;
signal \N__50997\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50991\ : std_logic;
signal \N__50986\ : std_logic;
signal \N__50985\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50983\ : std_logic;
signal \N__50982\ : std_logic;
signal \N__50979\ : std_logic;
signal \N__50976\ : std_logic;
signal \N__50973\ : std_logic;
signal \N__50970\ : std_logic;
signal \N__50967\ : std_logic;
signal \N__50964\ : std_logic;
signal \N__50961\ : std_logic;
signal \N__50956\ : std_logic;
signal \N__50953\ : std_logic;
signal \N__50950\ : std_logic;
signal \N__50943\ : std_logic;
signal \N__50940\ : std_logic;
signal \N__50939\ : std_logic;
signal \N__50938\ : std_logic;
signal \N__50935\ : std_logic;
signal \N__50932\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50930\ : std_logic;
signal \N__50929\ : std_logic;
signal \N__50928\ : std_logic;
signal \N__50925\ : std_logic;
signal \N__50914\ : std_logic;
signal \N__50907\ : std_logic;
signal \N__50904\ : std_logic;
signal \N__50903\ : std_logic;
signal \N__50900\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50898\ : std_logic;
signal \N__50897\ : std_logic;
signal \N__50896\ : std_logic;
signal \N__50893\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50889\ : std_logic;
signal \N__50884\ : std_logic;
signal \N__50883\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50881\ : std_logic;
signal \N__50880\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50878\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50861\ : std_logic;
signal \N__50858\ : std_logic;
signal \N__50855\ : std_logic;
signal \N__50852\ : std_logic;
signal \N__50851\ : std_logic;
signal \N__50848\ : std_logic;
signal \N__50845\ : std_logic;
signal \N__50840\ : std_logic;
signal \N__50837\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50831\ : std_logic;
signal \N__50828\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50816\ : std_logic;
signal \N__50815\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50811\ : std_logic;
signal \N__50808\ : std_logic;
signal \N__50805\ : std_logic;
signal \N__50802\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50787\ : std_logic;
signal \N__50784\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50769\ : std_logic;
signal \N__50766\ : std_logic;
signal \N__50763\ : std_logic;
signal \N__50758\ : std_logic;
signal \N__50755\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50747\ : std_logic;
signal \N__50742\ : std_logic;
signal \N__50739\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50719\ : std_logic;
signal \N__50718\ : std_logic;
signal \N__50717\ : std_logic;
signal \N__50716\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50707\ : std_logic;
signal \N__50696\ : std_logic;
signal \N__50689\ : std_logic;
signal \N__50682\ : std_logic;
signal \N__50667\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50655\ : std_logic;
signal \N__50652\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50646\ : std_logic;
signal \N__50643\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50629\ : std_logic;
signal \N__50624\ : std_logic;
signal \N__50609\ : std_logic;
signal \N__50606\ : std_logic;
signal \N__50603\ : std_logic;
signal \N__50600\ : std_logic;
signal \N__50597\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50593\ : std_logic;
signal \N__50590\ : std_logic;
signal \N__50587\ : std_logic;
signal \N__50584\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50570\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50564\ : std_logic;
signal \N__50561\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50545\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50542\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50531\ : std_logic;
signal \N__50530\ : std_logic;
signal \N__50529\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50508\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50492\ : std_logic;
signal \N__50489\ : std_logic;
signal \N__50488\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50483\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50468\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50452\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50440\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50420\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50382\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50374\ : std_logic;
signal \N__50367\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50346\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50331\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50328\ : std_logic;
signal \N__50327\ : std_logic;
signal \N__50324\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50280\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50229\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50225\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50221\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50209\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50196\ : std_logic;
signal \N__50189\ : std_logic;
signal \N__50186\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50180\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50168\ : std_logic;
signal \N__50161\ : std_logic;
signal \N__50156\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50144\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50117\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50111\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50072\ : std_logic;
signal \N__50069\ : std_logic;
signal \N__50066\ : std_logic;
signal \N__50063\ : std_logic;
signal \N__50062\ : std_logic;
signal \N__50061\ : std_logic;
signal \N__50060\ : std_logic;
signal \N__50059\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50057\ : std_logic;
signal \N__50056\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50054\ : std_logic;
signal \N__50053\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50051\ : std_logic;
signal \N__50050\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50041\ : std_logic;
signal \N__50038\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50036\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50032\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50030\ : std_logic;
signal \N__50029\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50027\ : std_logic;
signal \N__50024\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50020\ : std_logic;
signal \N__50017\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49997\ : std_logic;
signal \N__49996\ : std_logic;
signal \N__49995\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49991\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49961\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49926\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49912\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49892\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49877\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49823\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49813\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49793\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49789\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49760\ : std_logic;
signal \N__49757\ : std_logic;
signal \N__49754\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49740\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49731\ : std_logic;
signal \N__49728\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49710\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49681\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49673\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49662\ : std_logic;
signal \N__49659\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49655\ : std_logic;
signal \N__49654\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49648\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49613\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49603\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49583\ : std_logic;
signal \N__49580\ : std_logic;
signal \N__49577\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49565\ : std_logic;
signal \N__49562\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49550\ : std_logic;
signal \N__49547\ : std_logic;
signal \N__49544\ : std_logic;
signal \N__49541\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49532\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49529\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49519\ : std_logic;
signal \N__49510\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49484\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49440\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49430\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49400\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49391\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49364\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49355\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49349\ : std_logic;
signal \N__49338\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49315\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49307\ : std_logic;
signal \N__49306\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49303\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49299\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49291\ : std_logic;
signal \N__49290\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49283\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49275\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49261\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49250\ : std_logic;
signal \N__49247\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49241\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49217\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49193\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49161\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49149\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49142\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49085\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49073\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49053\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49027\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48960\ : std_logic;
signal \N__48957\ : std_logic;
signal \N__48956\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48952\ : std_logic;
signal \N__48951\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48930\ : std_logic;
signal \N__48929\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48912\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48909\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48903\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48899\ : std_logic;
signal \N__48898\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48889\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48850\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48796\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48771\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48692\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48666\ : std_logic;
signal \N__48665\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48636\ : std_logic;
signal \N__48633\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48618\ : std_logic;
signal \N__48615\ : std_logic;
signal \N__48612\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48601\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48568\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48553\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48522\ : std_logic;
signal \N__48515\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48499\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48491\ : std_logic;
signal \N__48490\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48488\ : std_logic;
signal \N__48487\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48485\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48476\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48473\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48471\ : std_logic;
signal \N__48470\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48467\ : std_logic;
signal \N__48466\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48455\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48452\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48446\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48347\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48294\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48116\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48094\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48062\ : std_logic;
signal \N__48059\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48052\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48041\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48015\ : std_logic;
signal \N__48012\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47977\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47965\ : std_logic;
signal \N__47962\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47951\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47936\ : std_logic;
signal \N__47933\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47929\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47903\ : std_logic;
signal \N__47900\ : std_logic;
signal \N__47897\ : std_logic;
signal \N__47894\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47717\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47660\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47621\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47588\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47582\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47525\ : std_logic;
signal \N__47522\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47503\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47500\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47497\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47374\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47352\ : std_logic;
signal \N__47349\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47346\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47329\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47251\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47210\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47171\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47104\ : std_logic;
signal \N__47101\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46844\ : std_logic;
signal \N__46841\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46780\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46774\ : std_logic;
signal \N__46771\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46753\ : std_logic;
signal \N__46752\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46738\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46518\ : std_logic;
signal \N__46515\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46430\ : std_logic;
signal \N__46427\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46421\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46394\ : std_logic;
signal \N__46391\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46356\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46352\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46288\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46233\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46144\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46141\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46130\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46075\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45980\ : std_logic;
signal \N__45979\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45956\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45918\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45776\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45748\ : std_logic;
signal \N__45745\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45601\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45577\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45574\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45532\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45413\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45351\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45320\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45308\ : std_logic;
signal \N__45301\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45118\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45115\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45103\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45100\ : std_logic;
signal \N__45097\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45068\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45002\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44951\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44939\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44924\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44876\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44861\ : std_logic;
signal \N__44858\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44803\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44672\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44600\ : std_logic;
signal \N__44597\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44576\ : std_logic;
signal \N__44573\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44519\ : std_logic;
signal \N__44516\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44501\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44462\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44438\ : std_logic;
signal \N__44435\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44429\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44396\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44381\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44366\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44342\ : std_logic;
signal \N__44339\ : std_logic;
signal \N__44336\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44318\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44309\ : std_logic;
signal \N__44306\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44291\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44264\ : std_logic;
signal \N__44261\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44249\ : std_logic;
signal \N__44246\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44117\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44023\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43999\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43993\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43952\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43949\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43889\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43871\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43756\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43618\ : std_logic;
signal \N__43615\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43535\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43355\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43252\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43244\ : std_logic;
signal \N__43241\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43184\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43172\ : std_logic;
signal \N__43169\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43112\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43049\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43036\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43022\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42926\ : std_logic;
signal \N__42923\ : std_logic;
signal \N__42920\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42911\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42899\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42854\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42827\ : std_logic;
signal \N__42824\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42776\ : std_logic;
signal \N__42773\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42679\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42659\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42633\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42557\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42553\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42433\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42422\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42281\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42211\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42170\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42167\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42158\ : std_logic;
signal \N__42157\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42146\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42142\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42067\ : std_logic;
signal \N__42064\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42014\ : std_logic;
signal \N__42013\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41983\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41911\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41893\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41884\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41608\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41605\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41572\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41291\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41240\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41195\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41051\ : std_logic;
signal \N__41048\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41033\ : std_logic;
signal \N__41030\ : std_logic;
signal \N__41027\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40978\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40931\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40904\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40877\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40646\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40624\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40592\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40537\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40429\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40385\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40357\ : std_logic;
signal \N__40354\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40297\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40295\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40286\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40255\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40180\ : std_logic;
signal \N__40177\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40006\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39920\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39899\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39772\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39749\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39638\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39602\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39559\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39194\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39098\ : std_logic;
signal \N__39095\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39071\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38990\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38963\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38872\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38863\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38717\ : std_logic;
signal \N__38714\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38705\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38684\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38663\ : std_logic;
signal \N__38660\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38521\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38246\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38144\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38126\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37673\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37505\ : std_logic;
signal \N__37502\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37420\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37348\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37334\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37268\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37202\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37175\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36668\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36578\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36350\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35690\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35486\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35216\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34868\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34196\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33866\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33745\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33398\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26062\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal cs_rpi2flash_c : std_logic;
signal clk_c : std_logic;
signal \pll128M2_inst.pll_clk64_0\ : std_logic;
signal \pll128M2_inst.pll_clk128\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \sRAM_pointer_write_cry_0\ : std_logic;
signal \sRAM_pointer_write_cry_1\ : std_logic;
signal \sRAM_pointer_write_cry_2\ : std_logic;
signal \sRAM_pointer_write_cry_3\ : std_logic;
signal \sRAM_pointer_write_cry_4\ : std_logic;
signal \sRAM_pointer_write_cry_5\ : std_logic;
signal \sRAM_pointer_write_cry_6\ : std_logic;
signal \sRAM_pointer_write_cry_7\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \sRAM_pointer_write_cry_8\ : std_logic;
signal \sRAM_pointer_write_cry_9\ : std_logic;
signal \sRAM_pointer_write_cry_10\ : std_logic;
signal \sRAM_pointer_write_cry_11\ : std_logic;
signal \sRAM_pointer_write_cry_12\ : std_logic;
signal \sRAM_pointer_write_cry_13\ : std_logic;
signal \sRAM_pointer_write_cry_14\ : std_logic;
signal \sRAM_pointer_write_cry_15\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \sRAM_pointer_write_cry_16\ : std_logic;
signal \sRAM_pointer_write_cry_17\ : std_logic;
signal \N_1487_g\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_1531_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1\ : std_logic;
signal button_mode_c : std_logic;
signal \button_mode_ibuf_RNIN5KZ0Z7\ : std_logic;
signal \DAC_cs_c\ : std_logic;
signal \bfn_3_6_0_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_s_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_s_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0\ : std_logic;
signal \bfn_3_8_0_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_6\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_1531\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_start_iZ0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_start_i_i\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_48_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_36\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_150_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_48\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1414_cascade_\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1415_cascade_\ : std_logic;
signal \DAC_mosi_c\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1421_cascade_\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1422\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6\ : std_logic;
signal \DAC_sclk_c\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_1737\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_1737_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_1540\ : std_logic;
signal \spi_master_inst.ss_start_i\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1411\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1418\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6\ : std_logic;
signal \spi_master_inst.o_sclk_RNIH6AC\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3\ : std_logic;
signal \spi_mosi_ready64_prevZ0Z2\ : std_logic;
signal \spi_mosi_ready64_prevZ0\ : std_logic;
signal \spi_mosi_ready64_prevZ0Z3\ : std_logic;
signal \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_\ : std_logic;
signal \bfn_6_12_0_\ : std_logic;
signal \sEETrigCounterZ0Z_1\ : std_logic;
signal un8_trig_prev_0_cry_0 : std_logic;
signal \sEETrigCounterZ0Z_2\ : std_logic;
signal un8_trig_prev_0_cry_1 : std_logic;
signal \sEETrigCounterZ0Z_3\ : std_logic;
signal un8_trig_prev_0_cry_2 : std_logic;
signal \sEETrigCounterZ0Z_4\ : std_logic;
signal un8_trig_prev_0_cry_3 : std_logic;
signal \sEETrigCounterZ0Z_5\ : std_logic;
signal un8_trig_prev_0_cry_4 : std_logic;
signal \sEETrigCounterZ0Z_6\ : std_logic;
signal un8_trig_prev_0_cry_5 : std_logic;
signal \sEETrigCounterZ0Z_7\ : std_logic;
signal un8_trig_prev_0_cry_6 : std_logic;
signal un8_trig_prev_0_cry_7 : std_logic;
signal \bfn_6_13_0_\ : std_logic;
signal un8_trig_prev_0_cry_8 : std_logic;
signal un8_trig_prev_0_cry_9 : std_logic;
signal un8_trig_prev_0_cry_10 : std_logic;
signal un8_trig_prev_0_cry_11 : std_logic;
signal un8_trig_prev_0_cry_12 : std_logic;
signal un8_trig_prev_0_cry_13 : std_logic;
signal un8_trig_prev_0_cry_14 : std_logic;
signal \sEETrigCounterZ0Z_10\ : std_logic;
signal \sEETrigCounterZ0Z_11\ : std_logic;
signal \sEETrigCounterZ0Z_12\ : std_logic;
signal \sEETrigCounterZ0Z_13\ : std_logic;
signal \sEETrigCounterZ0Z_14\ : std_logic;
signal \sEETrigCounterZ0Z_15\ : std_logic;
signal \sEETrigCounterZ0Z_8\ : std_logic;
signal \sEETrigCounterZ0Z_9\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_6\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_5\ : std_logic;
signal \N_316_cascade_\ : std_logic;
signal \N_317_cascade_\ : std_logic;
signal \sAddress_RNI8U0V1Z0Z_1_cascade_\ : std_logic;
signal \sAddress_RNI8U0V1Z0Z_1\ : std_logic;
signal \N_454_cascade_\ : std_logic;
signal \N_346_i_cascade_\ : std_logic;
signal \un1_spointer11_8_0_0_a2_1_cascade_\ : std_logic;
signal \sAddress_RNI7G5E2Z0Z_6\ : std_logic;
signal \sAddressZ0Z_7\ : std_logic;
signal \sAddressZ0Z_6\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5\ : std_logic;
signal \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\ : std_logic;
signal spi_mosi_ready : std_logic;
signal \spi_mosi_ready_prevZ0\ : std_logic;
signal \spi_mosi_ready_prevZ0Z2\ : std_logic;
signal \spi_mosi_ready_prevZ0Z3\ : std_logic;
signal un8_trig_prev_0 : std_logic;
signal un10_trig_prev_0 : std_logic;
signal \sTrigCounter_i_0\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal un10_trig_prev_1 : std_logic;
signal \sTrigCounter_i_1\ : std_logic;
signal un10_trig_prev_cry_0 : std_logic;
signal un10_trig_prev_2 : std_logic;
signal \sTrigCounter_i_2\ : std_logic;
signal un10_trig_prev_cry_1 : std_logic;
signal un10_trig_prev_3 : std_logic;
signal \sTrigCounter_i_3\ : std_logic;
signal un10_trig_prev_cry_2 : std_logic;
signal un10_trig_prev_4 : std_logic;
signal \sTrigCounter_i_4\ : std_logic;
signal un10_trig_prev_cry_3 : std_logic;
signal un10_trig_prev_5 : std_logic;
signal \sTrigCounter_i_5\ : std_logic;
signal un10_trig_prev_cry_4 : std_logic;
signal un10_trig_prev_6 : std_logic;
signal \sTrigCounter_i_6\ : std_logic;
signal un10_trig_prev_cry_5 : std_logic;
signal un10_trig_prev_7 : std_logic;
signal \sTrigCounter_i_7\ : std_logic;
signal un10_trig_prev_cry_6 : std_logic;
signal un10_trig_prev_cry_7 : std_logic;
signal un10_trig_prev_8 : std_logic;
signal \sTrigCounter_i_8\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal un10_trig_prev_9 : std_logic;
signal \sTrigCounter_i_9\ : std_logic;
signal un10_trig_prev_cry_8 : std_logic;
signal un10_trig_prev_10 : std_logic;
signal \sTrigCounter_i_10\ : std_logic;
signal un10_trig_prev_cry_9 : std_logic;
signal un10_trig_prev_11 : std_logic;
signal \sTrigCounter_i_11\ : std_logic;
signal un10_trig_prev_cry_10 : std_logic;
signal un10_trig_prev_12 : std_logic;
signal \sTrigCounter_i_12\ : std_logic;
signal un10_trig_prev_cry_11 : std_logic;
signal un10_trig_prev_13 : std_logic;
signal \sTrigCounter_i_13\ : std_logic;
signal un10_trig_prev_cry_12 : std_logic;
signal un10_trig_prev_14 : std_logic;
signal \sTrigCounter_i_14\ : std_logic;
signal un10_trig_prev_cry_13 : std_logic;
signal un10_trig_prev_15 : std_logic;
signal \sTrigCounter_i_15\ : std_logic;
signal un10_trig_prev_cry_14 : std_logic;
signal un10_trig_prev_cry_15 : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \N_173\ : std_logic;
signal \INVspi_slave_inst.rx_done_neg_sclk_iC_net\ : std_logic;
signal \sEEADC_freqZ0Z_4\ : std_logic;
signal un3_trig_0 : std_logic;
signal \sEEADC_freqZ0Z_5\ : std_logic;
signal spi_mosi_rpi_c : std_logic;
signal spi_mosi_ft_c : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7\ : std_logic;
signal \sDAC_mem_11_1_sqmuxa\ : std_logic;
signal \N_344_cascade_\ : std_logic;
signal \sDAC_mem_35_1_sqmuxa\ : std_logic;
signal \sEESingleCont_RNOZ0Z_0\ : std_logic;
signal \sEESingleContZ0\ : std_logic;
signal \N_1631\ : std_logic;
signal \sEETrigInternal_3_iv_0_0_i_0\ : std_logic;
signal \spi_slave_inst.rx_done_neg_sclk_iZ0\ : std_logic;
signal \spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541\ : std_logic;
signal \spi_slave_inst.rx_done_reg1_iZ0\ : std_logic;
signal \N_319_cascade_\ : std_logic;
signal \sAddress_RNI9IH12_2Z0Z_1\ : std_logic;
signal \spi_slave_inst.rx_done_reg2_iZ0\ : std_logic;
signal \spi_slave_inst.rx_done_reg3_iZ0\ : std_logic;
signal \spi_slave_inst.rx_ready_i_RNOZ0Z_0\ : std_logic;
signal \sPointer_RNI5LBD1Z0Z_0_cascade_\ : std_logic;
signal \sDAC_mem_17_1_sqmuxa_0_a2_0_a2_1_0\ : std_logic;
signal \sAddressZ0Z_4\ : std_logic;
signal \sAddress_RNIP2UK1Z0Z_4_cascade_\ : std_logic;
signal trig_rpi_c : std_logic;
signal trig_ext_c : std_logic;
signal trig_ft_c : std_logic;
signal \trig_prevZ0\ : std_logic;
signal \g3_0_cascade_\ : std_logic;
signal \sAddress_RNI70I7Z0Z_1_cascade_\ : std_logic;
signal g1_i_a4_0_0 : std_logic;
signal \N_8_mux\ : std_logic;
signal \un10_trig_prev_cry_15_THRU_CO\ : std_logic;
signal \N_178\ : std_logic;
signal un1_scounter_i_0 : std_logic;
signal \N_178_cascade_\ : std_logic;
signal \N_96\ : std_logic;
signal \N_77_cascade_\ : std_logic;
signal \sPeriod_prevZ0\ : std_logic;
signal un1_reset_rpi_inv_2_0 : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \un1_sTrigCounter_cry_0\ : std_logic;
signal \sTrigCounterZ0Z_2\ : std_logic;
signal \un1_sTrigCounter_cry_1\ : std_logic;
signal \sTrigCounterZ0Z_3\ : std_logic;
signal \un1_sTrigCounter_cry_2\ : std_logic;
signal \sTrigCounterZ0Z_4\ : std_logic;
signal \un1_sTrigCounter_cry_3\ : std_logic;
signal \sTrigCounterZ0Z_5\ : std_logic;
signal \un1_sTrigCounter_cry_4\ : std_logic;
signal \sTrigCounterZ0Z_6\ : std_logic;
signal \un1_sTrigCounter_cry_5\ : std_logic;
signal \sTrigCounterZ0Z_7\ : std_logic;
signal \un1_sTrigCounter_cry_6\ : std_logic;
signal \un1_sTrigCounter_cry_7\ : std_logic;
signal \sTrigCounterZ0Z_8\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \sTrigCounterZ0Z_9\ : std_logic;
signal \un1_sTrigCounter_cry_8\ : std_logic;
signal \sTrigCounterZ0Z_10\ : std_logic;
signal \un1_sTrigCounter_cry_9\ : std_logic;
signal \sTrigCounterZ0Z_11\ : std_logic;
signal \un1_sTrigCounter_cry_10\ : std_logic;
signal \sTrigCounterZ0Z_12\ : std_logic;
signal \un1_sTrigCounter_cry_11\ : std_logic;
signal \sTrigCounterZ0Z_13\ : std_logic;
signal \un1_sTrigCounter_cry_12\ : std_logic;
signal \sTrigCounterZ0Z_14\ : std_logic;
signal \un1_sTrigCounter_cry_13\ : std_logic;
signal \un1_sTrigCounter_cry_14\ : std_logic;
signal \sTrigCounterZ0Z_15\ : std_logic;
signal \N_82_i\ : std_logic;
signal \sDAC_mem_29_1_sqmuxa\ : std_logic;
signal \sEEPon_1_sqmuxa\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10\ : std_logic;
signal \sDAC_mem_38_1_sqmuxa\ : std_logic;
signal \sAddress_RNI6VH7_3Z0Z_1\ : std_logic;
signal \sAddress_RNI6VH7_3Z0Z_1_cascade_\ : std_logic;
signal \sDAC_mem_10_1_sqmuxa\ : std_logic;
signal \N_326_cascade_\ : std_logic;
signal \LED_ACQ_obuf_RNOZ0\ : std_logic;
signal \sAddress_RNIAM2A_0Z0Z_1_cascade_\ : std_logic;
signal \N_445_cascade_\ : std_logic;
signal \sAddress_RNI6VH7_5Z0Z_1\ : std_logic;
signal \N_445\ : std_logic;
signal \N_316\ : std_logic;
signal un1_spointer11_0 : std_logic;
signal \sAddress_RNI6VH7_2Z0Z_1\ : std_logic;
signal \sEETrigInternalZ0\ : std_logic;
signal g3_0 : std_logic;
signal \sEETrigInternal_prevZ0\ : std_logic;
signal \LED_MODE_c\ : std_logic;
signal \N_831_16_cascade_\ : std_logic;
signal \N_319\ : std_logic;
signal \g0_13_cascade_\ : std_logic;
signal g0_1_0 : std_logic;
signal g0_15_0 : std_logic;
signal g0_13_1 : std_logic;
signal g0_17_0 : std_logic;
signal \N_326\ : std_logic;
signal g0_16_0 : std_logic;
signal g1_i_a4_6 : std_logic;
signal \g1_i_a4_5_cascade_\ : std_logic;
signal un1_reset_rpi_inv_2_0_o2_5 : std_logic;
signal \g1_i_a4_9_cascade_\ : std_logic;
signal \sEETrigInternal_prev_RNIH3OJZ0Z1\ : std_logic;
signal g0_0_1 : std_logic;
signal g0_16 : std_logic;
signal g0_11 : std_logic;
signal g0_14 : std_logic;
signal \sDAC_mem_30_1_sqmuxa\ : std_logic;
signal \sEEPonZ0Z_0\ : std_logic;
signal \sEEPon_i_0\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \sEEPonZ0Z_1\ : std_logic;
signal \sEEPon_i_1\ : std_logic;
signal un7_spon_cry_0 : std_logic;
signal \sEEPonZ0Z_2\ : std_logic;
signal \sEEPon_i_2\ : std_logic;
signal un7_spon_cry_1 : std_logic;
signal \sEEPonZ0Z_3\ : std_logic;
signal \sEEPon_i_3\ : std_logic;
signal un7_spon_cry_2 : std_logic;
signal \sEEPonZ0Z_4\ : std_logic;
signal \sEEPon_i_4\ : std_logic;
signal un7_spon_cry_3 : std_logic;
signal \sEEPonZ0Z_5\ : std_logic;
signal \sEEPon_i_5\ : std_logic;
signal un7_spon_cry_4 : std_logic;
signal \sEEPonZ0Z_6\ : std_logic;
signal \sEEPon_i_6\ : std_logic;
signal un7_spon_cry_5 : std_logic;
signal \sEEPonZ0Z_7\ : std_logic;
signal \sEEPon_i_7\ : std_logic;
signal un7_spon_cry_6 : std_logic;
signal un7_spon_cry_7 : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal un7_spon_cry_8 : std_logic;
signal un7_spon_cry_9 : std_logic;
signal un7_spon_cry_10 : std_logic;
signal un7_spon_cry_11 : std_logic;
signal un7_spon_cry_12 : std_logic;
signal un7_spon_cry_13 : std_logic;
signal un7_spon_cry_14 : std_logic;
signal un7_spon_cry_15 : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal un7_spon_cry_16 : std_logic;
signal un7_spon_cry_17 : std_logic;
signal un7_spon_cry_18 : std_logic;
signal un7_spon_cry_19 : std_logic;
signal un7_spon_cry_20 : std_logic;
signal un7_spon_cry_21 : std_logic;
signal un7_spon_cry_22 : std_logic;
signal un7_spon_cry_23 : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \pon_obuf_RNOZ0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_1\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_10\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_11\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_13\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_14\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_15\ : std_logic;
signal \sDAC_mem_42_1_sqmuxa\ : std_logic;
signal \sDAC_mem_14_1_sqmuxa\ : std_logic;
signal \sAddress_RNI9IH12Z0Z_0\ : std_logic;
signal \sAddress_RNI9IH12_1Z0Z_2\ : std_logic;
signal \sDAC_mem_15_1_sqmuxa\ : std_logic;
signal un21_trig_prev_21_5 : std_logic;
signal \op_gt_op_gt_un13_striginternallto23_5_cascade_\ : std_logic;
signal un1_reset_rpi_inv_2_0_o2_2 : std_logic;
signal g0_13_0 : std_logic;
signal un21_trig_prev_21_4 : std_logic;
signal g0_6 : std_logic;
signal \N_99\ : std_logic;
signal op_gt_op_gt_un13_striginternallto23_3 : std_logic;
signal \N_831_16\ : std_logic;
signal op_gt_op_gt_un13_striginternallto23_6 : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_158_7\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spi_start_iZ0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_158_7_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0\ : std_logic;
signal g2_6 : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_i6_3\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_i6\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_3\ : std_logic;
signal \spi_slave_inst.un23_i_ssn_3_cascade_\ : std_logic;
signal \spi_slave_inst.un23_i_ssn_cascade_\ : std_logic;
signal g0_10 : std_logic;
signal g0_10_0 : std_logic;
signal \sDAC_mem_31_1_sqmuxa\ : std_logic;
signal \sAddress_RNIA6242_4Z0Z_0\ : std_logic;
signal \sAddress_RNIA6242Z0Z_0\ : std_logic;
signal \LED3_c_i\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15\ : std_logic;
signal \sDAC_dataZ0Z_0\ : std_logic;
signal \sDAC_dataZ0Z_1\ : std_logic;
signal \sDAC_dataZ0Z_11\ : std_logic;
signal \sDAC_dataZ0Z_12\ : std_logic;
signal \sDAC_dataZ0Z_13\ : std_logic;
signal \sDAC_dataZ0Z_14\ : std_logic;
signal \sDAC_dataZ0Z_15\ : std_logic;
signal \sAddress_RNIETI62Z0Z_1\ : std_logic;
signal \sEEPeriodZ0Z_0\ : std_logic;
signal \sEEPeriod_i_0\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \sEEPeriodZ0Z_1\ : std_logic;
signal \sEEPeriod_i_1\ : std_logic;
signal un4_speriod_cry_0 : std_logic;
signal \sEEPeriodZ0Z_2\ : std_logic;
signal \sEEPeriod_i_2\ : std_logic;
signal un4_speriod_cry_1 : std_logic;
signal \sEEPeriodZ0Z_3\ : std_logic;
signal \sEEPeriod_i_3\ : std_logic;
signal un4_speriod_cry_2 : std_logic;
signal \sEEPeriodZ0Z_4\ : std_logic;
signal \sEEPeriod_i_4\ : std_logic;
signal un4_speriod_cry_3 : std_logic;
signal \sEEPeriodZ0Z_5\ : std_logic;
signal \sEEPeriod_i_5\ : std_logic;
signal un4_speriod_cry_4 : std_logic;
signal \sEEPeriodZ0Z_6\ : std_logic;
signal \sEEPeriod_i_6\ : std_logic;
signal un4_speriod_cry_5 : std_logic;
signal \sEEPeriodZ0Z_7\ : std_logic;
signal \sEEPeriod_i_7\ : std_logic;
signal un4_speriod_cry_6 : std_logic;
signal un4_speriod_cry_7 : std_logic;
signal \sEEPeriodZ0Z_8\ : std_logic;
signal \sEEPeriod_i_8\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \sEEPeriodZ0Z_9\ : std_logic;
signal \sEEPeriod_i_9\ : std_logic;
signal un4_speriod_cry_8 : std_logic;
signal \sEEPeriodZ0Z_10\ : std_logic;
signal \sEEPeriod_i_10\ : std_logic;
signal un4_speriod_cry_9 : std_logic;
signal \sEEPeriodZ0Z_11\ : std_logic;
signal \sEEPeriod_i_11\ : std_logic;
signal un4_speriod_cry_10 : std_logic;
signal \sEEPeriodZ0Z_12\ : std_logic;
signal \sEEPeriod_i_12\ : std_logic;
signal un4_speriod_cry_11 : std_logic;
signal \sEEPeriodZ0Z_13\ : std_logic;
signal \sEEPeriod_i_13\ : std_logic;
signal un4_speriod_cry_12 : std_logic;
signal \sEEPeriodZ0Z_14\ : std_logic;
signal \sEEPeriod_i_14\ : std_logic;
signal un4_speriod_cry_13 : std_logic;
signal \sEEPeriodZ0Z_15\ : std_logic;
signal \sEEPeriod_i_15\ : std_logic;
signal un4_speriod_cry_14 : std_logic;
signal un4_speriod_cry_15 : std_logic;
signal \sEEPeriodZ0Z_16\ : std_logic;
signal \sEEPeriod_i_16\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \sEEPeriodZ0Z_17\ : std_logic;
signal \sEEPeriod_i_17\ : std_logic;
signal un4_speriod_cry_16 : std_logic;
signal \sEEPeriodZ0Z_18\ : std_logic;
signal \sEEPeriod_i_18\ : std_logic;
signal un4_speriod_cry_17 : std_logic;
signal \sEEPeriodZ0Z_19\ : std_logic;
signal \sEEPeriod_i_19\ : std_logic;
signal un4_speriod_cry_18 : std_logic;
signal \sEEPeriodZ0Z_20\ : std_logic;
signal \sEEPeriod_i_20\ : std_logic;
signal un4_speriod_cry_19 : std_logic;
signal \sEEPeriodZ0Z_21\ : std_logic;
signal \sEEPeriod_i_21\ : std_logic;
signal un4_speriod_cry_20 : std_logic;
signal \sEEPeriodZ0Z_22\ : std_logic;
signal \sEEPeriod_i_22\ : std_logic;
signal un4_speriod_cry_21 : std_logic;
signal \sEEPeriodZ0Z_23\ : std_logic;
signal \sEEPeriod_i_23\ : std_logic;
signal un4_speriod_cry_22 : std_logic;
signal un4_speriod_cry_23 : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal un1_spointer11_2_0_0_a2_6 : std_logic;
signal un1_spointer11_2_0_0_a2_1 : std_logic;
signal \sTrigInternalZ0\ : std_logic;
signal op_gt_op_gt_un13_striginternal_0 : std_logic;
signal \un4_speriod_cry_23_THRU_CO\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \sCounter_cry_0\ : std_logic;
signal \sCounter_cry_1\ : std_logic;
signal \sCounter_cry_2\ : std_logic;
signal \sCounter_cry_3\ : std_logic;
signal \sCounter_cry_4\ : std_logic;
signal \sCounter_cry_5\ : std_logic;
signal \sCounter_cry_6\ : std_logic;
signal \sCounter_cry_7\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \sCounter_cry_8\ : std_logic;
signal \sCounter_cry_9\ : std_logic;
signal \sCounter_cry_10\ : std_logic;
signal \sCounter_cry_11\ : std_logic;
signal \sCounter_cry_12\ : std_logic;
signal \sCounter_cry_13\ : std_logic;
signal \sCounter_cry_14\ : std_logic;
signal \sCounter_cry_15\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \sCounter_cry_16\ : std_logic;
signal \sCounter_cry_17\ : std_logic;
signal \sCounter_cry_18\ : std_logic;
signal \sCounter_cry_19\ : std_logic;
signal \sCounter_cry_20\ : std_logic;
signal \sCounter_cry_21\ : std_logic;
signal \LED_ACQ_c_i\ : std_logic;
signal \sCounter_cry_22\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7\ : std_logic;
signal un1_spointer11_5_0_2 : std_logic;
signal \sAddress_RNIA6242_3Z0Z_0\ : std_logic;
signal \sEEDelayACQZ0Z_0\ : std_logic;
signal \sEEDelayACQ_i_0\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \sEEDelayACQZ0Z_1\ : std_logic;
signal \sEEDelayACQ_i_1\ : std_logic;
signal un4_sacqtime_cry_0 : std_logic;
signal \sEEDelayACQZ0Z_2\ : std_logic;
signal \sEEDelayACQ_i_2\ : std_logic;
signal un4_sacqtime_cry_1 : std_logic;
signal \sEEDelayACQZ0Z_3\ : std_logic;
signal \sEEDelayACQ_i_3\ : std_logic;
signal un4_sacqtime_cry_2 : std_logic;
signal \sEEDelayACQZ0Z_4\ : std_logic;
signal \sEEDelayACQ_i_4\ : std_logic;
signal un4_sacqtime_cry_3 : std_logic;
signal \sEEDelayACQZ0Z_5\ : std_logic;
signal \sEEDelayACQ_i_5\ : std_logic;
signal un4_sacqtime_cry_4 : std_logic;
signal \sEEDelayACQZ0Z_6\ : std_logic;
signal \sEEDelayACQ_i_6\ : std_logic;
signal un4_sacqtime_cry_5 : std_logic;
signal \sEEDelayACQZ0Z_7\ : std_logic;
signal \sEEDelayACQ_i_7\ : std_logic;
signal un4_sacqtime_cry_6 : std_logic;
signal un4_sacqtime_cry_7 : std_logic;
signal \sEEDelayACQZ0Z_8\ : std_logic;
signal \sEEDelayACQ_i_8\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \sEEDelayACQZ0Z_9\ : std_logic;
signal \sEEDelayACQ_i_9\ : std_logic;
signal un4_sacqtime_cry_8 : std_logic;
signal \sEEDelayACQZ0Z_10\ : std_logic;
signal \sEEDelayACQ_i_10\ : std_logic;
signal un4_sacqtime_cry_9 : std_logic;
signal \sEEDelayACQZ0Z_11\ : std_logic;
signal \sEEDelayACQ_i_11\ : std_logic;
signal un4_sacqtime_cry_10 : std_logic;
signal \sEEDelayACQZ0Z_12\ : std_logic;
signal \sEEDelayACQ_i_12\ : std_logic;
signal un4_sacqtime_cry_11 : std_logic;
signal \sEEDelayACQZ0Z_13\ : std_logic;
signal \sEEDelayACQ_i_13\ : std_logic;
signal un4_sacqtime_cry_12 : std_logic;
signal \sEEDelayACQZ0Z_14\ : std_logic;
signal \sEEDelayACQ_i_14\ : std_logic;
signal un4_sacqtime_cry_13 : std_logic;
signal \sEEDelayACQZ0Z_15\ : std_logic;
signal \sEEDelayACQ_i_15\ : std_logic;
signal un4_sacqtime_cry_14 : std_logic;
signal un4_sacqtime_cry_15 : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal un4_sacqtime_cry_16 : std_logic;
signal un4_sacqtime_cry_17 : std_logic;
signal un4_sacqtime_cry_18 : std_logic;
signal un4_sacqtime_cry_19 : std_logic;
signal g1_i_a4_4 : std_logic;
signal un4_sacqtime_cry_20 : std_logic;
signal un4_sacqtime_cry_21 : std_logic;
signal g0_4_0 : std_logic;
signal un4_sacqtime_cry_22 : std_logic;
signal un4_sacqtime_cry_23 : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal spi_sclk_ft_c : std_logic;
signal spi_sclk_rpi_c : std_logic;
signal spi_sclk : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_12\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9\ : std_logic;
signal \sDAC_mem_35Z0Z_3\ : std_logic;
signal \sDAC_data_2_6_bm_1_6_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_3\ : std_logic;
signal \sDAC_mem_8Z0Z_3\ : std_logic;
signal \sDAC_data_2_20_am_1_6_cascade_\ : std_logic;
signal \sDAC_mem_10Z0Z_3\ : std_logic;
signal \sDAC_mem_42Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_6_cascade_\ : std_logic;
signal \sDAC_mem_11Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_6\ : std_logic;
signal \sDAC_mem_2Z0Z_3\ : std_logic;
signal \sDAC_mem_7Z0Z_1\ : std_logic;
signal un1_spointer11_2_0_0_a2_5 : std_logic;
signal \N_183\ : std_logic;
signal \sPointerZ0Z_1\ : std_logic;
signal \sPointerZ0Z_0\ : std_logic;
signal \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1\ : std_logic;
signal \N_1624\ : std_logic;
signal \sDAC_mem_34Z0Z_3\ : std_logic;
signal \sDAC_mem_34_1_sqmuxa\ : std_logic;
signal \sDAC_mem_39Z0Z_1\ : std_logic;
signal \sDAC_mem_39_1_sqmuxa\ : std_logic;
signal \sEEPoffZ0Z_0\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \sEEPoffZ0Z_1\ : std_logic;
signal un1_spoff_cry_0 : std_logic;
signal \sEEPoffZ0Z_2\ : std_logic;
signal un1_spoff_cry_1 : std_logic;
signal \sEEPoffZ0Z_3\ : std_logic;
signal un1_spoff_cry_2 : std_logic;
signal \sEEPoffZ0Z_4\ : std_logic;
signal un1_spoff_cry_3 : std_logic;
signal \sEEPoffZ0Z_5\ : std_logic;
signal un1_spoff_cry_4 : std_logic;
signal \sEEPoffZ0Z_6\ : std_logic;
signal un1_spoff_cry_5 : std_logic;
signal \sEEPoffZ0Z_7\ : std_logic;
signal un1_spoff_cry_6 : std_logic;
signal un1_spoff_cry_7 : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal un1_spoff_cry_8 : std_logic;
signal \sEEPoffZ0Z_10\ : std_logic;
signal un1_spoff_cry_9 : std_logic;
signal un1_spoff_cry_10 : std_logic;
signal un1_spoff_cry_11 : std_logic;
signal un1_spoff_cry_12 : std_logic;
signal un1_spoff_cry_13 : std_logic;
signal un1_spoff_cry_14 : std_logic;
signal un1_spoff_cry_15 : std_logic;
signal \sCounter_i_16\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \sCounter_i_17\ : std_logic;
signal un1_spoff_cry_16 : std_logic;
signal \sCounter_i_18\ : std_logic;
signal un1_spoff_cry_17 : std_logic;
signal \sCounter_i_19\ : std_logic;
signal un1_spoff_cry_18 : std_logic;
signal \sCounter_i_20\ : std_logic;
signal un1_spoff_cry_19 : std_logic;
signal \sCounter_i_21\ : std_logic;
signal un1_spoff_cry_20 : std_logic;
signal \sCounter_i_22\ : std_logic;
signal un1_spoff_cry_21 : std_logic;
signal \sCounter_i_23\ : std_logic;
signal un1_spoff_cry_22 : std_logic;
signal un1_spoff_cry_23 : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \N_1683_i\ : std_logic;
signal \sbuttonModeStatusZ0\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_0\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_18\ : std_logic;
signal \sAddress_RNIA6242_1Z0Z_0\ : std_logic;
signal \sAddress_RNIA6242_0Z0Z_0\ : std_logic;
signal \sEEPoffZ0Z_11\ : std_logic;
signal \sEEPoffZ0Z_12\ : std_logic;
signal \sEEPoffZ0Z_13\ : std_logic;
signal \sEEPoffZ0Z_14\ : std_logic;
signal \sEEPoffZ0Z_15\ : std_logic;
signal \sEEPoffZ0Z_8\ : std_logic;
signal \sEEPoffZ0Z_9\ : std_logic;
signal \sAddress_RNIA6242_2Z0Z_0\ : std_logic;
signal \un4_sacqtime_cry_23_c_RNI2CQMZ0\ : std_logic;
signal \ADC5_c\ : std_logic;
signal \RAM_DATA_1Z0Z_5\ : std_logic;
signal \ADC1_c\ : std_logic;
signal \RAM_DATA_1Z0Z_1\ : std_logic;
signal \ADC9_c\ : std_logic;
signal \RAM_DATA_1Z0Z_10\ : std_logic;
signal top_tour1_c : std_logic;
signal \RAM_DATA_1Z0Z_11\ : std_logic;
signal \sTrigCounterZ0Z_0\ : std_logic;
signal \RAM_DATA_1Z0Z_13\ : std_logic;
signal \sTrigCounterZ0Z_1\ : std_logic;
signal \RAM_DATA_1Z0Z_14\ : std_logic;
signal \ADC2_c\ : std_logic;
signal \RAM_DATA_1Z0Z_2\ : std_logic;
signal \ADC6_c\ : std_logic;
signal \RAM_DATA_1Z0Z_6\ : std_logic;
signal \ADC0_c\ : std_logic;
signal \RAM_DATA_1Z0Z_0\ : std_logic;
signal \sDAC_mem_40Z0Z_3\ : std_logic;
signal \sDAC_mem_40_1_sqmuxa\ : std_logic;
signal \sDAC_mem_8_1_sqmuxa\ : std_logic;
signal \N_317\ : std_logic;
signal \sAddress_RNI6VH7_4Z0Z_1\ : std_logic;
signal \sAddress_RNI70I7Z0Z_1\ : std_logic;
signal \sAddress_RNIAM2A_0Z0Z_1\ : std_logic;
signal \sDAC_data_2_32_ns_1_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_6\ : std_logic;
signal \sDAC_data_2_14_ns_1_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_6\ : std_logic;
signal \sDAC_data_2_41_ns_1_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_6\ : std_logic;
signal \sDAC_data_2_6_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_6\ : std_logic;
signal \sDAC_mem_34Z0Z_5\ : std_logic;
signal \sDAC_mem_2Z0Z_5\ : std_logic;
signal \sDAC_mem_35Z0Z_5\ : std_logic;
signal \sDAC_data_2_6_bm_1_8_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_5\ : std_logic;
signal \sDAC_mem_42Z0Z_5\ : std_logic;
signal \sDAC_mem_10Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_8_cascade_\ : std_logic;
signal \sDAC_mem_11Z0Z_5\ : std_logic;
signal \sDAC_mem_40Z0Z_5\ : std_logic;
signal \sDAC_mem_8Z0Z_5\ : std_logic;
signal \sDAC_data_2_20_am_1_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_8\ : std_logic;
signal \sDAC_data_2_14_ns_1_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_8_cascade_\ : std_logic;
signal \sDAC_data_2_8_cascade_\ : std_logic;
signal \sDAC_data_2_32_ns_1_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_8_cascade_\ : std_logic;
signal \sDAC_data_2_41_ns_1_8\ : std_logic;
signal \sDAC_mem_34Z0Z_1\ : std_logic;
signal \sDAC_mem_2Z0Z_1\ : std_logic;
signal \sDAC_mem_3Z0Z_1\ : std_logic;
signal \sDAC_mem_35Z0Z_1\ : std_logic;
signal \sDAC_data_2_6_bm_1_4_cascade_\ : std_logic;
signal \sDAC_mem_42Z0Z_1\ : std_logic;
signal \sDAC_mem_10Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_4_cascade_\ : std_logic;
signal \sDAC_mem_11Z0Z_1\ : std_logic;
signal \sDAC_mem_40Z0Z_1\ : std_logic;
signal \sDAC_mem_8Z0Z_1\ : std_logic;
signal \sDAC_data_2_20_am_1_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_4\ : std_logic;
signal \sDAC_mem_15Z0Z_0\ : std_logic;
signal \sDAC_mem_14Z0Z_0\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_2_24_ns_1_4\ : std_logic;
signal \sDAC_mem_15Z0Z_1\ : std_logic;
signal \sDAC_mem_14Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_4\ : std_logic;
signal \sDAC_mem_12Z0Z_0\ : std_logic;
signal \sDAC_mem_12Z0Z_1\ : std_logic;
signal \sDAC_mem_31Z0Z_5\ : std_logic;
signal \sDAC_mem_30Z0Z_5\ : std_logic;
signal \sDAC_mem_29Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_8\ : std_logic;
signal \sDAC_mem_28Z0Z_5\ : std_logic;
signal \sDAC_mem_24Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_9_cascade_\ : std_logic;
signal \sDAC_data_2_39_ns_1_9_cascade_\ : std_logic;
signal \sDAC_mem_26Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_9\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_7_cascade_\ : std_logic;
signal \sDAC_data_2_39_ns_1_7_cascade_\ : std_logic;
signal \sDAC_mem_26Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_7\ : std_logic;
signal \sDAC_mem_29Z0Z_4\ : std_logic;
signal \sDAC_mem_28Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_7\ : std_logic;
signal \sDAC_mem_30Z0Z_4\ : std_logic;
signal \sDAC_mem_31Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_7\ : std_logic;
signal \sDAC_mem_24Z0Z_4\ : std_logic;
signal \sDAC_data_2_39_ns_1_8\ : std_logic;
signal \sDAC_mem_26Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_4\ : std_logic;
signal \sDAC_data_2_39_ns_1_4_cascade_\ : std_logic;
signal \sDAC_mem_28Z0Z_1\ : std_logic;
signal \sDAC_mem_29Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_4\ : std_logic;
signal \sDAC_mem_31Z0Z_1\ : std_logic;
signal \sDAC_mem_30Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_4\ : std_logic;
signal \sDAC_mem_24Z0Z_1\ : std_logic;
signal \sDAC_mem_24_1_sqmuxa\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_5\ : std_logic;
signal \sDAC_mem_26Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_8\ : std_logic;
signal \sDAC_mem_26Z0Z_5\ : std_logic;
signal \sDAC_mem_26_1_sqmuxa\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_clk_iZ0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.div_clk_iZ0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.falling_count_start_iZ0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.falling_count_start_i_i\ : std_logic;
signal \sCounter_i_0\ : std_logic;
signal \bfn_13_14_0_\ : std_logic;
signal \sCounter_i_1\ : std_logic;
signal un1_sacqtime_cry_0 : std_logic;
signal \sCounter_i_2\ : std_logic;
signal un1_sacqtime_cry_1 : std_logic;
signal \sCounter_i_3\ : std_logic;
signal un1_sacqtime_cry_2 : std_logic;
signal \sCounter_i_4\ : std_logic;
signal un1_sacqtime_cry_3 : std_logic;
signal \sCounter_i_5\ : std_logic;
signal un1_sacqtime_cry_4 : std_logic;
signal \sCounter_i_6\ : std_logic;
signal un1_sacqtime_cry_5 : std_logic;
signal \sCounter_i_7\ : std_logic;
signal un1_sacqtime_cry_6 : std_logic;
signal un1_sacqtime_cry_7 : std_logic;
signal \sCounter_i_8\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \sCounter_i_9\ : std_logic;
signal un1_sacqtime_cry_8 : std_logic;
signal \sCounter_i_10\ : std_logic;
signal un1_sacqtime_cry_9 : std_logic;
signal \sCounter_i_11\ : std_logic;
signal un1_sacqtime_cry_10 : std_logic;
signal \sCounter_i_12\ : std_logic;
signal un1_sacqtime_cry_11 : std_logic;
signal \sCounter_i_13\ : std_logic;
signal un1_sacqtime_cry_12 : std_logic;
signal \sCounter_i_14\ : std_logic;
signal un1_sacqtime_cry_13 : std_logic;
signal \sCounter_i_15\ : std_logic;
signal un1_sacqtime_cry_14 : std_logic;
signal un1_sacqtime_cry_15 : std_logic;
signal un1_sacqtime_cry_16_sf : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal un1_sacqtime_cry_17_sf : std_logic;
signal un1_sacqtime_cry_16 : std_logic;
signal un1_sacqtime_cry_18_sf : std_logic;
signal un1_sacqtime_cry_17 : std_logic;
signal un1_sacqtime_cry_19_sf : std_logic;
signal un1_sacqtime_cry_18 : std_logic;
signal un1_sacqtime_cry_20_sf : std_logic;
signal un1_sacqtime_cry_19 : std_logic;
signal un1_sacqtime_cry_21_sf : std_logic;
signal un1_sacqtime_cry_20 : std_logic;
signal un1_sacqtime_cry_22_sf : std_logic;
signal un1_sacqtime_cry_21 : std_logic;
signal un1_sacqtime_cry_23_sf : std_logic;
signal un1_sacqtime_cry_22 : std_logic;
signal un1_sacqtime_cry_23 : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \sADC_clk_prevZ0\ : std_logic;
signal \N_71_cascade_\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \sRAM_pointer_read_cry_0\ : std_logic;
signal \sRAM_pointer_read_cry_1\ : std_logic;
signal \sRAM_pointer_read_cry_2\ : std_logic;
signal \sRAM_pointer_read_cry_3\ : std_logic;
signal \sRAM_pointer_read_cry_4\ : std_logic;
signal \sRAM_pointer_read_cry_5\ : std_logic;
signal \sRAM_pointer_read_cry_6\ : std_logic;
signal \sRAM_pointer_read_cry_7\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \sRAM_pointer_read_cry_8\ : std_logic;
signal \sRAM_pointer_read_cry_9\ : std_logic;
signal \sRAM_pointer_read_cry_10\ : std_logic;
signal \sRAM_pointer_read_cry_11\ : std_logic;
signal \sRAM_pointer_read_cry_12\ : std_logic;
signal \sRAM_pointer_read_cry_13\ : std_logic;
signal \sRAM_pointer_read_cry_14\ : std_logic;
signal \sRAM_pointer_read_cry_15\ : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \sRAM_pointer_read_cry_16\ : std_logic;
signal \sRAM_pointer_read_cry_17\ : std_logic;
signal \N_28_g\ : std_logic;
signal \sDAC_mem_36_1_sqmuxa\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_6\ : std_logic;
signal \sDAC_mem_18Z0Z_3\ : std_logic;
signal \sDAC_mem_18Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_8\ : std_logic;
signal \sDAC_mem_18Z0Z_5\ : std_logic;
signal \sDAC_mem_18Z0Z_6\ : std_logic;
signal \sDAC_mem_18_1_sqmuxa\ : std_logic;
signal \sDAC_mem_15Z0Z_4\ : std_logic;
signal \sDAC_mem_14Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_8_cascade_\ : std_logic;
signal \sDAC_data_2_24_ns_1_8\ : std_logic;
signal \sDAC_mem_15Z0Z_5\ : std_logic;
signal \sDAC_mem_14Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_8\ : std_logic;
signal \sDAC_mem_12Z0Z_4\ : std_logic;
signal \sDAC_mem_12Z0Z_5\ : std_logic;
signal \sDAC_mem_38Z0Z_2\ : std_logic;
signal \sDAC_mem_39Z0Z_2\ : std_logic;
signal \sDAC_data_2_13_bm_1_5_cascade_\ : std_logic;
signal \sDAC_mem_6Z0Z_2\ : std_logic;
signal \sDAC_mem_38Z0Z_3\ : std_logic;
signal \sDAC_mem_39Z0Z_3\ : std_logic;
signal \sDAC_data_2_13_bm_1_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_6\ : std_logic;
signal \sDAC_mem_6Z0Z_3\ : std_logic;
signal \sDAC_mem_38Z0Z_4\ : std_logic;
signal \sDAC_mem_39Z0Z_4\ : std_logic;
signal \sDAC_data_2_13_bm_1_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_28Z0Z_6\ : std_logic;
signal \sDAC_mem_16Z0Z_3\ : std_logic;
signal \sDAC_mem_16Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_28Z0Z_8\ : std_logic;
signal \sDAC_mem_16Z0Z_5\ : std_logic;
signal \sDAC_mem_16Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_2_41_ns_1_4\ : std_logic;
signal \sDAC_data_2_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_4\ : std_logic;
signal \sDAC_data_2_14_ns_1_4\ : std_logic;
signal \sDAC_data_2_32_ns_1_4\ : std_logic;
signal \sDAC_mem_15Z0Z_2\ : std_logic;
signal \sDAC_mem_14Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_5_cascade_\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_6_cascade_\ : std_logic;
signal \sDAC_data_2_24_ns_1_6\ : std_logic;
signal \sDAC_mem_15Z0Z_3\ : std_logic;
signal \sDAC_mem_14Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_6\ : std_logic;
signal \sDAC_mem_12Z0Z_2\ : std_logic;
signal \sDAC_mem_12Z0Z_3\ : std_logic;
signal \sEEACQZ0Z_0\ : std_logic;
signal \sEEACQ_i_0\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \sEEACQZ0Z_1\ : std_logic;
signal \sEEACQ_i_1\ : std_logic;
signal un5_sdacdyn_cry_0 : std_logic;
signal \sEEACQZ0Z_2\ : std_logic;
signal \sEEACQ_i_2\ : std_logic;
signal un5_sdacdyn_cry_1 : std_logic;
signal \sEEACQZ0Z_3\ : std_logic;
signal \sEEACQ_i_3\ : std_logic;
signal un5_sdacdyn_cry_2 : std_logic;
signal \sEEACQZ0Z_4\ : std_logic;
signal \sEEACQ_i_4\ : std_logic;
signal un5_sdacdyn_cry_3 : std_logic;
signal \sEEACQZ0Z_5\ : std_logic;
signal \sEEACQ_i_5\ : std_logic;
signal un5_sdacdyn_cry_4 : std_logic;
signal \sEEACQZ0Z_6\ : std_logic;
signal \sEEACQ_i_6\ : std_logic;
signal un5_sdacdyn_cry_5 : std_logic;
signal \sEEACQZ0Z_7\ : std_logic;
signal \sEEACQ_i_7\ : std_logic;
signal un5_sdacdyn_cry_6 : std_logic;
signal un5_sdacdyn_cry_7 : std_logic;
signal \sEEACQZ0Z_8\ : std_logic;
signal \sEEACQ_i_8\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \sEEACQZ0Z_9\ : std_logic;
signal \sEEACQ_i_9\ : std_logic;
signal un5_sdacdyn_cry_8 : std_logic;
signal \sEEACQZ0Z_10\ : std_logic;
signal \sEEACQ_i_10\ : std_logic;
signal un5_sdacdyn_cry_9 : std_logic;
signal \sEEACQZ0Z_11\ : std_logic;
signal \sEEACQ_i_11\ : std_logic;
signal un5_sdacdyn_cry_10 : std_logic;
signal \sEEACQZ0Z_12\ : std_logic;
signal \sEEACQ_i_12\ : std_logic;
signal un5_sdacdyn_cry_11 : std_logic;
signal \sEEACQZ0Z_13\ : std_logic;
signal \sEEACQ_i_13\ : std_logic;
signal un5_sdacdyn_cry_12 : std_logic;
signal \sEEACQZ0Z_14\ : std_logic;
signal \sEEACQ_i_14\ : std_logic;
signal un5_sdacdyn_cry_13 : std_logic;
signal \sEEACQZ0Z_15\ : std_logic;
signal \sEEACQ_i_15\ : std_logic;
signal un5_sdacdyn_cry_14 : std_logic;
signal un5_sdacdyn_cry_15 : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal un5_sdacdyn_cry_16 : std_logic;
signal un5_sdacdyn_cry_17 : std_logic;
signal un5_sdacdyn_cry_18 : std_logic;
signal un5_sdacdyn_cry_19 : std_logic;
signal un5_sdacdyn_cry_20 : std_logic;
signal un5_sdacdyn_cry_21 : std_logic;
signal un5_sdacdyn_cry_22 : std_logic;
signal un5_sdacdyn_cry_23 : std_logic;
signal \N_106\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \sDAC_mem_24Z0Z_7\ : std_logic;
signal \sDAC_mem_26Z0Z_7\ : std_logic;
signal \sDAC_dataZ0Z_10\ : std_logic;
signal \sDAC_mem_24Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_5\ : std_logic;
signal \sDAC_mem_24Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_8\ : std_logic;
signal \sDAC_mem_29Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_9\ : std_logic;
signal \sDAC_mem_28Z0Z_6\ : std_logic;
signal \sDAC_mem_31Z0Z_0\ : std_logic;
signal \sDAC_mem_30Z0Z_0\ : std_logic;
signal \sDAC_mem_31Z0Z_3\ : std_logic;
signal \sDAC_mem_30Z0Z_3\ : std_logic;
signal \sDAC_mem_31Z0Z_6\ : std_logic;
signal \sDAC_mem_30Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_9\ : std_logic;
signal \sDAC_mem_16Z0Z_0\ : std_logic;
signal \sDAC_mem_16Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_28Z0Z_4\ : std_logic;
signal \sDAC_mem_16Z0Z_2\ : std_logic;
signal \sDAC_mem_27Z0Z_1\ : std_logic;
signal \sDAC_mem_27Z0Z_2\ : std_logic;
signal \sDAC_mem_27Z0Z_4\ : std_logic;
signal \sDAC_mem_27Z0Z_5\ : std_logic;
signal \sDAC_mem_27Z0Z_6\ : std_logic;
signal \sDAC_mem_27Z0Z_7\ : std_logic;
signal \sDAC_mem_27_1_sqmuxa\ : std_logic;
signal \sEEPonPoffZ0Z_0\ : std_logic;
signal un7_spon_0 : std_logic;
signal \sEEPonPoff_i_0\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal un7_spon_1 : std_logic;
signal \sEEPonPoffZ0Z_1\ : std_logic;
signal \sEEPonPoff_i_1\ : std_logic;
signal un4_spoff_cry_0 : std_logic;
signal \sEEPonPoffZ0Z_2\ : std_logic;
signal un7_spon_2 : std_logic;
signal \sEEPonPoff_i_2\ : std_logic;
signal un4_spoff_cry_1 : std_logic;
signal \sEEPonPoffZ0Z_3\ : std_logic;
signal un7_spon_3 : std_logic;
signal \sEEPonPoff_i_3\ : std_logic;
signal un4_spoff_cry_2 : std_logic;
signal \sEEPonPoffZ0Z_4\ : std_logic;
signal un7_spon_4 : std_logic;
signal \sEEPonPoff_i_4\ : std_logic;
signal un4_spoff_cry_3 : std_logic;
signal \sEEPonPoffZ0Z_5\ : std_logic;
signal un7_spon_5 : std_logic;
signal \sEEPonPoff_i_5\ : std_logic;
signal un4_spoff_cry_4 : std_logic;
signal \sEEPonPoffZ0Z_6\ : std_logic;
signal un7_spon_6 : std_logic;
signal \sEEPonPoff_i_6\ : std_logic;
signal un4_spoff_cry_5 : std_logic;
signal un7_spon_7 : std_logic;
signal \sEEPonPoffZ0Z_7\ : std_logic;
signal \sEEPonPoff_i_7\ : std_logic;
signal un4_spoff_cry_6 : std_logic;
signal un4_spoff_cry_7 : std_logic;
signal un7_spon_8 : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal un7_spon_9 : std_logic;
signal un4_spoff_cry_8 : std_logic;
signal un7_spon_10 : std_logic;
signal un4_spoff_cry_9 : std_logic;
signal un4_spoff_cry_10 : std_logic;
signal un7_spon_12 : std_logic;
signal un4_spoff_cry_11 : std_logic;
signal un7_spon_13 : std_logic;
signal un4_spoff_cry_12 : std_logic;
signal un7_spon_14 : std_logic;
signal un4_spoff_cry_13 : std_logic;
signal un7_spon_15 : std_logic;
signal un4_spoff_cry_14 : std_logic;
signal un4_spoff_cry_15 : std_logic;
signal un7_spon_16 : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal un7_spon_17 : std_logic;
signal un4_spoff_cry_16 : std_logic;
signal un7_spon_18 : std_logic;
signal un4_spoff_cry_17 : std_logic;
signal un4_spoff_cry_18 : std_logic;
signal un4_spoff_cry_19 : std_logic;
signal un4_spoff_cry_20 : std_logic;
signal un7_spon_22 : std_logic;
signal un4_spoff_cry_21 : std_logic;
signal un7_spon_23 : std_logic;
signal un4_spoff_cry_22 : std_logic;
signal un4_spoff_cry_23 : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \un4_spoff_cry_23_THRU_CO\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_3\ : std_logic;
signal \sDAC_dataZ0Z_4\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_4\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_7\ : std_logic;
signal \sDAC_dataZ0Z_8\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_9\ : std_logic;
signal \sEEDACZ0Z_1\ : std_logic;
signal \sEEDACZ0Z_3\ : std_logic;
signal \sEEDACZ0Z_5\ : std_logic;
signal \sEEDACZ0Z_7\ : std_logic;
signal \sEEDAC_1_sqmuxa\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_28Z0Z_7\ : std_logic;
signal \sDAC_data_2_32_ns_1_7\ : std_logic;
signal \sDAC_data_2_14_ns_1_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_7\ : std_logic;
signal \sDAC_data_2_41_ns_1_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_7\ : std_logic;
signal \sEEDACZ0Z_4\ : std_logic;
signal \sDAC_data_2_7_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_7\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_9_cascade_\ : std_logic;
signal \sEEDACZ0Z_6\ : std_logic;
signal \sDAC_data_2_9_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_9\ : std_logic;
signal \sDAC_data_2_14_ns_1_9\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_9\ : std_logic;
signal \sDAC_data_RNO_28Z0Z_9\ : std_logic;
signal \sDAC_data_2_32_ns_1_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_9\ : std_logic;
signal \sDAC_data_2_41_ns_1_9\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_8\ : std_logic;
signal \sDAC_mem_20Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_9\ : std_logic;
signal \sDAC_mem_20Z0Z_6\ : std_logic;
signal \sDAC_mem_22Z0Z_0\ : std_logic;
signal \sDAC_mem_22Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_4\ : std_logic;
signal \sDAC_mem_22Z0Z_2\ : std_logic;
signal \sDAC_mem_22Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_6\ : std_logic;
signal \sDAC_mem_36Z0Z_4\ : std_logic;
signal \sDAC_data_2_13_am_1_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_7\ : std_logic;
signal \sDAC_mem_4Z0Z_4\ : std_logic;
signal \sDAC_mem_36Z0Z_5\ : std_logic;
signal \sDAC_data_2_13_am_1_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_8\ : std_logic;
signal \sDAC_mem_38Z0Z_5\ : std_logic;
signal \sDAC_mem_39Z0Z_5\ : std_logic;
signal \sDAC_data_2_13_bm_1_8_cascade_\ : std_logic;
signal \sDAC_mem_7Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_8\ : std_logic;
signal \sDAC_mem_6Z0Z_5\ : std_logic;
signal \sDAC_mem_38Z0Z_6\ : std_logic;
signal \sDAC_data_2_13_bm_1_9_cascade_\ : std_logic;
signal \sDAC_mem_39Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_9\ : std_logic;
signal \sDAC_mem_6Z0Z_6\ : std_logic;
signal \sDAC_mem_40Z0Z_7\ : std_logic;
signal \sDAC_mem_8Z0Z_7\ : std_logic;
signal \sDAC_data_2_20_am_1_10_cascade_\ : std_logic;
signal \sDAC_mem_36Z0Z_6\ : std_logic;
signal \sDAC_data_2_13_am_1_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_9\ : std_logic;
signal \sDAC_mem_4Z0Z_6\ : std_logic;
signal \sDAC_mem_38Z0Z_7\ : std_logic;
signal \sDAC_mem_39Z0Z_7\ : std_logic;
signal \sDAC_data_2_13_bm_1_10_cascade_\ : std_logic;
signal \sDAC_mem_7Z0Z_7\ : std_logic;
signal \sDAC_mem_38Z0Z_0\ : std_logic;
signal \sDAC_mem_39Z0Z_0\ : std_logic;
signal \sDAC_data_2_13_bm_1_3_cascade_\ : std_logic;
signal \sDAC_mem_7Z0Z_0\ : std_logic;
signal \sDAC_mem_38Z0Z_1\ : std_logic;
signal \sDAC_data_2_13_bm_1_4\ : std_logic;
signal \sDAC_mem_34Z0Z_7\ : std_logic;
signal \sDAC_mem_2Z0Z_7\ : std_logic;
signal \sDAC_mem_2_1_sqmuxa\ : std_logic;
signal \sDAC_mem_12Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_10_cascade_\ : std_logic;
signal \sDAC_mem_15Z0Z_7\ : std_logic;
signal \sDAC_mem_14Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_10\ : std_logic;
signal \sDAC_mem_42Z0Z_7\ : std_logic;
signal \sDAC_mem_10Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_10_cascade_\ : std_logic;
signal \sDAC_mem_11Z0Z_7\ : std_logic;
signal \sDAC_data_2_24_ns_1_10\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_10_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_10\ : std_logic;
signal un7_spon_20 : std_logic;
signal un7_spon_19 : std_logic;
signal un7_spon_21 : std_logic;
signal un7_spon_11 : std_logic;
signal g0_12 : std_logic;
signal \sDAC_data_RNO_2Z0Z_10\ : std_logic;
signal \sDAC_data_2_41_ns_1_10_cascade_\ : std_logic;
signal \sDAC_data_2_10\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_17\ : std_logic;
signal \sDAC_mem_22Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_28Z0Z_10_cascade_\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_10\ : std_logic;
signal \sDAC_data_2_32_ns_1_10_cascade_\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_10\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_10\ : std_logic;
signal \sDAC_mem_18Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_10\ : std_logic;
signal \sDAC_mem_16Z0Z_7\ : std_logic;
signal \sDAC_mem_16_1_sqmuxa\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_10\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_10\ : std_logic;
signal \sDAC_mem_31Z0Z_7\ : std_logic;
signal \sDAC_mem_30Z0Z_7\ : std_logic;
signal \sDAC_mem_29Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_10\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_10_cascade_\ : std_logic;
signal \sDAC_data_2_39_ns_1_10\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_10\ : std_logic;
signal \sDAC_mem_28Z0Z_7\ : std_logic;
signal \sDAC_mem_27Z0Z_0\ : std_logic;
signal \sDAC_mem_26Z0Z_0\ : std_logic;
signal \sDAC_mem_24Z0Z_0\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_3\ : std_logic;
signal \sDAC_data_2_39_ns_1_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_7\ : std_logic;
signal \sDAC_mem_22Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_8\ : std_logic;
signal \sDAC_mem_22Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_9\ : std_logic;
signal \sDAC_mem_22Z0Z_6\ : std_logic;
signal \sDAC_mem_22_1_sqmuxa\ : std_logic;
signal \sDAC_mem_29Z0Z_0\ : std_logic;
signal \sDAC_mem_28Z0Z_0\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_3\ : std_logic;
signal \sDAC_mem_29Z0Z_3\ : std_logic;
signal \sDAC_mem_28Z0Z_3\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_14_cascade_\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_13\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_22\ : std_logic;
signal \sEEPonPoff_1_sqmuxa_0_a3_0_a2_1\ : std_logic;
signal \sPointer_RNI5LBD1Z0Z_0\ : std_logic;
signal \sEEPonPoff_1_sqmuxa\ : std_logic;
signal \RAM_nWE_0_i\ : std_logic;
signal \sRead_data_RNOZ0Z_0_cascade_\ : std_logic;
signal \ADC_clk_c\ : std_logic;
signal \sRead_dataZ0\ : std_logic;
signal spi_data_miso_0_sqmuxa_2_i_o2_4 : std_logic;
signal spi_data_miso_0_sqmuxa_2_i_o2_5 : std_logic;
signal \ADC3_c\ : std_logic;
signal \RAM_DATA_1Z0Z_3\ : std_logic;
signal \sDAC_mem_19Z0Z_4\ : std_logic;
signal \sDAC_mem_19Z0Z_5\ : std_logic;
signal \sDAC_mem_19Z0Z_6\ : std_logic;
signal \sDAC_mem_19Z0Z_7\ : std_logic;
signal \sDAC_mem_21Z0Z_5\ : std_logic;
signal \sDAC_mem_21Z0Z_6\ : std_logic;
signal \sDAC_mem_21Z0Z_7\ : std_logic;
signal \sDAC_mem_21_1_sqmuxa\ : std_logic;
signal \sDAC_mem_34Z0Z_4\ : std_logic;
signal \sDAC_mem_2Z0Z_4\ : std_logic;
signal \sDAC_mem_35Z0Z_4\ : std_logic;
signal \sDAC_data_2_6_bm_1_7_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_7\ : std_logic;
signal \sDAC_mem_40Z0Z_4\ : std_logic;
signal \sDAC_mem_8Z0Z_4\ : std_logic;
signal \sDAC_data_2_20_am_1_7_cascade_\ : std_logic;
signal \sDAC_data_2_24_ns_1_7\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_7\ : std_logic;
signal \sDAC_mem_11Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_7\ : std_logic;
signal \sDAC_mem_42Z0Z_4\ : std_logic;
signal \sDAC_mem_10Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_7\ : std_logic;
signal \sDAC_mem_34Z0Z_6\ : std_logic;
signal \sDAC_mem_2Z0Z_6\ : std_logic;
signal \sDAC_mem_35Z0Z_6\ : std_logic;
signal \sDAC_data_2_6_bm_1_9_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_9\ : std_logic;
signal \sDAC_mem_42Z0Z_6\ : std_logic;
signal \sDAC_mem_10Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_9_cascade_\ : std_logic;
signal \sDAC_mem_11Z0Z_6\ : std_logic;
signal \sDAC_mem_40Z0Z_6\ : std_logic;
signal \sDAC_mem_8Z0Z_6\ : std_logic;
signal \sDAC_data_2_20_am_1_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_9\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_9\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_9_cascade_\ : std_logic;
signal \sDAC_mem_32Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_9\ : std_logic;
signal \sDAC_mem_21Z0Z_0\ : std_logic;
signal \sDAC_mem_21Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_4\ : std_logic;
signal \sDAC_mem_21Z0Z_2\ : std_logic;
signal \sDAC_mem_21Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_6\ : std_logic;
signal \sDAC_mem_21Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_7\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \sDAC_mem_pointer_0_cry_1\ : std_logic;
signal \sDAC_mem_pointer_0_cry_2\ : std_logic;
signal \sDAC_mem_pointer_0_cry_3\ : std_logic;
signal \sDAC_mem_pointer_0_cry_4\ : std_logic;
signal \sDAC_mem_34Z0Z_2\ : std_logic;
signal \sDAC_mem_2Z0Z_2\ : std_logic;
signal \sDAC_mem_35Z0Z_2\ : std_logic;
signal \sDAC_data_2_6_bm_1_5_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_2\ : std_logic;
signal \sDAC_mem_42Z0Z_2\ : std_logic;
signal \sDAC_mem_10Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_5_cascade_\ : std_logic;
signal \sDAC_mem_11Z0Z_2\ : std_logic;
signal \sDAC_mem_40Z0Z_2\ : std_logic;
signal \sDAC_mem_8Z0Z_2\ : std_logic;
signal \sDAC_data_2_20_am_1_5_cascade_\ : std_logic;
signal \sDAC_data_2_24_ns_1_5\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_5_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_5\ : std_logic;
signal \sDAC_mem_34Z0Z_0\ : std_logic;
signal \sDAC_mem_2Z0Z_0\ : std_logic;
signal \sDAC_mem_35Z0Z_0\ : std_logic;
signal \sDAC_data_2_6_bm_1_3_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_0\ : std_logic;
signal \sDAC_mem_42Z0Z_0\ : std_logic;
signal \sDAC_mem_10Z0Z_0\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_3_cascade_\ : std_logic;
signal \sDAC_mem_11Z0Z_0\ : std_logic;
signal \sDAC_mem_40Z0Z_0\ : std_logic;
signal \sDAC_mem_8Z0Z_0\ : std_logic;
signal \sDAC_data_2_20_am_1_3_cascade_\ : std_logic;
signal \sDAC_data_2_24_ns_1_3\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_3\ : std_logic;
signal \N_333\ : std_logic;
signal \sDAC_mem_19Z0Z_0\ : std_logic;
signal \sDAC_mem_18Z0Z_0\ : std_logic;
signal \sDAC_mem_19Z0Z_1\ : std_logic;
signal \sDAC_mem_18Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_4\ : std_logic;
signal \sDAC_mem_19Z0Z_2\ : std_logic;
signal \sDAC_mem_18Z0Z_2\ : std_logic;
signal \sDAC_mem_19Z0Z_3\ : std_logic;
signal \sDAC_mem_19_1_sqmuxa\ : std_logic;
signal \sDAC_mem_35Z0Z_7\ : std_logic;
signal \sDAC_data_2_6_bm_1_10\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_10_cascade_\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_10\ : std_logic;
signal \sDAC_data_2_14_ns_1_10_cascade_\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_10\ : std_logic;
signal \sDAC_mem_36Z0Z_7\ : std_logic;
signal \sDAC_data_2_13_am_1_10_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_10\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_10\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_10\ : std_logic;
signal \bfn_16_13_0_\ : std_logic;
signal \button_debounce_counterZ0Z_2\ : std_logic;
signal un1_button_debounce_counter_cry_1 : std_logic;
signal \button_debounce_counterZ0Z_3\ : std_logic;
signal un1_button_debounce_counter_cry_2 : std_logic;
signal \button_debounce_counterZ0Z_4\ : std_logic;
signal un1_button_debounce_counter_cry_3 : std_logic;
signal \button_debounce_counterZ0Z_5\ : std_logic;
signal un1_button_debounce_counter_cry_4 : std_logic;
signal \button_debounce_counterZ0Z_6\ : std_logic;
signal un1_button_debounce_counter_cry_5 : std_logic;
signal un1_button_debounce_counter_cry_6 : std_logic;
signal un1_button_debounce_counter_cry_7 : std_logic;
signal un1_button_debounce_counter_cry_8 : std_logic;
signal \bfn_16_14_0_\ : std_logic;
signal un1_button_debounce_counter_cry_9 : std_logic;
signal un1_button_debounce_counter_cry_10 : std_logic;
signal un1_button_debounce_counter_cry_11 : std_logic;
signal un1_button_debounce_counter_cry_12 : std_logic;
signal un1_button_debounce_counter_cry_13 : std_logic;
signal \button_debounce_counterZ0Z_15\ : std_logic;
signal un1_button_debounce_counter_cry_14 : std_logic;
signal \button_debounce_counterZ0Z_16\ : std_logic;
signal un1_button_debounce_counter_cry_15 : std_logic;
signal un1_button_debounce_counter_cry_16 : std_logic;
signal \button_debounce_counterZ0Z_17\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \button_debounce_counterZ0Z_18\ : std_logic;
signal un1_button_debounce_counter_cry_17 : std_logic;
signal \button_debounce_counterZ0Z_19\ : std_logic;
signal un1_button_debounce_counter_cry_18 : std_logic;
signal \button_debounce_counterZ0Z_20\ : std_logic;
signal un1_button_debounce_counter_cry_19 : std_logic;
signal \button_debounce_counterZ0Z_21\ : std_logic;
signal un1_button_debounce_counter_cry_20 : std_logic;
signal \button_debounce_counterZ0Z_22\ : std_logic;
signal un1_button_debounce_counter_cry_21 : std_logic;
signal un1_button_debounce_counter_cry_22 : std_logic;
signal \un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO\ : std_logic;
signal \un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \button_debounce_counterZ0Z_23\ : std_logic;
signal \LED3_c_0\ : std_logic;
signal \sRAM_pointer_readZ0Z_5\ : std_logic;
signal \sRAM_pointer_writeZ0Z_5\ : std_logic;
signal \RAM_ADD_c_5\ : std_logic;
signal \sRAM_pointer_readZ0Z_0\ : std_logic;
signal \sRAM_pointer_writeZ0Z_0\ : std_logic;
signal \RAM_ADD_c_0\ : std_logic;
signal \sRAM_pointer_readZ0Z_10\ : std_logic;
signal \sRAM_pointer_writeZ0Z_10\ : std_logic;
signal \RAM_ADD_c_10\ : std_logic;
signal \sRAM_pointer_readZ0Z_11\ : std_logic;
signal \sRAM_pointer_writeZ0Z_11\ : std_logic;
signal \RAM_ADD_c_11\ : std_logic;
signal \sRAM_pointer_writeZ0Z_12\ : std_logic;
signal \sRAM_pointer_readZ0Z_12\ : std_logic;
signal \RAM_ADD_c_12\ : std_logic;
signal \sRAM_pointer_readZ0Z_13\ : std_logic;
signal \sRAM_pointer_writeZ0Z_13\ : std_logic;
signal \RAM_ADD_c_13\ : std_logic;
signal \sRAM_pointer_writeZ0Z_14\ : std_logic;
signal \sRAM_pointer_readZ0Z_14\ : std_logic;
signal \RAM_ADD_c_14\ : std_logic;
signal \sRAM_pointer_readZ0Z_15\ : std_logic;
signal \sRAM_pointer_writeZ0Z_15\ : std_logic;
signal \RAM_ADD_c_15\ : std_logic;
signal \sRAM_pointer_readZ0Z_16\ : std_logic;
signal \sRAM_pointer_writeZ0Z_16\ : std_logic;
signal \RAM_ADD_c_16\ : std_logic;
signal \sRAM_pointer_writeZ0Z_17\ : std_logic;
signal \sRAM_pointer_readZ0Z_17\ : std_logic;
signal \RAM_ADD_c_17\ : std_logic;
signal \sRAM_pointer_writeZ0Z_18\ : std_logic;
signal \sRAM_pointer_readZ0Z_18\ : std_logic;
signal \RAM_ADD_c_18\ : std_logic;
signal \sRAM_pointer_writeZ0Z_9\ : std_logic;
signal \sRAM_pointer_readZ0Z_9\ : std_logic;
signal \RAM_ADD_c_9\ : std_logic;
signal \sRAM_pointer_writeZ0Z_7\ : std_logic;
signal \sRAM_pointer_readZ0Z_7\ : std_logic;
signal \RAM_ADD_c_7\ : std_logic;
signal \sRAM_pointer_readZ0Z_2\ : std_logic;
signal \sRAM_pointer_writeZ0Z_2\ : std_logic;
signal \RAM_ADD_c_2\ : std_logic;
signal \sRAM_pointer_writeZ0Z_1\ : std_logic;
signal \sRAM_pointer_readZ0Z_1\ : std_logic;
signal \RAM_ADD_c_1\ : std_logic;
signal \sRAM_pointer_writeZ0Z_6\ : std_logic;
signal \sRAM_pointer_readZ0Z_6\ : std_logic;
signal \RAM_ADD_c_6\ : std_logic;
signal \ADC4_c\ : std_logic;
signal \RAM_DATA_1Z0Z_4\ : std_logic;
signal \sDAC_mem_4Z0Z_5\ : std_logic;
signal \sDAC_mem_4Z0Z_7\ : std_logic;
signal \sDAC_mem_20Z0Z_0\ : std_logic;
signal \sDAC_mem_20Z0Z_1\ : std_logic;
signal \sDAC_mem_20Z0Z_2\ : std_logic;
signal \sDAC_mem_20Z0Z_3\ : std_logic;
signal \sDAC_mem_20Z0Z_4\ : std_logic;
signal \sDAC_mem_20Z0Z_7\ : std_logic;
signal \sDAC_mem_20_1_sqmuxa\ : std_logic;
signal \sDAC_mem_6Z0Z_0\ : std_logic;
signal \sDAC_mem_6Z0Z_1\ : std_logic;
signal \sDAC_mem_6Z0Z_4\ : std_logic;
signal \sDAC_mem_6Z0Z_7\ : std_logic;
signal \sDAC_mem_6_1_sqmuxa\ : std_logic;
signal \sDAC_mem_23Z0Z_0\ : std_logic;
signal \sDAC_mem_23Z0Z_1\ : std_logic;
signal \sDAC_mem_23Z0Z_2\ : std_logic;
signal \sDAC_mem_23Z0Z_3\ : std_logic;
signal \sDAC_mem_23Z0Z_4\ : std_logic;
signal \sDAC_mem_23Z0Z_5\ : std_logic;
signal \sDAC_mem_23Z0Z_6\ : std_logic;
signal \sDAC_mem_23Z0Z_7\ : std_logic;
signal \sDAC_mem_23_1_sqmuxa\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_6_cascade_\ : std_logic;
signal \sDAC_mem_32Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_7\ : std_logic;
signal \sDAC_mem_32Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_8\ : std_logic;
signal \sDAC_mem_9Z0Z_0\ : std_logic;
signal \sDAC_mem_9Z0Z_1\ : std_logic;
signal \sDAC_mem_9Z0Z_2\ : std_logic;
signal \sDAC_mem_9Z0Z_3\ : std_logic;
signal \sDAC_mem_9Z0Z_4\ : std_logic;
signal \sDAC_mem_9Z0Z_5\ : std_logic;
signal \sDAC_mem_9Z0Z_6\ : std_logic;
signal \sDAC_mem_9Z0Z_7\ : std_logic;
signal \sDAC_mem_15Z0Z_6\ : std_logic;
signal \sDAC_mem_14Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_9\ : std_logic;
signal \sDAC_data_2_24_ns_1_9\ : std_logic;
signal \sDAC_mem_12Z0Z_6\ : std_logic;
signal \sDAC_mem_12_1_sqmuxa\ : std_logic;
signal \op_le_op_le_un15_sdacdynlt4_cascade_\ : std_logic;
signal un17_sdacdyn_1 : std_logic;
signal \sDAC_mem_pointerZ0Z_7\ : std_logic;
signal \sDAC_mem_pointerZ0Z_6\ : std_logic;
signal un17_sdacdyn_0 : std_logic;
signal \sDAC_data_RNO_5Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_5_cascade_\ : std_logic;
signal \sEEDACZ0Z_2\ : std_logic;
signal \sDAC_data_2_5_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_5\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_5\ : std_logic;
signal \sDAC_data_2_14_ns_1_5\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_28Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_5\ : std_logic;
signal \sDAC_data_2_32_ns_1_5_cascade_\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_5_cascade_\ : std_logic;
signal \sDAC_data_2_41_ns_1_5\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \sEEDACZ0Z_0\ : std_logic;
signal \sDAC_data_2_3_cascade_\ : std_logic;
signal \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\ : std_logic;
signal \sDAC_dataZ0Z_3\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_3\ : std_logic;
signal \sDAC_mem_pointerZ0Z_4\ : std_logic;
signal \sDAC_mem_pointerZ0Z_3\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_3\ : std_logic;
signal \sDAC_data_2_41_ns_1_3\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_3\ : std_logic;
signal \sDAC_data_2_14_ns_1_3\ : std_logic;
signal \sDAC_data_RNO_28Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_3\ : std_logic;
signal \sDAC_data_2_32_ns_1_3\ : std_logic;
signal \sDAC_data_2_39_ns_1_5\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_5\ : std_logic;
signal \sDAC_mem_29Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_5\ : std_logic;
signal \sDAC_mem_24Z0Z_3\ : std_logic;
signal \sDAC_mem_pointerZ0Z_1\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_6_cascade_\ : std_logic;
signal \sDAC_mem_pointerZ0Z_2\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_6\ : std_logic;
signal \sDAC_data_2_39_ns_1_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_6\ : std_logic;
signal \sDAC_mem_28Z0Z_2\ : std_logic;
signal \sDAC_mem_28_1_sqmuxa\ : std_logic;
signal \sDAC_mem_30Z0Z_2\ : std_logic;
signal \sDAC_mem_31Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_5\ : std_logic;
signal \sDAC_mem_26Z0Z_3\ : std_logic;
signal \sDAC_mem_27Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_6\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5\ : std_logic;
signal \sDAC_mem_17Z0Z_0\ : std_logic;
signal \sDAC_mem_17Z0Z_1\ : std_logic;
signal \sDAC_mem_17Z0Z_2\ : std_logic;
signal \sDAC_mem_17Z0Z_3\ : std_logic;
signal \sDAC_mem_17Z0Z_4\ : std_logic;
signal \sDAC_mem_17Z0Z_5\ : std_logic;
signal \sDAC_mem_17Z0Z_6\ : std_logic;
signal \sDAC_mem_17Z0Z_7\ : std_logic;
signal \RAM_DATA_in_14\ : std_logic;
signal \RAM_DATA_in_6\ : std_logic;
signal \button_debounce_counterZ0Z_13\ : std_logic;
signal \button_debounce_counterZ0Z_12\ : std_logic;
signal \button_debounce_counterZ0Z_14\ : std_logic;
signal \button_debounce_counterZ0Z_11\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_15\ : std_logic;
signal \button_debounce_counterZ0Z_9\ : std_logic;
signal \button_debounce_counterZ0Z_7\ : std_logic;
signal \button_debounce_counterZ0Z_10\ : std_logic;
signal \button_debounce_counterZ0Z_8\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_16\ : std_logic;
signal \RAM_DATA_in_0\ : std_logic;
signal \RAM_DATA_in_8\ : std_logic;
signal \RAM_DATA_in_12\ : std_logic;
signal \RAM_DATA_in_4\ : std_logic;
signal \sEEPointerResetZ0\ : std_logic;
signal \un4_sacqtime_cry_23_c_RNITTSZ0Z3_cascade_\ : std_logic;
signal \N_28\ : std_logic;
signal \sSPI_MSB0LSBZ0Z1\ : std_logic;
signal \spi_mosi_ready_prev3_RNILKERZ0\ : std_logic;
signal \RAM_DATA_cl_11Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_12Z0Z_15\ : std_logic;
signal \sCounterRAMZ0Z_0\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \sCounterRAMZ0Z_1\ : std_logic;
signal \sCounterRAM_cry_0\ : std_logic;
signal \sCounterRAMZ0Z_2\ : std_logic;
signal \sCounterRAM_cry_1\ : std_logic;
signal \sCounterRAMZ0Z_3\ : std_logic;
signal \sCounterRAM_cry_2\ : std_logic;
signal \sCounterRAMZ0Z_4\ : std_logic;
signal \sCounterRAM_cry_3\ : std_logic;
signal \sCounterRAMZ0Z_5\ : std_logic;
signal \sCounterRAM_cry_4\ : std_logic;
signal \sCounterRAMZ0Z_6\ : std_logic;
signal \sCounterRAM_cry_5\ : std_logic;
signal \N_70_i\ : std_logic;
signal \sCounterRAM_cry_6\ : std_logic;
signal \sCounterRAMZ0Z_7\ : std_logic;
signal \RAM_DATA_cl_6Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_7Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_8Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_9Z0Z_15\ : std_logic;
signal \RAM_DATA_clZ0Z_15\ : std_logic;
signal \RAM_DATA_1Z0Z_7\ : std_logic;
signal \sDAC_mem_41Z0Z_4\ : std_logic;
signal \sDAC_mem_36Z0Z_3\ : std_logic;
signal \sDAC_mem_4Z0Z_3\ : std_logic;
signal \sDAC_data_2_13_am_1_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_6\ : std_logic;
signal \sDAC_mem_32Z0Z_5\ : std_logic;
signal \sDAC_mem_32Z0Z_7\ : std_logic;
signal \sDAC_mem_41Z0Z_0\ : std_logic;
signal \sDAC_mem_41Z0Z_1\ : std_logic;
signal \sDAC_mem_41Z0Z_2\ : std_logic;
signal \sDAC_mem_41Z0Z_3\ : std_logic;
signal \sDAC_mem_41Z0Z_5\ : std_logic;
signal \sDAC_mem_41Z0Z_6\ : std_logic;
signal \sDAC_mem_41Z0Z_7\ : std_logic;
signal \sDAC_mem_9_1_sqmuxa\ : std_logic;
signal \sDAC_mem_41_1_sqmuxa\ : std_logic;
signal \sAddress_RNI6VH7_6Z0Z_1\ : std_logic;
signal \sAddress_RNI6VH7_6Z0Z_1_cascade_\ : std_logic;
signal \sAddressZ0Z_5\ : std_logic;
signal \sAddress_RNIP2UK1Z0Z_4\ : std_logic;
signal \sAddressZ0Z_2\ : std_logic;
signal \sAddressZ0Z_1\ : std_logic;
signal \sAddressZ0Z_3\ : std_logic;
signal \sAddressZ0Z_0\ : std_logic;
signal \sAddress_RNIAM2A_1Z0Z_1\ : std_logic;
signal \sAddress_RNIAM2A_1Z0Z_1_cascade_\ : std_logic;
signal \sAddress_RNIVREN1Z0Z_4\ : std_logic;
signal \sDAC_mem_17_1_sqmuxa\ : std_logic;
signal \sDAC_mem_37Z0Z_3\ : std_logic;
signal \sDAC_mem_37Z0Z_4\ : std_logic;
signal \sDAC_mem_37Z0Z_5\ : std_logic;
signal \sDAC_mem_37Z0Z_6\ : std_logic;
signal \sDAC_mem_37Z0Z_7\ : std_logic;
signal \sDAC_mem_37_1_sqmuxa\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_4\ : std_logic;
signal \sDAC_mem_32Z0Z_0\ : std_logic;
signal \sDAC_mem_32Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_5_cascade_\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_5\ : std_logic;
signal \sDAC_mem_32Z0Z_2\ : std_logic;
signal \sDAC_mem_32_1_sqmuxa\ : std_logic;
signal \sDAC_mem_36Z0Z_0\ : std_logic;
signal \sDAC_mem_37Z0Z_0\ : std_logic;
signal \sDAC_data_2_13_am_1_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_3\ : std_logic;
signal \sDAC_mem_4Z0Z_0\ : std_logic;
signal \sDAC_mem_36Z0Z_1\ : std_logic;
signal \sDAC_data_2_13_am_1_4_cascade_\ : std_logic;
signal \sDAC_mem_37Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_4\ : std_logic;
signal \sDAC_mem_4Z0Z_1\ : std_logic;
signal \sDAC_mem_4_1_sqmuxa\ : std_logic;
signal \sDAC_mem_pointerZ0Z_5\ : std_logic;
signal \sDAC_mem_36Z0Z_2\ : std_logic;
signal \sDAC_mem_4Z0Z_2\ : std_logic;
signal \sDAC_mem_pointerZ0Z_0\ : std_logic;
signal \sDAC_mem_37Z0Z_2\ : std_logic;
signal \sDAC_data_2_13_am_1_5_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_5\ : std_logic;
signal \sDAC_mem_25Z0Z_5\ : std_logic;
signal \sDAC_mem_25Z0Z_2\ : std_logic;
signal \sDAC_mem_25Z0Z_3\ : std_logic;
signal \sDAC_mem_25Z0Z_4\ : std_logic;
signal \sDAC_mem_25Z0Z_0\ : std_logic;
signal \sDAC_mem_25Z0Z_6\ : std_logic;
signal \sDAC_mem_25Z0Z_7\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1\ : std_logic;
signal \spi_slave_inst.un23_i_ssn\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2\ : std_logic;
signal \spi_data_misoZ0Z_0\ : std_logic;
signal \spi_data_misoZ0Z_4\ : std_logic;
signal \spi_data_misoZ0Z_6\ : std_logic;
signal \spi_slave_inst.un4_i_wr\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \sCounterADC_cry_0\ : std_logic;
signal \sCounterADC_cry_1\ : std_logic;
signal \sCounterADC_cry_2\ : std_logic;
signal \sCounterADCZ0Z_4\ : std_logic;
signal \sCounterADC_cry_3\ : std_logic;
signal \sCounterADCZ0Z_5\ : std_logic;
signal \sCounterADC_cry_4\ : std_logic;
signal \sCounterADC_cry_5\ : std_logic;
signal \sCounterADC_cry_6\ : std_logic;
signal \RAM_DATA_in_5\ : std_logic;
signal \RAM_DATA_in_13\ : std_logic;
signal \spi_data_misoZ0Z_5\ : std_logic;
signal \RAM_DATA_in_15\ : std_logic;
signal \RAM_DATA_in_7\ : std_logic;
signal \spi_data_misoZ0Z_7\ : std_logic;
signal \RAM_DATA_in_3\ : std_logic;
signal \RAM_DATA_in_11\ : std_logic;
signal \spi_data_misoZ0Z_3\ : std_logic;
signal \RAM_DATA_in_10\ : std_logic;
signal \RAM_DATA_in_2\ : std_logic;
signal \spi_data_misoZ0Z_2\ : std_logic;
signal \RAM_DATA_in_1\ : std_logic;
signal \RAM_DATA_in_9\ : std_logic;
signal \N_75\ : std_logic;
signal \spi_data_misoZ0Z_1\ : std_logic;
signal \sSPI_MSB0LSB1_RNIGRPGZ0Z4\ : std_logic;
signal \sRAM_pointer_writeZ0Z_8\ : std_logic;
signal \sRAM_pointer_readZ0Z_8\ : std_logic;
signal \RAM_ADD_c_8\ : std_logic;
signal \sRAM_pointer_writeZ0Z_4\ : std_logic;
signal \sRAM_pointer_readZ0Z_4\ : std_logic;
signal \RAM_ADD_c_4\ : std_logic;
signal \sRAM_pointer_writeZ0Z_3\ : std_logic;
signal \un1_sacqtime_cry_23_THRU_CO\ : std_logic;
signal \sRAM_pointer_readZ0Z_3\ : std_logic;
signal \un4_sacqtime_cry_23_THRU_CO\ : std_logic;
signal \RAM_ADD_c_3\ : std_logic;
signal \N_67_i\ : std_logic;
signal \RAM_DATA_cl_13Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_14Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_15Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_1Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_10Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_3Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_4Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_2Z0Z_15\ : std_logic;
signal \GNDG0\ : std_logic;
signal op_eq_scounterdac10_g : std_logic;
signal \sDAC_dataZ0Z_2\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_ready_iZ0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_2\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2\ : std_logic;
signal \sDAC_mem_7Z0Z_2\ : std_logic;
signal \sDAC_mem_7Z0Z_3\ : std_logic;
signal \sDAC_mem_7Z0Z_4\ : std_logic;
signal \sDAC_mem_7Z0Z_6\ : std_logic;
signal \sDAC_mem_7_1_sqmuxa\ : std_logic;
signal \sDAC_mem_3Z0Z_7\ : std_logic;
signal \sDAC_mem_3_1_sqmuxa\ : std_logic;
signal \sDAC_mem_1Z0Z_0\ : std_logic;
signal \sDAC_mem_1Z0Z_1\ : std_logic;
signal \sDAC_mem_1Z0Z_2\ : std_logic;
signal \sDAC_mem_1Z0Z_3\ : std_logic;
signal \sDAC_mem_1Z0Z_4\ : std_logic;
signal \sDAC_mem_1Z0Z_5\ : std_logic;
signal \sDAC_mem_1Z0Z_6\ : std_logic;
signal \sDAC_mem_1Z0Z_7\ : std_logic;
signal \sDAC_mem_1_1_sqmuxa\ : std_logic;
signal \sDAC_mem_33Z0Z_0\ : std_logic;
signal \sDAC_mem_33Z0Z_1\ : std_logic;
signal \sDAC_mem_33Z0Z_2\ : std_logic;
signal \sDAC_mem_33Z0Z_3\ : std_logic;
signal \sDAC_mem_33Z0Z_4\ : std_logic;
signal \sDAC_mem_33Z0Z_5\ : std_logic;
signal \sDAC_mem_33Z0Z_6\ : std_logic;
signal \sDAC_mem_33Z0Z_7\ : std_logic;
signal \sDAC_mem_33_1_sqmuxa\ : std_logic;
signal \sDAC_mem_5Z0Z_0\ : std_logic;
signal \sDAC_mem_5Z0Z_1\ : std_logic;
signal \sDAC_mem_5Z0Z_2\ : std_logic;
signal \sDAC_mem_5Z0Z_3\ : std_logic;
signal \sDAC_mem_5Z0Z_4\ : std_logic;
signal \sDAC_mem_5Z0Z_5\ : std_logic;
signal \sDAC_mem_5Z0Z_6\ : std_logic;
signal \sDAC_mem_5Z0Z_7\ : std_logic;
signal \sDAC_mem_5_1_sqmuxa\ : std_logic;
signal \sDAC_mem_13Z0Z_0\ : std_logic;
signal \sDAC_mem_13Z0Z_1\ : std_logic;
signal \sDAC_mem_13Z0Z_2\ : std_logic;
signal \sDAC_mem_13Z0Z_3\ : std_logic;
signal spi_data_mosi_4 : std_logic;
signal \sDAC_mem_13Z0Z_4\ : std_logic;
signal spi_data_mosi_5 : std_logic;
signal \sDAC_mem_13Z0Z_5\ : std_logic;
signal \sDAC_mem_13Z0Z_6\ : std_logic;
signal \sDAC_mem_13Z0Z_7\ : std_logic;
signal \sDAC_mem_13_1_sqmuxa\ : std_logic;
signal \spi_slave_inst.tx_ready_iZ0\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_0\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_2\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_2\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_1\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_1\ : std_logic;
signal \button_debounce_counterZ0Z_1\ : std_logic;
signal \button_debounce_counterZ0Z_0\ : std_logic;
signal \N_3154_g\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_6\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_6\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_5\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_5\ : std_logic;
signal spi_data_mosi_2 : std_logic;
signal \sCounterADCZ0Z_2\ : std_logic;
signal \sEEADC_freqZ0Z_2\ : std_logic;
signal \sCounterADCZ0Z_3\ : std_logic;
signal \un11_sacqtime_NE_3\ : std_logic;
signal \un11_sacqtime_NE_0_0_cascade_\ : std_logic;
signal \un11_sacqtime_NE_0\ : std_logic;
signal spi_data_mosi_3 : std_logic;
signal \sEEADC_freqZ0Z_3\ : std_logic;
signal \sCounterADCZ0Z_1\ : std_logic;
signal \sCounterADCZ0Z_0\ : std_logic;
signal \un11_sacqtime_NE_1\ : std_logic;
signal spi_data_mosi_0 : std_logic;
signal \sEEADC_freqZ0Z_0\ : std_logic;
signal \sEEADC_freqZ0Z_1\ : std_logic;
signal \sCounterADCZ0Z_7\ : std_logic;
signal \sCounterADCZ0Z_6\ : std_logic;
signal \un11_sacqtime_NE_2\ : std_logic;
signal \ADC7_c\ : std_logic;
signal \RAM_DATA_1Z0Z_8\ : std_logic;
signal \ADC8_c\ : std_logic;
signal \RAM_DATA_1Z0Z_9\ : std_logic;
signal top_tour2_c : std_logic;
signal \RAM_DATA_1Z0Z_12\ : std_logic;
signal spi_miso_ft_c : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_8\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8\ : std_logic;
signal \sDAC_spi_startZ0\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_\ : std_logic;
signal spi_select_c : std_logic;
signal spi_cs_ft_c : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_\ : std_logic;
signal spi_cs_rpi_c : std_logic;
signal \spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1\ : std_logic;
signal \spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3\ : std_logic;
signal \spi_slave_inst.N_1393_cascade_\ : std_logic;
signal spi_miso : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_0\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0_cascade_\ : std_logic;
signal \spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2\ : std_logic;
signal \spi_slave_inst.N_1396\ : std_logic;
signal \N_23_mux_cascade_\ : std_logic;
signal \N_25_mux_cascade_\ : std_logic;
signal m15_1 : std_logic;
signal op_eq_scounterdac10 : std_logic;
signal m8_2 : std_logic;
signal \N_23_mux\ : std_logic;
signal \N_30_mux_cascade_\ : std_logic;
signal \N_25_mux\ : std_logic;
signal \N_32_mux\ : std_logic;
signal \sCounterDACZ0Z_0\ : std_logic;
signal \sCounterDACZ0Z_1\ : std_logic;
signal \bfn_20_10_0_\ : std_logic;
signal \sCounterDACZ0Z_2\ : std_logic;
signal un2_scounterdac_cry_1 : std_logic;
signal \sCounterDACZ0Z_3\ : std_logic;
signal un2_scounterdac_cry_2 : std_logic;
signal \sCounterDACZ0Z_4\ : std_logic;
signal un2_scounterdac_cry_3 : std_logic;
signal \sCounterDACZ0Z_5\ : std_logic;
signal un2_scounterdac_cry_4 : std_logic;
signal \sCounterDACZ0Z_6\ : std_logic;
signal \un2_scounterdac_cry_5_THRU_CO\ : std_logic;
signal un2_scounterdac_cry_5 : std_logic;
signal \sCounterDACZ0Z_7\ : std_logic;
signal un2_scounterdac_cry_6 : std_logic;
signal \N_30_mux\ : std_logic;
signal \sCounterDACZ0Z_8\ : std_logic;
signal un2_scounterdac_cry_7 : std_logic;
signal un2_scounterdac_cry_8 : std_logic;
signal \bfn_20_11_0_\ : std_logic;
signal \sCounterDACZ0Z_9\ : std_logic;
signal pll_clk64_0_g : std_logic;
signal \spi_slave_inst.un23_i_ssn_3\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.rx_done_pos_sclk_iZ0\ : std_logic;
signal spi_sclk_g : std_logic;
signal \spi_slave_inst.spi_cs_iZ0\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_7\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_7\ : std_logic;
signal spi_data_mosi_6 : std_logic;
signal \sEEADC_freqZ0Z_6\ : std_logic;
signal spi_data_mosi_7 : std_logic;
signal \sEEADC_freqZ0Z_7\ : std_logic;
signal \sEEADC_freq_1_sqmuxa\ : std_logic;
signal \N_71\ : std_logic;
signal \LED3_c\ : std_logic;
signal \un4_sacqtime_cry_23_c_RNITTSZ0Z3\ : std_logic;
signal \RAM_DATA_cl_5Z0Z_15\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0\ : std_logic;
signal \bfn_22_7_0_\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1\ : std_logic;
signal \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2\ : std_logic;
signal \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3\ : std_logic;
signal \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5\ : std_logic;
signal \spi_slave_inst.spi_csZ0\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_i6\ : std_logic;
signal \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\ : std_logic;
signal \spi_slave_inst.tx_done_neg_sclk_iZ0\ : std_logic;
signal \spi_slave_inst.tx_done_reg1_iZ0\ : std_logic;
signal \spi_slave_inst.tx_done_reg3_iZ0\ : std_logic;
signal \spi_slave_inst.tx_done_reg2_iZ0\ : std_logic;
signal \spi_slave_inst.un4_tx_done_reg2_i\ : std_logic;
signal spi_data_mosi_1 : std_logic;
signal \sDAC_mem_25Z0Z_1\ : std_logic;
signal \sDAC_mem_25_1_sqmuxa\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \RAM_DATA_1Z0Z_15\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal pll_clk128_g : std_logic;
signal \N_31_i\ : std_logic;
signal \LED3_c_i_g\ : std_logic;

signal \RAM_ADD_wire\ : std_logic_vector(18 downto 0);
signal spi_mosi_rpi_wire : std_logic;
signal spi_sclk_rpi_wire : std_logic;
signal spi_miso_ft_wire : std_logic;
signal \ADC5_wire\ : std_logic;
signal \LED_ACQ_wire\ : std_logic;
signal reset_rpi_wire : std_logic;
signal trig_rpi_wire : std_logic;
signal \ADC2_wire\ : std_logic;
signal \DAC_mosi_wire\ : std_logic;
signal \RAM_nWE_wire\ : std_logic;
signal \ADC0_wire\ : std_logic;
signal \RAM_nLB_wire\ : std_logic;
signal spi_select_wire : std_logic;
signal \RAM_nCE_wire\ : std_logic;
signal spi_sclk_flash_wire : std_logic;
signal \ADC3_wire\ : std_logic;
signal pon_wire : std_logic;
signal \DAC_sclk_wire\ : std_logic;
signal \ADC1_wire\ : std_logic;
signal spi_cs_flash_wire : std_logic;
signal trig_ext_wire : std_logic;
signal top_tour1_wire : std_logic;
signal \LED_MODE_wire\ : std_logic;
signal \RAM_nUB_wire\ : std_logic;
signal \DAC_cs_wire\ : std_logic;
signal \ADC8_wire\ : std_logic;
signal \ADC_clk_wire\ : std_logic;
signal spi_miso_rpi_wire : std_logic;
signal poff_wire : std_logic;
signal \ADC4_wire\ : std_logic;
signal \ADC6_wire\ : std_logic;
signal \ADC7_wire\ : std_logic;
signal button_mode_wire : std_logic;
signal spi_sclk_ft_wire : std_logic;
signal trig_ft_wire : std_logic;
signal \ADC9_wire\ : std_logic;
signal cs_rpi2flash_wire : std_logic;
signal \LED3_wire\ : std_logic;
signal spi_mosi_ft_wire : std_logic;
signal \RAM_nOE_wire\ : std_logic;
signal clk_wire : std_logic;
signal top_tour2_wire : std_logic;
signal spi_cs_rpi_wire : std_logic;
signal spi_cs_ft_wire : std_logic;
signal spi_mosi_flash_wire : std_logic;
signal \pll128M2_inst.pll128M2_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    RAM_ADD <= \RAM_ADD_wire\;
    spi_mosi_rpi_wire <= spi_mosi_rpi;
    spi_sclk_rpi_wire <= spi_sclk_rpi;
    spi_miso_ft <= spi_miso_ft_wire;
    \ADC5_wire\ <= ADC5;
    LED_ACQ <= \LED_ACQ_wire\;
    reset_rpi_wire <= reset_rpi;
    trig_rpi_wire <= trig_rpi;
    \ADC2_wire\ <= ADC2;
    DAC_mosi <= \DAC_mosi_wire\;
    RAM_nWE <= \RAM_nWE_wire\;
    \ADC0_wire\ <= ADC0;
    RAM_nLB <= \RAM_nLB_wire\;
    spi_select_wire <= spi_select;
    RAM_nCE <= \RAM_nCE_wire\;
    spi_sclk_flash <= spi_sclk_flash_wire;
    \ADC3_wire\ <= ADC3;
    pon <= pon_wire;
    DAC_sclk <= \DAC_sclk_wire\;
    \ADC1_wire\ <= ADC1;
    spi_cs_flash <= spi_cs_flash_wire;
    trig_ext_wire <= trig_ext;
    top_tour1_wire <= top_tour1;
    LED_MODE <= \LED_MODE_wire\;
    RAM_nUB <= \RAM_nUB_wire\;
    DAC_cs <= \DAC_cs_wire\;
    \ADC8_wire\ <= ADC8;
    ADC_clk <= \ADC_clk_wire\;
    spi_miso_rpi <= spi_miso_rpi_wire;
    poff <= poff_wire;
    \ADC4_wire\ <= ADC4;
    \ADC6_wire\ <= ADC6;
    \ADC7_wire\ <= ADC7;
    button_mode_wire <= button_mode;
    spi_sclk_ft_wire <= spi_sclk_ft;
    trig_ft_wire <= trig_ft;
    \ADC9_wire\ <= ADC9;
    cs_rpi2flash_wire <= cs_rpi2flash;
    LED3 <= \LED3_wire\;
    spi_mosi_ft_wire <= spi_mosi_ft;
    RAM_nOE <= \RAM_nOE_wire\;
    clk_wire <= clk;
    top_tour2_wire <= top_tour2;
    spi_cs_rpi_wire <= spi_cs_rpi;
    spi_cs_ft_wire <= spi_cs_ft;
    spi_mosi_flash <= spi_mosi_flash_wire;
    \pll128M2_inst.pll128M2_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll128M2_inst.pll128M2_inst\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1010100",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \pll128M2_inst.pll_clk64_0\,
            REFERENCECLK => \N__20270\,
            RESETB => \N__49049\,
            BYPASS => \GNDG0\,
            PLLOUTCOREA => \pll128M2_inst.pll_clk128\,
            SDI => \GNDG0\,
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll128M2_inst.pll128M2_inst_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => \GNDG0\,
            PLLOUTGLOBALA => OPEN,
            SCLK => \GNDG0\
        );

    \RAM_ADD_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53520\,
            DIN => \N__53519\,
            DOUT => \N__53518\,
            PACKAGEPIN => \RAM_ADD_wire\(5)
        );

    \RAM_ADD_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53520\,
            PADOUT => \N__53519\,
            PADIN => \N__53518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35216\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_mosi_rpi_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53511\,
            DIN => \N__53510\,
            DOUT => \N__53509\,
            PACKAGEPIN => spi_mosi_rpi_wire
        );

    \spi_mosi_rpi_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53511\,
            PADOUT => \N__53510\,
            PADIN => \N__53509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_mosi_rpi_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_sclk_rpi_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53502\,
            DIN => \N__53501\,
            DOUT => \N__53500\,
            PACKAGEPIN => spi_sclk_rpi_wire
        );

    \spi_sclk_rpi_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53502\,
            PADOUT => \N__53501\,
            PADIN => \N__53500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_sclk_rpi_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_miso_ft_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53493\,
            DIN => \N__53492\,
            DOUT => \N__53491\,
            PACKAGEPIN => spi_miso_ft_wire
        );

    \spi_miso_ft_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53493\,
            PADOUT => \N__53492\,
            PADIN => \N__53491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__47600\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC5_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53484\,
            DIN => \N__53483\,
            DOUT => \N__53482\,
            PACKAGEPIN => \ADC5_wire\
        );

    \ADC5_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53484\,
            PADOUT => \N__53483\,
            PADIN => \N__53482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC5_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_ACQ_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53475\,
            DIN => \N__53474\,
            DOUT => \N__53473\,
            PACKAGEPIN => \LED_ACQ_wire\
        );

    \LED_ACQ_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53475\,
            PADOUT => \N__53474\,
            PADIN => \N__53473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23318\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \reset_rpi_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53466\,
            DIN => \N__53465\,
            DOUT => \N__53464\,
            PACKAGEPIN => reset_rpi_wire
        );

    \reset_rpi_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53466\,
            PADOUT => \N__53465\,
            PADIN => \N__53464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \LED3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53457\,
            DIN => \N__53456\,
            DOUT => \N__53455\,
            PACKAGEPIN => RAM_DATA(6)
        );

    \RAM_DATA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53457\,
            PADOUT => \N__53456\,
            PADIN => \N__53455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__43172\,
            DIN0 => \RAM_DATA_in_6\,
            DOUT0 => \N__26861\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53448\,
            DIN => \N__53447\,
            DOUT => \N__53446\,
            PACKAGEPIN => \RAM_ADD_wire\(9)
        );

    \RAM_ADD_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53448\,
            PADOUT => \N__53447\,
            PADIN => \N__53446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36218\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53439\,
            DIN => \N__53438\,
            DOUT => \N__53437\,
            PACKAGEPIN => RAM_DATA(11)
        );

    \RAM_DATA_iobuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53439\,
            PADOUT => \N__53438\,
            PADIN => \N__53437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__39428\,
            DIN0 => \RAM_DATA_in_11\,
            DOUT0 => \N__26594\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \trig_rpi_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53430\,
            DIN => \N__53429\,
            DOUT => \N__53428\,
            PACKAGEPIN => trig_rpi_wire
        );

    \trig_rpi_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53430\,
            PADOUT => \N__53429\,
            PADIN => \N__53428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => trig_rpi_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53421\,
            DIN => \N__53420\,
            DOUT => \N__53419\,
            PACKAGEPIN => RAM_DATA(0)
        );

    \RAM_DATA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53421\,
            PADOUT => \N__53420\,
            PADIN => \N__53419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__39071\,
            DIN0 => \RAM_DATA_in_0\,
            DOUT0 => \N__26822\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53412\,
            DIN => \N__53411\,
            DOUT => \N__53410\,
            PACKAGEPIN => \ADC2_wire\
        );

    \ADC2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53412\,
            PADOUT => \N__53411\,
            PADIN => \N__53410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC2_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53403\,
            DIN => \N__53402\,
            DOUT => \N__53401\,
            PACKAGEPIN => \RAM_ADD_wire\(18)
        );

    \RAM_ADD_obuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53403\,
            PADOUT => \N__53402\,
            PADIN => \N__53401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36290\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53394\,
            DIN => \N__53393\,
            DOUT => \N__53392\,
            PACKAGEPIN => \RAM_ADD_wire\(2)
        );

    \RAM_ADD_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53394\,
            PADOUT => \N__53393\,
            PADIN => \N__53392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36089\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DAC_mosi_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53385\,
            DIN => \N__53384\,
            DOUT => \N__53383\,
            PACKAGEPIN => \DAC_mosi_wire\
        );

    \DAC_mosi_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53385\,
            PADOUT => \N__53384\,
            PADIN => \N__53383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20810\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53376\,
            DIN => \N__53375\,
            DOUT => \N__53374\,
            PACKAGEPIN => \RAM_ADD_wire\(13)
        );

    \RAM_ADD_obuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53376\,
            PADOUT => \N__53375\,
            PADIN => \N__53374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35594\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_nWE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53367\,
            DIN => \N__53366\,
            DOUT => \N__53365\,
            PACKAGEPIN => \RAM_nWE_wire\
        );

    \RAM_nWE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53367\,
            PADOUT => \N__53366\,
            PADIN => \N__53365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33671\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53358\,
            DIN => \N__53357\,
            DOUT => \N__53356\,
            PACKAGEPIN => RAM_DATA(7)
        );

    \RAM_DATA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53358\,
            PADOUT => \N__53357\,
            PADIN => \N__53356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__39755\,
            DIN0 => \RAM_DATA_in_7\,
            DOUT0 => \N__39701\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC0_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53349\,
            DIN => \N__53348\,
            DOUT => \N__53347\,
            PACKAGEPIN => \ADC0_wire\
        );

    \ADC0_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53349\,
            PADOUT => \N__53348\,
            PADIN => \N__53347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC0_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_nLB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53340\,
            DIN => \N__53339\,
            DOUT => \N__53338\,
            PACKAGEPIN => \RAM_nLB_wire\
        );

    \RAM_nLB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53340\,
            PADOUT => \N__53339\,
            PADIN => \N__53338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53331\,
            DIN => \N__53330\,
            DOUT => \N__53329\,
            PACKAGEPIN => RAM_DATA(10)
        );

    \RAM_DATA_iobuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53331\,
            PADOUT => \N__53330\,
            PADIN => \N__53329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__39461\,
            DIN0 => \RAM_DATA_in_10\,
            DOUT0 => \N__26627\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53322\,
            DIN => \N__53321\,
            DOUT => \N__53320\,
            PACKAGEPIN => RAM_DATA(1)
        );

    \RAM_DATA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53322\,
            PADOUT => \N__53321\,
            PADIN => \N__53320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__44015\,
            DIN0 => \RAM_DATA_in_1\,
            DOUT0 => \N__26660\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_select_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53313\,
            DIN => \N__53312\,
            DOUT => \N__53311\,
            PACKAGEPIN => spi_select_wire
        );

    \spi_select_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53313\,
            PADOUT => \N__53312\,
            PADIN => \N__53311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_select_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_nCE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53304\,
            DIN => \N__53303\,
            DOUT => \N__53302\,
            PACKAGEPIN => \RAM_nCE_wire\
        );

    \RAM_nCE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53304\,
            PADOUT => \N__53303\,
            PADIN => \N__53302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_sclk_flash_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53295\,
            DIN => \N__53294\,
            DOUT => \N__53293\,
            PACKAGEPIN => spi_sclk_flash_wire
        );

    \spi_sclk_flash_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53295\,
            PADOUT => \N__53294\,
            PADIN => \N__53293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53286\,
            DIN => \N__53285\,
            DOUT => \N__53284\,
            PACKAGEPIN => \RAM_ADD_wire\(3)
        );

    \RAM_ADD_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53286\,
            PADOUT => \N__53285\,
            PADIN => \N__53284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__43244\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53277\,
            DIN => \N__53276\,
            DOUT => \N__53275\,
            PACKAGEPIN => \RAM_ADD_wire\(12)
        );

    \RAM_ADD_obuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53277\,
            PADOUT => \N__53276\,
            PADIN => \N__53275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35660\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53268\,
            DIN => \N__53267\,
            DOUT => \N__53266\,
            PACKAGEPIN => \ADC3_wire\
        );

    \ADC3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53268\,
            PADOUT => \N__53267\,
            PADIN => \N__53266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53259\,
            DIN => \N__53258\,
            DOUT => \N__53257\,
            PACKAGEPIN => RAM_DATA(15)
        );

    \RAM_DATA_iobuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53259\,
            PADOUT => \N__53258\,
            PADIN => \N__53257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__43142\,
            DIN0 => \RAM_DATA_in_15\,
            DOUT0 => \N__52367\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pon_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53250\,
            DIN => \N__53249\,
            DOUT => \N__53248\,
            PACKAGEPIN => pon_wire
        );

    \pon_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53250\,
            PADOUT => \N__53249\,
            PADIN => \N__53248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24014\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DAC_sclk_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53241\,
            DIN => \N__53240\,
            DOUT => \N__53239\,
            PACKAGEPIN => \DAC_sclk_wire\
        );

    \DAC_sclk_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53241\,
            PADOUT => \N__53240\,
            PADIN => \N__53239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20888\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53232\,
            DIN => \N__53231\,
            DOUT => \N__53230\,
            PACKAGEPIN => RAM_DATA(4)
        );

    \RAM_DATA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53232\,
            PADOUT => \N__53231\,
            PADIN => \N__53230\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__39785\,
            DIN0 => \RAM_DATA_in_4\,
            DOUT0 => \N__35930\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53223\,
            DIN => \N__53222\,
            DOUT => \N__53221\,
            PACKAGEPIN => \ADC1_wire\
        );

    \ADC1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53223\,
            PADOUT => \N__53222\,
            PADIN => \N__53221\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_cs_flash_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53214\,
            DIN => \N__53213\,
            DOUT => \N__53212\,
            PACKAGEPIN => spi_cs_flash_wire
        );

    \spi_cs_flash_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53214\,
            PADOUT => \N__53213\,
            PADIN => \N__53212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \trig_ext_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53205\,
            DIN => \N__53204\,
            DOUT => \N__53203\,
            PACKAGEPIN => trig_ext_wire
        );

    \trig_ext_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53205\,
            PADOUT => \N__53204\,
            PADIN => \N__53203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => trig_ext_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53196\,
            DIN => \N__53195\,
            DOUT => \N__53194\,
            PACKAGEPIN => \RAM_ADD_wire\(6)
        );

    \RAM_ADD_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53196\,
            PADOUT => \N__53195\,
            PADIN => \N__53194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35972\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \top_tour1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53187\,
            DIN => \N__53186\,
            DOUT => \N__53185\,
            PACKAGEPIN => top_tour1_wire
        );

    \top_tour1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53187\,
            PADOUT => \N__53186\,
            PADIN => \N__53185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => top_tour1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53178\,
            DIN => \N__53177\,
            DOUT => \N__53176\,
            PACKAGEPIN => \RAM_ADD_wire\(17)
        );

    \RAM_ADD_obuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53178\,
            PADOUT => \N__53177\,
            PADIN => \N__53176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36356\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53169\,
            DIN => \N__53168\,
            DOUT => \N__53167\,
            PACKAGEPIN => \RAM_ADD_wire\(0)
        );

    \RAM_ADD_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53169\,
            PADOUT => \N__53168\,
            PADIN => \N__53167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35861\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_MODE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53160\,
            DIN => \N__53159\,
            DOUT => \N__53158\,
            PACKAGEPIN => \LED_MODE_wire\
        );

    \LED_MODE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53160\,
            PADOUT => \N__53159\,
            PADIN => \N__53158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23618\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_nUB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53151\,
            DIN => \N__53150\,
            DOUT => \N__53149\,
            PACKAGEPIN => \RAM_nUB_wire\
        );

    \RAM_nUB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53151\,
            PADOUT => \N__53150\,
            PADIN => \N__53149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53142\,
            DIN => \N__53141\,
            DOUT => \N__53140\,
            PACKAGEPIN => \RAM_ADD_wire\(11)
        );

    \RAM_ADD_obuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53142\,
            PADOUT => \N__53141\,
            PADIN => \N__53140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35726\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53133\,
            DIN => \N__53132\,
            DOUT => \N__53131\,
            PACKAGEPIN => RAM_DATA(14)
        );

    \RAM_DATA_iobuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53133\,
            PADOUT => \N__53132\,
            PADIN => \N__53131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__43988\,
            DIN0 => \RAM_DATA_in_14\,
            DOUT0 => \N__26933\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DAC_cs_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53124\,
            DIN => \N__53123\,
            DOUT => \N__53122\,
            PACKAGEPIN => \DAC_cs_wire\
        );

    \DAC_cs_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53124\,
            PADOUT => \N__53123\,
            PADIN => \N__53122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20471\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC8_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53115\,
            DIN => \N__53114\,
            DOUT => \N__53113\,
            PACKAGEPIN => \ADC8_wire\
        );

    \ADC8_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53115\,
            PADOUT => \N__53114\,
            PADIN => \N__53113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC8_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53106\,
            DIN => \N__53105\,
            DOUT => \N__53104\,
            PACKAGEPIN => RAM_DATA(5)
        );

    \RAM_DATA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53106\,
            PADOUT => \N__53105\,
            PADIN => \N__53104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__43190\,
            DIN0 => \RAM_DATA_in_5\,
            DOUT0 => \N__26702\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC_clk_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53097\,
            DIN => \N__53096\,
            DOUT => \N__53095\,
            PACKAGEPIN => \ADC_clk_wire\
        );

    \ADC_clk_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53097\,
            PADOUT => \N__53096\,
            PADIN => \N__53095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34028\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_miso_rpi_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53088\,
            DIN => \N__53087\,
            DOUT => \N__53086\,
            PACKAGEPIN => spi_miso_rpi_wire
        );

    \spi_miso_rpi_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53088\,
            PADOUT => \N__53087\,
            PADIN => \N__53086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__20294\,
            DIN0 => OPEN,
            DOUT0 => \N__47798\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53079\,
            DIN => \N__53078\,
            DOUT => \N__53077\,
            PACKAGEPIN => \RAM_ADD_wire\(7)
        );

    \RAM_ADD_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53079\,
            PADOUT => \N__53078\,
            PADIN => \N__53077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36152\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \poff_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53070\,
            DIN => \N__53069\,
            DOUT => \N__53068\,
            PACKAGEPIN => poff_wire
        );

    \poff_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53070\,
            PADOUT => \N__53069\,
            PADIN => \N__53068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__26423\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC4_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53061\,
            DIN => \N__53060\,
            DOUT => \N__53059\,
            PACKAGEPIN => \ADC4_wire\
        );

    \ADC4_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53061\,
            PADOUT => \N__53060\,
            PADIN => \N__53059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC4_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC6_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53052\,
            DIN => \N__53051\,
            DOUT => \N__53050\,
            PACKAGEPIN => \ADC6_wire\
        );

    \ADC6_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53052\,
            PADOUT => \N__53051\,
            PADIN => \N__53050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC6_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53043\,
            DIN => \N__53042\,
            DOUT => \N__53041\,
            PACKAGEPIN => \RAM_ADD_wire\(16)
        );

    \RAM_ADD_obuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53043\,
            PADOUT => \N__53042\,
            PADIN => \N__53041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35381\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53034\,
            DIN => \N__53033\,
            DOUT => \N__53032\,
            PACKAGEPIN => \RAM_ADD_wire\(1)
        );

    \RAM_ADD_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53034\,
            PADOUT => \N__53033\,
            PADIN => \N__53032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__36029\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC7_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53025\,
            DIN => \N__53024\,
            DOUT => \N__53023\,
            PACKAGEPIN => \ADC7_wire\
        );

    \ADC7_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53025\,
            PADOUT => \N__53024\,
            PADIN => \N__53023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC7_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \button_mode_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53016\,
            DIN => \N__53015\,
            DOUT => \N__53014\,
            PACKAGEPIN => button_mode_wire
        );

    \button_mode_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53016\,
            PADOUT => \N__53015\,
            PADIN => \N__53014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => button_mode_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_sclk_ft_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53007\,
            DIN => \N__53006\,
            DOUT => \N__53005\,
            PACKAGEPIN => spi_sclk_ft_wire
        );

    \spi_sclk_ft_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53007\,
            PADOUT => \N__53006\,
            PADIN => \N__53005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_sclk_ft_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52998\,
            DIN => \N__52997\,
            DOUT => \N__52996\,
            PACKAGEPIN => RAM_DATA(8)
        );

    \RAM_DATA_iobuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__52998\,
            PADOUT => \N__52997\,
            PADIN => \N__52996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__39101\,
            DIN0 => \RAM_DATA_in_8\,
            DOUT0 => \N__47702\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52989\,
            DIN => \N__52988\,
            DOUT => \N__52987\,
            PACKAGEPIN => \RAM_ADD_wire\(10)
        );

    \RAM_ADD_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__52989\,
            PADOUT => \N__52988\,
            PADIN => \N__52987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35798\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52980\,
            DIN => \N__52979\,
            DOUT => \N__52978\,
            PACKAGEPIN => RAM_DATA(13)
        );

    \RAM_DATA_iobuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__52980\,
            PADOUT => \N__52979\,
            PADIN => \N__52978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__48815\,
            DIN0 => \RAM_DATA_in_13\,
            DOUT0 => \N__26546\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \trig_ft_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52971\,
            DIN => \N__52970\,
            DOUT => \N__52969\,
            PACKAGEPIN => trig_ft_wire
        );

    \trig_ft_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52971\,
            PADOUT => \N__52970\,
            PADIN => \N__52969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => trig_ft_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC9_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52962\,
            DIN => \N__52961\,
            DOUT => \N__52960\,
            PACKAGEPIN => \ADC9_wire\
        );

    \ADC9_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52962\,
            PADOUT => \N__52961\,
            PADIN => \N__52960\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC9_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52953\,
            DIN => \N__52952\,
            DOUT => \N__52951\,
            PACKAGEPIN => RAM_DATA(2)
        );

    \RAM_DATA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__52953\,
            PADOUT => \N__52952\,
            PADIN => \N__52951\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__39725\,
            DIN0 => \RAM_DATA_in_2\,
            DOUT0 => \N__26894\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \cs_rpi2flash_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52944\,
            DIN => \N__52943\,
            DOUT => \N__52942\,
            PACKAGEPIN => cs_rpi2flash_wire
        );

    \cs_rpi2flash_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52944\,
            PADOUT => \N__52943\,
            PADIN => \N__52942\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => cs_rpi2flash_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52935\,
            DIN => \N__52934\,
            DOUT => \N__52933\,
            PACKAGEPIN => \LED3_wire\
        );

    \LED3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__52935\,
            PADOUT => \N__52934\,
            PADIN => \N__52933\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__49419\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_mosi_ft_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52926\,
            DIN => \N__52925\,
            DOUT => \N__52924\,
            PACKAGEPIN => spi_mosi_ft_wire
        );

    \spi_mosi_ft_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52926\,
            PADOUT => \N__52925\,
            PADIN => \N__52924\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_mosi_ft_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_nOE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52917\,
            DIN => \N__52916\,
            DOUT => \N__52915\,
            PACKAGEPIN => \RAM_nOE_wire\
        );

    \RAM_nOE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__52917\,
            PADOUT => \N__52916\,
            PADIN => \N__52915\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52908\,
            DIN => \N__52907\,
            DOUT => \N__52906\,
            PACKAGEPIN => \RAM_ADD_wire\(4)
        );

    \RAM_ADD_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__52908\,
            PADOUT => \N__52907\,
            PADIN => \N__52906\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__43538\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52899\,
            DIN => \N__52898\,
            DOUT => \N__52897\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52899\,
            PADOUT => \N__52898\,
            PADIN => \N__52897\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \top_tour2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52890\,
            DIN => \N__52889\,
            DOUT => \N__52888\,
            PACKAGEPIN => top_tour2_wire
        );

    \top_tour2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52890\,
            PADOUT => \N__52889\,
            PADIN => \N__52888\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => top_tour2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_cs_rpi_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52881\,
            DIN => \N__52880\,
            DOUT => \N__52879\,
            PACKAGEPIN => spi_cs_rpi_wire
        );

    \spi_cs_rpi_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52881\,
            PADOUT => \N__52880\,
            PADIN => \N__52879\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_cs_rpi_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52872\,
            DIN => \N__52871\,
            DOUT => \N__52870\,
            PACKAGEPIN => \RAM_ADD_wire\(15)
        );

    \RAM_ADD_obuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__52872\,
            PADOUT => \N__52871\,
            PADIN => \N__52870\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35453\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52863\,
            DIN => \N__52862\,
            DOUT => \N__52861\,
            PACKAGEPIN => RAM_DATA(9)
        );

    \RAM_DATA_iobuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__52863\,
            PADOUT => \N__52862\,
            PADIN => \N__52861\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__43115\,
            DIN0 => \RAM_DATA_in_9\,
            DOUT0 => \N__47657\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52854\,
            DIN => \N__52853\,
            DOUT => \N__52852\,
            PACKAGEPIN => \RAM_ADD_wire\(8)
        );

    \RAM_ADD_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__52854\,
            PADOUT => \N__52853\,
            PADIN => \N__52852\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__43610\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52845\,
            DIN => \N__52844\,
            DOUT => \N__52843\,
            PACKAGEPIN => RAM_DATA(12)
        );

    \RAM_DATA_iobuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__52845\,
            PADOUT => \N__52844\,
            PADIN => \N__52843\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__44075\,
            DIN0 => \RAM_DATA_in_12\,
            DOUT0 => \N__47618\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52836\,
            DIN => \N__52835\,
            DOUT => \N__52834\,
            PACKAGEPIN => RAM_DATA(3)
        );

    \RAM_DATA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__52836\,
            PADOUT => \N__52835\,
            PADIN => \N__52834\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__44045\,
            DIN0 => \RAM_DATA_in_3\,
            DOUT0 => \N__33944\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_cs_ft_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52827\,
            DIN => \N__52826\,
            DOUT => \N__52825\,
            PACKAGEPIN => spi_cs_ft_wire
        );

    \spi_cs_ft_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__52827\,
            PADOUT => \N__52826\,
            PADIN => \N__52825\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_cs_ft_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_mosi_flash_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52818\,
            DIN => \N__52817\,
            DOUT => \N__52816\,
            PACKAGEPIN => spi_mosi_flash_wire
        );

    \spi_mosi_flash_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__52818\,
            PADOUT => \N__52817\,
            PADIN => \N__52816\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__52809\,
            DIN => \N__52808\,
            DOUT => \N__52807\,
            PACKAGEPIN => \RAM_ADD_wire\(14)
        );

    \RAM_ADD_obuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__52809\,
            PADOUT => \N__52808\,
            PADIN => \N__52807\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35528\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__12567\ : InMux
    port map (
            O => \N__52790\,
            I => \N__52770\
        );

    \I__12566\ : InMux
    port map (
            O => \N__52789\,
            I => \N__52770\
        );

    \I__12565\ : InMux
    port map (
            O => \N__52788\,
            I => \N__52770\
        );

    \I__12564\ : InMux
    port map (
            O => \N__52787\,
            I => \N__52770\
        );

    \I__12563\ : CascadeMux
    port map (
            O => \N__52786\,
            I => \N__52760\
        );

    \I__12562\ : CascadeMux
    port map (
            O => \N__52785\,
            I => \N__52756\
        );

    \I__12561\ : CascadeMux
    port map (
            O => \N__52784\,
            I => \N__52752\
        );

    \I__12560\ : CascadeMux
    port map (
            O => \N__52783\,
            I => \N__52748\
        );

    \I__12559\ : CascadeMux
    port map (
            O => \N__52782\,
            I => \N__52739\
        );

    \I__12558\ : InMux
    port map (
            O => \N__52781\,
            I => \N__52731\
        );

    \I__12557\ : InMux
    port map (
            O => \N__52780\,
            I => \N__52731\
        );

    \I__12556\ : InMux
    port map (
            O => \N__52779\,
            I => \N__52731\
        );

    \I__12555\ : LocalMux
    port map (
            O => \N__52770\,
            I => \N__52728\
        );

    \I__12554\ : InMux
    port map (
            O => \N__52769\,
            I => \N__52721\
        );

    \I__12553\ : InMux
    port map (
            O => \N__52768\,
            I => \N__52721\
        );

    \I__12552\ : InMux
    port map (
            O => \N__52767\,
            I => \N__52721\
        );

    \I__12551\ : InMux
    port map (
            O => \N__52766\,
            I => \N__52712\
        );

    \I__12550\ : InMux
    port map (
            O => \N__52765\,
            I => \N__52712\
        );

    \I__12549\ : InMux
    port map (
            O => \N__52764\,
            I => \N__52712\
        );

    \I__12548\ : InMux
    port map (
            O => \N__52763\,
            I => \N__52712\
        );

    \I__12547\ : InMux
    port map (
            O => \N__52760\,
            I => \N__52688\
        );

    \I__12546\ : InMux
    port map (
            O => \N__52759\,
            I => \N__52688\
        );

    \I__12545\ : InMux
    port map (
            O => \N__52756\,
            I => \N__52688\
        );

    \I__12544\ : InMux
    port map (
            O => \N__52755\,
            I => \N__52688\
        );

    \I__12543\ : InMux
    port map (
            O => \N__52752\,
            I => \N__52688\
        );

    \I__12542\ : InMux
    port map (
            O => \N__52751\,
            I => \N__52688\
        );

    \I__12541\ : InMux
    port map (
            O => \N__52748\,
            I => \N__52688\
        );

    \I__12540\ : InMux
    port map (
            O => \N__52747\,
            I => \N__52688\
        );

    \I__12539\ : CascadeMux
    port map (
            O => \N__52746\,
            I => \N__52685\
        );

    \I__12538\ : CascadeMux
    port map (
            O => \N__52745\,
            I => \N__52681\
        );

    \I__12537\ : CascadeMux
    port map (
            O => \N__52744\,
            I => \N__52677\
        );

    \I__12536\ : CascadeMux
    port map (
            O => \N__52743\,
            I => \N__52673\
        );

    \I__12535\ : InMux
    port map (
            O => \N__52742\,
            I => \N__52661\
        );

    \I__12534\ : InMux
    port map (
            O => \N__52739\,
            I => \N__52661\
        );

    \I__12533\ : InMux
    port map (
            O => \N__52738\,
            I => \N__52661\
        );

    \I__12532\ : LocalMux
    port map (
            O => \N__52731\,
            I => \N__52658\
        );

    \I__12531\ : Span4Mux_h
    port map (
            O => \N__52728\,
            I => \N__52651\
        );

    \I__12530\ : LocalMux
    port map (
            O => \N__52721\,
            I => \N__52651\
        );

    \I__12529\ : LocalMux
    port map (
            O => \N__52712\,
            I => \N__52651\
        );

    \I__12528\ : CascadeMux
    port map (
            O => \N__52711\,
            I => \N__52646\
        );

    \I__12527\ : CascadeMux
    port map (
            O => \N__52710\,
            I => \N__52643\
        );

    \I__12526\ : CascadeMux
    port map (
            O => \N__52709\,
            I => \N__52640\
        );

    \I__12525\ : CascadeMux
    port map (
            O => \N__52708\,
            I => \N__52636\
        );

    \I__12524\ : CascadeMux
    port map (
            O => \N__52707\,
            I => \N__52633\
        );

    \I__12523\ : CascadeMux
    port map (
            O => \N__52706\,
            I => \N__52630\
        );

    \I__12522\ : CascadeMux
    port map (
            O => \N__52705\,
            I => \N__52627\
        );

    \I__12521\ : LocalMux
    port map (
            O => \N__52688\,
            I => \N__52620\
        );

    \I__12520\ : InMux
    port map (
            O => \N__52685\,
            I => \N__52603\
        );

    \I__12519\ : InMux
    port map (
            O => \N__52684\,
            I => \N__52603\
        );

    \I__12518\ : InMux
    port map (
            O => \N__52681\,
            I => \N__52603\
        );

    \I__12517\ : InMux
    port map (
            O => \N__52680\,
            I => \N__52603\
        );

    \I__12516\ : InMux
    port map (
            O => \N__52677\,
            I => \N__52603\
        );

    \I__12515\ : InMux
    port map (
            O => \N__52676\,
            I => \N__52603\
        );

    \I__12514\ : InMux
    port map (
            O => \N__52673\,
            I => \N__52603\
        );

    \I__12513\ : InMux
    port map (
            O => \N__52672\,
            I => \N__52603\
        );

    \I__12512\ : CascadeMux
    port map (
            O => \N__52671\,
            I => \N__52599\
        );

    \I__12511\ : CascadeMux
    port map (
            O => \N__52670\,
            I => \N__52595\
        );

    \I__12510\ : CascadeMux
    port map (
            O => \N__52669\,
            I => \N__52591\
        );

    \I__12509\ : CascadeMux
    port map (
            O => \N__52668\,
            I => \N__52587\
        );

    \I__12508\ : LocalMux
    port map (
            O => \N__52661\,
            I => \N__52579\
        );

    \I__12507\ : Span4Mux_v
    port map (
            O => \N__52658\,
            I => \N__52579\
        );

    \I__12506\ : Span4Mux_v
    port map (
            O => \N__52651\,
            I => \N__52579\
        );

    \I__12505\ : InMux
    port map (
            O => \N__52650\,
            I => \N__52574\
        );

    \I__12504\ : InMux
    port map (
            O => \N__52649\,
            I => \N__52574\
        );

    \I__12503\ : InMux
    port map (
            O => \N__52646\,
            I => \N__52563\
        );

    \I__12502\ : InMux
    port map (
            O => \N__52643\,
            I => \N__52563\
        );

    \I__12501\ : InMux
    port map (
            O => \N__52640\,
            I => \N__52563\
        );

    \I__12500\ : InMux
    port map (
            O => \N__52639\,
            I => \N__52552\
        );

    \I__12499\ : InMux
    port map (
            O => \N__52636\,
            I => \N__52552\
        );

    \I__12498\ : InMux
    port map (
            O => \N__52633\,
            I => \N__52552\
        );

    \I__12497\ : InMux
    port map (
            O => \N__52630\,
            I => \N__52552\
        );

    \I__12496\ : InMux
    port map (
            O => \N__52627\,
            I => \N__52552\
        );

    \I__12495\ : CascadeMux
    port map (
            O => \N__52626\,
            I => \N__52549\
        );

    \I__12494\ : CascadeMux
    port map (
            O => \N__52625\,
            I => \N__52545\
        );

    \I__12493\ : CascadeMux
    port map (
            O => \N__52624\,
            I => \N__52541\
        );

    \I__12492\ : CascadeMux
    port map (
            O => \N__52623\,
            I => \N__52537\
        );

    \I__12491\ : Span4Mux_v
    port map (
            O => \N__52620\,
            I => \N__52531\
        );

    \I__12490\ : LocalMux
    port map (
            O => \N__52603\,
            I => \N__52531\
        );

    \I__12489\ : InMux
    port map (
            O => \N__52602\,
            I => \N__52514\
        );

    \I__12488\ : InMux
    port map (
            O => \N__52599\,
            I => \N__52514\
        );

    \I__12487\ : InMux
    port map (
            O => \N__52598\,
            I => \N__52514\
        );

    \I__12486\ : InMux
    port map (
            O => \N__52595\,
            I => \N__52514\
        );

    \I__12485\ : InMux
    port map (
            O => \N__52594\,
            I => \N__52514\
        );

    \I__12484\ : InMux
    port map (
            O => \N__52591\,
            I => \N__52514\
        );

    \I__12483\ : InMux
    port map (
            O => \N__52590\,
            I => \N__52514\
        );

    \I__12482\ : InMux
    port map (
            O => \N__52587\,
            I => \N__52514\
        );

    \I__12481\ : CascadeMux
    port map (
            O => \N__52586\,
            I => \N__52511\
        );

    \I__12480\ : Span4Mux_v
    port map (
            O => \N__52579\,
            I => \N__52507\
        );

    \I__12479\ : LocalMux
    port map (
            O => \N__52574\,
            I => \N__52504\
        );

    \I__12478\ : CascadeMux
    port map (
            O => \N__52573\,
            I => \N__52500\
        );

    \I__12477\ : CascadeMux
    port map (
            O => \N__52572\,
            I => \N__52496\
        );

    \I__12476\ : CascadeMux
    port map (
            O => \N__52571\,
            I => \N__52492\
        );

    \I__12475\ : CascadeMux
    port map (
            O => \N__52570\,
            I => \N__52488\
        );

    \I__12474\ : LocalMux
    port map (
            O => \N__52563\,
            I => \N__52485\
        );

    \I__12473\ : LocalMux
    port map (
            O => \N__52552\,
            I => \N__52482\
        );

    \I__12472\ : InMux
    port map (
            O => \N__52549\,
            I => \N__52465\
        );

    \I__12471\ : InMux
    port map (
            O => \N__52548\,
            I => \N__52465\
        );

    \I__12470\ : InMux
    port map (
            O => \N__52545\,
            I => \N__52465\
        );

    \I__12469\ : InMux
    port map (
            O => \N__52544\,
            I => \N__52465\
        );

    \I__12468\ : InMux
    port map (
            O => \N__52541\,
            I => \N__52465\
        );

    \I__12467\ : InMux
    port map (
            O => \N__52540\,
            I => \N__52465\
        );

    \I__12466\ : InMux
    port map (
            O => \N__52537\,
            I => \N__52465\
        );

    \I__12465\ : InMux
    port map (
            O => \N__52536\,
            I => \N__52465\
        );

    \I__12464\ : Span4Mux_h
    port map (
            O => \N__52531\,
            I => \N__52460\
        );

    \I__12463\ : LocalMux
    port map (
            O => \N__52514\,
            I => \N__52460\
        );

    \I__12462\ : InMux
    port map (
            O => \N__52511\,
            I => \N__52455\
        );

    \I__12461\ : InMux
    port map (
            O => \N__52510\,
            I => \N__52455\
        );

    \I__12460\ : Span4Mux_h
    port map (
            O => \N__52507\,
            I => \N__52450\
        );

    \I__12459\ : Span4Mux_v
    port map (
            O => \N__52504\,
            I => \N__52450\
        );

    \I__12458\ : InMux
    port map (
            O => \N__52503\,
            I => \N__52433\
        );

    \I__12457\ : InMux
    port map (
            O => \N__52500\,
            I => \N__52433\
        );

    \I__12456\ : InMux
    port map (
            O => \N__52499\,
            I => \N__52433\
        );

    \I__12455\ : InMux
    port map (
            O => \N__52496\,
            I => \N__52433\
        );

    \I__12454\ : InMux
    port map (
            O => \N__52495\,
            I => \N__52433\
        );

    \I__12453\ : InMux
    port map (
            O => \N__52492\,
            I => \N__52433\
        );

    \I__12452\ : InMux
    port map (
            O => \N__52491\,
            I => \N__52433\
        );

    \I__12451\ : InMux
    port map (
            O => \N__52488\,
            I => \N__52433\
        );

    \I__12450\ : Span4Mux_v
    port map (
            O => \N__52485\,
            I => \N__52428\
        );

    \I__12449\ : Span4Mux_v
    port map (
            O => \N__52482\,
            I => \N__52428\
        );

    \I__12448\ : LocalMux
    port map (
            O => \N__52465\,
            I => \N__52425\
        );

    \I__12447\ : Span4Mux_h
    port map (
            O => \N__52460\,
            I => \N__52420\
        );

    \I__12446\ : LocalMux
    port map (
            O => \N__52455\,
            I => \N__52420\
        );

    \I__12445\ : Span4Mux_h
    port map (
            O => \N__52450\,
            I => \N__52417\
        );

    \I__12444\ : LocalMux
    port map (
            O => \N__52433\,
            I => \N__52414\
        );

    \I__12443\ : Span4Mux_h
    port map (
            O => \N__52428\,
            I => \N__52409\
        );

    \I__12442\ : Span4Mux_v
    port map (
            O => \N__52425\,
            I => \N__52409\
        );

    \I__12441\ : Span4Mux_v
    port map (
            O => \N__52420\,
            I => \N__52405\
        );

    \I__12440\ : Span4Mux_h
    port map (
            O => \N__52417\,
            I => \N__52402\
        );

    \I__12439\ : Span4Mux_v
    port map (
            O => \N__52414\,
            I => \N__52399\
        );

    \I__12438\ : Span4Mux_h
    port map (
            O => \N__52409\,
            I => \N__52396\
        );

    \I__12437\ : InMux
    port map (
            O => \N__52408\,
            I => \N__52393\
        );

    \I__12436\ : Span4Mux_v
    port map (
            O => \N__52405\,
            I => \N__52390\
        );

    \I__12435\ : Span4Mux_v
    port map (
            O => \N__52402\,
            I => \N__52385\
        );

    \I__12434\ : Span4Mux_h
    port map (
            O => \N__52399\,
            I => \N__52385\
        );

    \I__12433\ : Span4Mux_h
    port map (
            O => \N__52396\,
            I => \N__52380\
        );

    \I__12432\ : LocalMux
    port map (
            O => \N__52393\,
            I => \N__52380\
        );

    \I__12431\ : Span4Mux_h
    port map (
            O => \N__52390\,
            I => \N__52377\
        );

    \I__12430\ : Span4Mux_h
    port map (
            O => \N__52385\,
            I => \N__52372\
        );

    \I__12429\ : Span4Mux_v
    port map (
            O => \N__52380\,
            I => \N__52372\
        );

    \I__12428\ : Odrv4
    port map (
            O => \N__52377\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12427\ : Odrv4
    port map (
            O => \N__52372\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12426\ : IoInMux
    port map (
            O => \N__52367\,
            I => \N__52364\
        );

    \I__12425\ : LocalMux
    port map (
            O => \N__52364\,
            I => \N__52361\
        );

    \I__12424\ : IoSpan4Mux
    port map (
            O => \N__52361\,
            I => \N__52358\
        );

    \I__12423\ : Span4Mux_s3_h
    port map (
            O => \N__52358\,
            I => \N__52355\
        );

    \I__12422\ : Span4Mux_v
    port map (
            O => \N__52355\,
            I => \N__52352\
        );

    \I__12421\ : Odrv4
    port map (
            O => \N__52352\,
            I => \RAM_DATA_1Z0Z_15\
        );

    \I__12420\ : ClkMux
    port map (
            O => \N__52349\,
            I => \N__51902\
        );

    \I__12419\ : ClkMux
    port map (
            O => \N__52348\,
            I => \N__51902\
        );

    \I__12418\ : ClkMux
    port map (
            O => \N__52347\,
            I => \N__51902\
        );

    \I__12417\ : ClkMux
    port map (
            O => \N__52346\,
            I => \N__51902\
        );

    \I__12416\ : ClkMux
    port map (
            O => \N__52345\,
            I => \N__51902\
        );

    \I__12415\ : ClkMux
    port map (
            O => \N__52344\,
            I => \N__51902\
        );

    \I__12414\ : ClkMux
    port map (
            O => \N__52343\,
            I => \N__51902\
        );

    \I__12413\ : ClkMux
    port map (
            O => \N__52342\,
            I => \N__51902\
        );

    \I__12412\ : ClkMux
    port map (
            O => \N__52341\,
            I => \N__51902\
        );

    \I__12411\ : ClkMux
    port map (
            O => \N__52340\,
            I => \N__51902\
        );

    \I__12410\ : ClkMux
    port map (
            O => \N__52339\,
            I => \N__51902\
        );

    \I__12409\ : ClkMux
    port map (
            O => \N__52338\,
            I => \N__51902\
        );

    \I__12408\ : ClkMux
    port map (
            O => \N__52337\,
            I => \N__51902\
        );

    \I__12407\ : ClkMux
    port map (
            O => \N__52336\,
            I => \N__51902\
        );

    \I__12406\ : ClkMux
    port map (
            O => \N__52335\,
            I => \N__51902\
        );

    \I__12405\ : ClkMux
    port map (
            O => \N__52334\,
            I => \N__51902\
        );

    \I__12404\ : ClkMux
    port map (
            O => \N__52333\,
            I => \N__51902\
        );

    \I__12403\ : ClkMux
    port map (
            O => \N__52332\,
            I => \N__51902\
        );

    \I__12402\ : ClkMux
    port map (
            O => \N__52331\,
            I => \N__51902\
        );

    \I__12401\ : ClkMux
    port map (
            O => \N__52330\,
            I => \N__51902\
        );

    \I__12400\ : ClkMux
    port map (
            O => \N__52329\,
            I => \N__51902\
        );

    \I__12399\ : ClkMux
    port map (
            O => \N__52328\,
            I => \N__51902\
        );

    \I__12398\ : ClkMux
    port map (
            O => \N__52327\,
            I => \N__51902\
        );

    \I__12397\ : ClkMux
    port map (
            O => \N__52326\,
            I => \N__51902\
        );

    \I__12396\ : ClkMux
    port map (
            O => \N__52325\,
            I => \N__51902\
        );

    \I__12395\ : ClkMux
    port map (
            O => \N__52324\,
            I => \N__51902\
        );

    \I__12394\ : ClkMux
    port map (
            O => \N__52323\,
            I => \N__51902\
        );

    \I__12393\ : ClkMux
    port map (
            O => \N__52322\,
            I => \N__51902\
        );

    \I__12392\ : ClkMux
    port map (
            O => \N__52321\,
            I => \N__51902\
        );

    \I__12391\ : ClkMux
    port map (
            O => \N__52320\,
            I => \N__51902\
        );

    \I__12390\ : ClkMux
    port map (
            O => \N__52319\,
            I => \N__51902\
        );

    \I__12389\ : ClkMux
    port map (
            O => \N__52318\,
            I => \N__51902\
        );

    \I__12388\ : ClkMux
    port map (
            O => \N__52317\,
            I => \N__51902\
        );

    \I__12387\ : ClkMux
    port map (
            O => \N__52316\,
            I => \N__51902\
        );

    \I__12386\ : ClkMux
    port map (
            O => \N__52315\,
            I => \N__51902\
        );

    \I__12385\ : ClkMux
    port map (
            O => \N__52314\,
            I => \N__51902\
        );

    \I__12384\ : ClkMux
    port map (
            O => \N__52313\,
            I => \N__51902\
        );

    \I__12383\ : ClkMux
    port map (
            O => \N__52312\,
            I => \N__51902\
        );

    \I__12382\ : ClkMux
    port map (
            O => \N__52311\,
            I => \N__51902\
        );

    \I__12381\ : ClkMux
    port map (
            O => \N__52310\,
            I => \N__51902\
        );

    \I__12380\ : ClkMux
    port map (
            O => \N__52309\,
            I => \N__51902\
        );

    \I__12379\ : ClkMux
    port map (
            O => \N__52308\,
            I => \N__51902\
        );

    \I__12378\ : ClkMux
    port map (
            O => \N__52307\,
            I => \N__51902\
        );

    \I__12377\ : ClkMux
    port map (
            O => \N__52306\,
            I => \N__51902\
        );

    \I__12376\ : ClkMux
    port map (
            O => \N__52305\,
            I => \N__51902\
        );

    \I__12375\ : ClkMux
    port map (
            O => \N__52304\,
            I => \N__51902\
        );

    \I__12374\ : ClkMux
    port map (
            O => \N__52303\,
            I => \N__51902\
        );

    \I__12373\ : ClkMux
    port map (
            O => \N__52302\,
            I => \N__51902\
        );

    \I__12372\ : ClkMux
    port map (
            O => \N__52301\,
            I => \N__51902\
        );

    \I__12371\ : ClkMux
    port map (
            O => \N__52300\,
            I => \N__51902\
        );

    \I__12370\ : ClkMux
    port map (
            O => \N__52299\,
            I => \N__51902\
        );

    \I__12369\ : ClkMux
    port map (
            O => \N__52298\,
            I => \N__51902\
        );

    \I__12368\ : ClkMux
    port map (
            O => \N__52297\,
            I => \N__51902\
        );

    \I__12367\ : ClkMux
    port map (
            O => \N__52296\,
            I => \N__51902\
        );

    \I__12366\ : ClkMux
    port map (
            O => \N__52295\,
            I => \N__51902\
        );

    \I__12365\ : ClkMux
    port map (
            O => \N__52294\,
            I => \N__51902\
        );

    \I__12364\ : ClkMux
    port map (
            O => \N__52293\,
            I => \N__51902\
        );

    \I__12363\ : ClkMux
    port map (
            O => \N__52292\,
            I => \N__51902\
        );

    \I__12362\ : ClkMux
    port map (
            O => \N__52291\,
            I => \N__51902\
        );

    \I__12361\ : ClkMux
    port map (
            O => \N__52290\,
            I => \N__51902\
        );

    \I__12360\ : ClkMux
    port map (
            O => \N__52289\,
            I => \N__51902\
        );

    \I__12359\ : ClkMux
    port map (
            O => \N__52288\,
            I => \N__51902\
        );

    \I__12358\ : ClkMux
    port map (
            O => \N__52287\,
            I => \N__51902\
        );

    \I__12357\ : ClkMux
    port map (
            O => \N__52286\,
            I => \N__51902\
        );

    \I__12356\ : ClkMux
    port map (
            O => \N__52285\,
            I => \N__51902\
        );

    \I__12355\ : ClkMux
    port map (
            O => \N__52284\,
            I => \N__51902\
        );

    \I__12354\ : ClkMux
    port map (
            O => \N__52283\,
            I => \N__51902\
        );

    \I__12353\ : ClkMux
    port map (
            O => \N__52282\,
            I => \N__51902\
        );

    \I__12352\ : ClkMux
    port map (
            O => \N__52281\,
            I => \N__51902\
        );

    \I__12351\ : ClkMux
    port map (
            O => \N__52280\,
            I => \N__51902\
        );

    \I__12350\ : ClkMux
    port map (
            O => \N__52279\,
            I => \N__51902\
        );

    \I__12349\ : ClkMux
    port map (
            O => \N__52278\,
            I => \N__51902\
        );

    \I__12348\ : ClkMux
    port map (
            O => \N__52277\,
            I => \N__51902\
        );

    \I__12347\ : ClkMux
    port map (
            O => \N__52276\,
            I => \N__51902\
        );

    \I__12346\ : ClkMux
    port map (
            O => \N__52275\,
            I => \N__51902\
        );

    \I__12345\ : ClkMux
    port map (
            O => \N__52274\,
            I => \N__51902\
        );

    \I__12344\ : ClkMux
    port map (
            O => \N__52273\,
            I => \N__51902\
        );

    \I__12343\ : ClkMux
    port map (
            O => \N__52272\,
            I => \N__51902\
        );

    \I__12342\ : ClkMux
    port map (
            O => \N__52271\,
            I => \N__51902\
        );

    \I__12341\ : ClkMux
    port map (
            O => \N__52270\,
            I => \N__51902\
        );

    \I__12340\ : ClkMux
    port map (
            O => \N__52269\,
            I => \N__51902\
        );

    \I__12339\ : ClkMux
    port map (
            O => \N__52268\,
            I => \N__51902\
        );

    \I__12338\ : ClkMux
    port map (
            O => \N__52267\,
            I => \N__51902\
        );

    \I__12337\ : ClkMux
    port map (
            O => \N__52266\,
            I => \N__51902\
        );

    \I__12336\ : ClkMux
    port map (
            O => \N__52265\,
            I => \N__51902\
        );

    \I__12335\ : ClkMux
    port map (
            O => \N__52264\,
            I => \N__51902\
        );

    \I__12334\ : ClkMux
    port map (
            O => \N__52263\,
            I => \N__51902\
        );

    \I__12333\ : ClkMux
    port map (
            O => \N__52262\,
            I => \N__51902\
        );

    \I__12332\ : ClkMux
    port map (
            O => \N__52261\,
            I => \N__51902\
        );

    \I__12331\ : ClkMux
    port map (
            O => \N__52260\,
            I => \N__51902\
        );

    \I__12330\ : ClkMux
    port map (
            O => \N__52259\,
            I => \N__51902\
        );

    \I__12329\ : ClkMux
    port map (
            O => \N__52258\,
            I => \N__51902\
        );

    \I__12328\ : ClkMux
    port map (
            O => \N__52257\,
            I => \N__51902\
        );

    \I__12327\ : ClkMux
    port map (
            O => \N__52256\,
            I => \N__51902\
        );

    \I__12326\ : ClkMux
    port map (
            O => \N__52255\,
            I => \N__51902\
        );

    \I__12325\ : ClkMux
    port map (
            O => \N__52254\,
            I => \N__51902\
        );

    \I__12324\ : ClkMux
    port map (
            O => \N__52253\,
            I => \N__51902\
        );

    \I__12323\ : ClkMux
    port map (
            O => \N__52252\,
            I => \N__51902\
        );

    \I__12322\ : ClkMux
    port map (
            O => \N__52251\,
            I => \N__51902\
        );

    \I__12321\ : ClkMux
    port map (
            O => \N__52250\,
            I => \N__51902\
        );

    \I__12320\ : ClkMux
    port map (
            O => \N__52249\,
            I => \N__51902\
        );

    \I__12319\ : ClkMux
    port map (
            O => \N__52248\,
            I => \N__51902\
        );

    \I__12318\ : ClkMux
    port map (
            O => \N__52247\,
            I => \N__51902\
        );

    \I__12317\ : ClkMux
    port map (
            O => \N__52246\,
            I => \N__51902\
        );

    \I__12316\ : ClkMux
    port map (
            O => \N__52245\,
            I => \N__51902\
        );

    \I__12315\ : ClkMux
    port map (
            O => \N__52244\,
            I => \N__51902\
        );

    \I__12314\ : ClkMux
    port map (
            O => \N__52243\,
            I => \N__51902\
        );

    \I__12313\ : ClkMux
    port map (
            O => \N__52242\,
            I => \N__51902\
        );

    \I__12312\ : ClkMux
    port map (
            O => \N__52241\,
            I => \N__51902\
        );

    \I__12311\ : ClkMux
    port map (
            O => \N__52240\,
            I => \N__51902\
        );

    \I__12310\ : ClkMux
    port map (
            O => \N__52239\,
            I => \N__51902\
        );

    \I__12309\ : ClkMux
    port map (
            O => \N__52238\,
            I => \N__51902\
        );

    \I__12308\ : ClkMux
    port map (
            O => \N__52237\,
            I => \N__51902\
        );

    \I__12307\ : ClkMux
    port map (
            O => \N__52236\,
            I => \N__51902\
        );

    \I__12306\ : ClkMux
    port map (
            O => \N__52235\,
            I => \N__51902\
        );

    \I__12305\ : ClkMux
    port map (
            O => \N__52234\,
            I => \N__51902\
        );

    \I__12304\ : ClkMux
    port map (
            O => \N__52233\,
            I => \N__51902\
        );

    \I__12303\ : ClkMux
    port map (
            O => \N__52232\,
            I => \N__51902\
        );

    \I__12302\ : ClkMux
    port map (
            O => \N__52231\,
            I => \N__51902\
        );

    \I__12301\ : ClkMux
    port map (
            O => \N__52230\,
            I => \N__51902\
        );

    \I__12300\ : ClkMux
    port map (
            O => \N__52229\,
            I => \N__51902\
        );

    \I__12299\ : ClkMux
    port map (
            O => \N__52228\,
            I => \N__51902\
        );

    \I__12298\ : ClkMux
    port map (
            O => \N__52227\,
            I => \N__51902\
        );

    \I__12297\ : ClkMux
    port map (
            O => \N__52226\,
            I => \N__51902\
        );

    \I__12296\ : ClkMux
    port map (
            O => \N__52225\,
            I => \N__51902\
        );

    \I__12295\ : ClkMux
    port map (
            O => \N__52224\,
            I => \N__51902\
        );

    \I__12294\ : ClkMux
    port map (
            O => \N__52223\,
            I => \N__51902\
        );

    \I__12293\ : ClkMux
    port map (
            O => \N__52222\,
            I => \N__51902\
        );

    \I__12292\ : ClkMux
    port map (
            O => \N__52221\,
            I => \N__51902\
        );

    \I__12291\ : ClkMux
    port map (
            O => \N__52220\,
            I => \N__51902\
        );

    \I__12290\ : ClkMux
    port map (
            O => \N__52219\,
            I => \N__51902\
        );

    \I__12289\ : ClkMux
    port map (
            O => \N__52218\,
            I => \N__51902\
        );

    \I__12288\ : ClkMux
    port map (
            O => \N__52217\,
            I => \N__51902\
        );

    \I__12287\ : ClkMux
    port map (
            O => \N__52216\,
            I => \N__51902\
        );

    \I__12286\ : ClkMux
    port map (
            O => \N__52215\,
            I => \N__51902\
        );

    \I__12285\ : ClkMux
    port map (
            O => \N__52214\,
            I => \N__51902\
        );

    \I__12284\ : ClkMux
    port map (
            O => \N__52213\,
            I => \N__51902\
        );

    \I__12283\ : ClkMux
    port map (
            O => \N__52212\,
            I => \N__51902\
        );

    \I__12282\ : ClkMux
    port map (
            O => \N__52211\,
            I => \N__51902\
        );

    \I__12281\ : ClkMux
    port map (
            O => \N__52210\,
            I => \N__51902\
        );

    \I__12280\ : ClkMux
    port map (
            O => \N__52209\,
            I => \N__51902\
        );

    \I__12279\ : ClkMux
    port map (
            O => \N__52208\,
            I => \N__51902\
        );

    \I__12278\ : ClkMux
    port map (
            O => \N__52207\,
            I => \N__51902\
        );

    \I__12277\ : ClkMux
    port map (
            O => \N__52206\,
            I => \N__51902\
        );

    \I__12276\ : ClkMux
    port map (
            O => \N__52205\,
            I => \N__51902\
        );

    \I__12275\ : ClkMux
    port map (
            O => \N__52204\,
            I => \N__51902\
        );

    \I__12274\ : ClkMux
    port map (
            O => \N__52203\,
            I => \N__51902\
        );

    \I__12273\ : ClkMux
    port map (
            O => \N__52202\,
            I => \N__51902\
        );

    \I__12272\ : ClkMux
    port map (
            O => \N__52201\,
            I => \N__51902\
        );

    \I__12271\ : GlobalMux
    port map (
            O => \N__51902\,
            I => \N__51899\
        );

    \I__12270\ : gio2CtrlBuf
    port map (
            O => \N__51899\,
            I => pll_clk128_g
        );

    \I__12269\ : CEMux
    port map (
            O => \N__51896\,
            I => \N__51891\
        );

    \I__12268\ : CEMux
    port map (
            O => \N__51895\,
            I => \N__51886\
        );

    \I__12267\ : CEMux
    port map (
            O => \N__51894\,
            I => \N__51883\
        );

    \I__12266\ : LocalMux
    port map (
            O => \N__51891\,
            I => \N__51879\
        );

    \I__12265\ : CEMux
    port map (
            O => \N__51890\,
            I => \N__51876\
        );

    \I__12264\ : CEMux
    port map (
            O => \N__51889\,
            I => \N__51873\
        );

    \I__12263\ : LocalMux
    port map (
            O => \N__51886\,
            I => \N__51869\
        );

    \I__12262\ : LocalMux
    port map (
            O => \N__51883\,
            I => \N__51866\
        );

    \I__12261\ : CEMux
    port map (
            O => \N__51882\,
            I => \N__51863\
        );

    \I__12260\ : Span4Mux_h
    port map (
            O => \N__51879\,
            I => \N__51858\
        );

    \I__12259\ : LocalMux
    port map (
            O => \N__51876\,
            I => \N__51858\
        );

    \I__12258\ : LocalMux
    port map (
            O => \N__51873\,
            I => \N__51855\
        );

    \I__12257\ : CEMux
    port map (
            O => \N__51872\,
            I => \N__51852\
        );

    \I__12256\ : Span4Mux_h
    port map (
            O => \N__51869\,
            I => \N__51849\
        );

    \I__12255\ : Span12Mux_s6_h
    port map (
            O => \N__51866\,
            I => \N__51844\
        );

    \I__12254\ : LocalMux
    port map (
            O => \N__51863\,
            I => \N__51844\
        );

    \I__12253\ : Span4Mux_h
    port map (
            O => \N__51858\,
            I => \N__51841\
        );

    \I__12252\ : Span4Mux_v
    port map (
            O => \N__51855\,
            I => \N__51836\
        );

    \I__12251\ : LocalMux
    port map (
            O => \N__51852\,
            I => \N__51836\
        );

    \I__12250\ : Odrv4
    port map (
            O => \N__51849\,
            I => \N_31_i\
        );

    \I__12249\ : Odrv12
    port map (
            O => \N__51844\,
            I => \N_31_i\
        );

    \I__12248\ : Odrv4
    port map (
            O => \N__51841\,
            I => \N_31_i\
        );

    \I__12247\ : Odrv4
    port map (
            O => \N__51836\,
            I => \N_31_i\
        );

    \I__12246\ : SRMux
    port map (
            O => \N__51827\,
            I => \N__51269\
        );

    \I__12245\ : SRMux
    port map (
            O => \N__51826\,
            I => \N__51269\
        );

    \I__12244\ : SRMux
    port map (
            O => \N__51825\,
            I => \N__51269\
        );

    \I__12243\ : SRMux
    port map (
            O => \N__51824\,
            I => \N__51269\
        );

    \I__12242\ : SRMux
    port map (
            O => \N__51823\,
            I => \N__51269\
        );

    \I__12241\ : SRMux
    port map (
            O => \N__51822\,
            I => \N__51269\
        );

    \I__12240\ : SRMux
    port map (
            O => \N__51821\,
            I => \N__51269\
        );

    \I__12239\ : SRMux
    port map (
            O => \N__51820\,
            I => \N__51269\
        );

    \I__12238\ : SRMux
    port map (
            O => \N__51819\,
            I => \N__51269\
        );

    \I__12237\ : SRMux
    port map (
            O => \N__51818\,
            I => \N__51269\
        );

    \I__12236\ : SRMux
    port map (
            O => \N__51817\,
            I => \N__51269\
        );

    \I__12235\ : SRMux
    port map (
            O => \N__51816\,
            I => \N__51269\
        );

    \I__12234\ : SRMux
    port map (
            O => \N__51815\,
            I => \N__51269\
        );

    \I__12233\ : SRMux
    port map (
            O => \N__51814\,
            I => \N__51269\
        );

    \I__12232\ : SRMux
    port map (
            O => \N__51813\,
            I => \N__51269\
        );

    \I__12231\ : SRMux
    port map (
            O => \N__51812\,
            I => \N__51269\
        );

    \I__12230\ : SRMux
    port map (
            O => \N__51811\,
            I => \N__51269\
        );

    \I__12229\ : SRMux
    port map (
            O => \N__51810\,
            I => \N__51269\
        );

    \I__12228\ : SRMux
    port map (
            O => \N__51809\,
            I => \N__51269\
        );

    \I__12227\ : SRMux
    port map (
            O => \N__51808\,
            I => \N__51269\
        );

    \I__12226\ : SRMux
    port map (
            O => \N__51807\,
            I => \N__51269\
        );

    \I__12225\ : SRMux
    port map (
            O => \N__51806\,
            I => \N__51269\
        );

    \I__12224\ : SRMux
    port map (
            O => \N__51805\,
            I => \N__51269\
        );

    \I__12223\ : SRMux
    port map (
            O => \N__51804\,
            I => \N__51269\
        );

    \I__12222\ : SRMux
    port map (
            O => \N__51803\,
            I => \N__51269\
        );

    \I__12221\ : SRMux
    port map (
            O => \N__51802\,
            I => \N__51269\
        );

    \I__12220\ : SRMux
    port map (
            O => \N__51801\,
            I => \N__51269\
        );

    \I__12219\ : SRMux
    port map (
            O => \N__51800\,
            I => \N__51269\
        );

    \I__12218\ : SRMux
    port map (
            O => \N__51799\,
            I => \N__51269\
        );

    \I__12217\ : SRMux
    port map (
            O => \N__51798\,
            I => \N__51269\
        );

    \I__12216\ : SRMux
    port map (
            O => \N__51797\,
            I => \N__51269\
        );

    \I__12215\ : SRMux
    port map (
            O => \N__51796\,
            I => \N__51269\
        );

    \I__12214\ : SRMux
    port map (
            O => \N__51795\,
            I => \N__51269\
        );

    \I__12213\ : SRMux
    port map (
            O => \N__51794\,
            I => \N__51269\
        );

    \I__12212\ : SRMux
    port map (
            O => \N__51793\,
            I => \N__51269\
        );

    \I__12211\ : SRMux
    port map (
            O => \N__51792\,
            I => \N__51269\
        );

    \I__12210\ : SRMux
    port map (
            O => \N__51791\,
            I => \N__51269\
        );

    \I__12209\ : SRMux
    port map (
            O => \N__51790\,
            I => \N__51269\
        );

    \I__12208\ : SRMux
    port map (
            O => \N__51789\,
            I => \N__51269\
        );

    \I__12207\ : SRMux
    port map (
            O => \N__51788\,
            I => \N__51269\
        );

    \I__12206\ : SRMux
    port map (
            O => \N__51787\,
            I => \N__51269\
        );

    \I__12205\ : SRMux
    port map (
            O => \N__51786\,
            I => \N__51269\
        );

    \I__12204\ : SRMux
    port map (
            O => \N__51785\,
            I => \N__51269\
        );

    \I__12203\ : SRMux
    port map (
            O => \N__51784\,
            I => \N__51269\
        );

    \I__12202\ : SRMux
    port map (
            O => \N__51783\,
            I => \N__51269\
        );

    \I__12201\ : SRMux
    port map (
            O => \N__51782\,
            I => \N__51269\
        );

    \I__12200\ : SRMux
    port map (
            O => \N__51781\,
            I => \N__51269\
        );

    \I__12199\ : SRMux
    port map (
            O => \N__51780\,
            I => \N__51269\
        );

    \I__12198\ : SRMux
    port map (
            O => \N__51779\,
            I => \N__51269\
        );

    \I__12197\ : SRMux
    port map (
            O => \N__51778\,
            I => \N__51269\
        );

    \I__12196\ : SRMux
    port map (
            O => \N__51777\,
            I => \N__51269\
        );

    \I__12195\ : SRMux
    port map (
            O => \N__51776\,
            I => \N__51269\
        );

    \I__12194\ : SRMux
    port map (
            O => \N__51775\,
            I => \N__51269\
        );

    \I__12193\ : SRMux
    port map (
            O => \N__51774\,
            I => \N__51269\
        );

    \I__12192\ : SRMux
    port map (
            O => \N__51773\,
            I => \N__51269\
        );

    \I__12191\ : SRMux
    port map (
            O => \N__51772\,
            I => \N__51269\
        );

    \I__12190\ : SRMux
    port map (
            O => \N__51771\,
            I => \N__51269\
        );

    \I__12189\ : SRMux
    port map (
            O => \N__51770\,
            I => \N__51269\
        );

    \I__12188\ : SRMux
    port map (
            O => \N__51769\,
            I => \N__51269\
        );

    \I__12187\ : SRMux
    port map (
            O => \N__51768\,
            I => \N__51269\
        );

    \I__12186\ : SRMux
    port map (
            O => \N__51767\,
            I => \N__51269\
        );

    \I__12185\ : SRMux
    port map (
            O => \N__51766\,
            I => \N__51269\
        );

    \I__12184\ : SRMux
    port map (
            O => \N__51765\,
            I => \N__51269\
        );

    \I__12183\ : SRMux
    port map (
            O => \N__51764\,
            I => \N__51269\
        );

    \I__12182\ : SRMux
    port map (
            O => \N__51763\,
            I => \N__51269\
        );

    \I__12181\ : SRMux
    port map (
            O => \N__51762\,
            I => \N__51269\
        );

    \I__12180\ : SRMux
    port map (
            O => \N__51761\,
            I => \N__51269\
        );

    \I__12179\ : SRMux
    port map (
            O => \N__51760\,
            I => \N__51269\
        );

    \I__12178\ : SRMux
    port map (
            O => \N__51759\,
            I => \N__51269\
        );

    \I__12177\ : SRMux
    port map (
            O => \N__51758\,
            I => \N__51269\
        );

    \I__12176\ : SRMux
    port map (
            O => \N__51757\,
            I => \N__51269\
        );

    \I__12175\ : SRMux
    port map (
            O => \N__51756\,
            I => \N__51269\
        );

    \I__12174\ : SRMux
    port map (
            O => \N__51755\,
            I => \N__51269\
        );

    \I__12173\ : SRMux
    port map (
            O => \N__51754\,
            I => \N__51269\
        );

    \I__12172\ : SRMux
    port map (
            O => \N__51753\,
            I => \N__51269\
        );

    \I__12171\ : SRMux
    port map (
            O => \N__51752\,
            I => \N__51269\
        );

    \I__12170\ : SRMux
    port map (
            O => \N__51751\,
            I => \N__51269\
        );

    \I__12169\ : SRMux
    port map (
            O => \N__51750\,
            I => \N__51269\
        );

    \I__12168\ : SRMux
    port map (
            O => \N__51749\,
            I => \N__51269\
        );

    \I__12167\ : SRMux
    port map (
            O => \N__51748\,
            I => \N__51269\
        );

    \I__12166\ : SRMux
    port map (
            O => \N__51747\,
            I => \N__51269\
        );

    \I__12165\ : SRMux
    port map (
            O => \N__51746\,
            I => \N__51269\
        );

    \I__12164\ : SRMux
    port map (
            O => \N__51745\,
            I => \N__51269\
        );

    \I__12163\ : SRMux
    port map (
            O => \N__51744\,
            I => \N__51269\
        );

    \I__12162\ : SRMux
    port map (
            O => \N__51743\,
            I => \N__51269\
        );

    \I__12161\ : SRMux
    port map (
            O => \N__51742\,
            I => \N__51269\
        );

    \I__12160\ : SRMux
    port map (
            O => \N__51741\,
            I => \N__51269\
        );

    \I__12159\ : SRMux
    port map (
            O => \N__51740\,
            I => \N__51269\
        );

    \I__12158\ : SRMux
    port map (
            O => \N__51739\,
            I => \N__51269\
        );

    \I__12157\ : SRMux
    port map (
            O => \N__51738\,
            I => \N__51269\
        );

    \I__12156\ : SRMux
    port map (
            O => \N__51737\,
            I => \N__51269\
        );

    \I__12155\ : SRMux
    port map (
            O => \N__51736\,
            I => \N__51269\
        );

    \I__12154\ : SRMux
    port map (
            O => \N__51735\,
            I => \N__51269\
        );

    \I__12153\ : SRMux
    port map (
            O => \N__51734\,
            I => \N__51269\
        );

    \I__12152\ : SRMux
    port map (
            O => \N__51733\,
            I => \N__51269\
        );

    \I__12151\ : SRMux
    port map (
            O => \N__51732\,
            I => \N__51269\
        );

    \I__12150\ : SRMux
    port map (
            O => \N__51731\,
            I => \N__51269\
        );

    \I__12149\ : SRMux
    port map (
            O => \N__51730\,
            I => \N__51269\
        );

    \I__12148\ : SRMux
    port map (
            O => \N__51729\,
            I => \N__51269\
        );

    \I__12147\ : SRMux
    port map (
            O => \N__51728\,
            I => \N__51269\
        );

    \I__12146\ : SRMux
    port map (
            O => \N__51727\,
            I => \N__51269\
        );

    \I__12145\ : SRMux
    port map (
            O => \N__51726\,
            I => \N__51269\
        );

    \I__12144\ : SRMux
    port map (
            O => \N__51725\,
            I => \N__51269\
        );

    \I__12143\ : SRMux
    port map (
            O => \N__51724\,
            I => \N__51269\
        );

    \I__12142\ : SRMux
    port map (
            O => \N__51723\,
            I => \N__51269\
        );

    \I__12141\ : SRMux
    port map (
            O => \N__51722\,
            I => \N__51269\
        );

    \I__12140\ : SRMux
    port map (
            O => \N__51721\,
            I => \N__51269\
        );

    \I__12139\ : SRMux
    port map (
            O => \N__51720\,
            I => \N__51269\
        );

    \I__12138\ : SRMux
    port map (
            O => \N__51719\,
            I => \N__51269\
        );

    \I__12137\ : SRMux
    port map (
            O => \N__51718\,
            I => \N__51269\
        );

    \I__12136\ : SRMux
    port map (
            O => \N__51717\,
            I => \N__51269\
        );

    \I__12135\ : SRMux
    port map (
            O => \N__51716\,
            I => \N__51269\
        );

    \I__12134\ : SRMux
    port map (
            O => \N__51715\,
            I => \N__51269\
        );

    \I__12133\ : SRMux
    port map (
            O => \N__51714\,
            I => \N__51269\
        );

    \I__12132\ : SRMux
    port map (
            O => \N__51713\,
            I => \N__51269\
        );

    \I__12131\ : SRMux
    port map (
            O => \N__51712\,
            I => \N__51269\
        );

    \I__12130\ : SRMux
    port map (
            O => \N__51711\,
            I => \N__51269\
        );

    \I__12129\ : SRMux
    port map (
            O => \N__51710\,
            I => \N__51269\
        );

    \I__12128\ : SRMux
    port map (
            O => \N__51709\,
            I => \N__51269\
        );

    \I__12127\ : SRMux
    port map (
            O => \N__51708\,
            I => \N__51269\
        );

    \I__12126\ : SRMux
    port map (
            O => \N__51707\,
            I => \N__51269\
        );

    \I__12125\ : SRMux
    port map (
            O => \N__51706\,
            I => \N__51269\
        );

    \I__12124\ : SRMux
    port map (
            O => \N__51705\,
            I => \N__51269\
        );

    \I__12123\ : SRMux
    port map (
            O => \N__51704\,
            I => \N__51269\
        );

    \I__12122\ : SRMux
    port map (
            O => \N__51703\,
            I => \N__51269\
        );

    \I__12121\ : SRMux
    port map (
            O => \N__51702\,
            I => \N__51269\
        );

    \I__12120\ : SRMux
    port map (
            O => \N__51701\,
            I => \N__51269\
        );

    \I__12119\ : SRMux
    port map (
            O => \N__51700\,
            I => \N__51269\
        );

    \I__12118\ : SRMux
    port map (
            O => \N__51699\,
            I => \N__51269\
        );

    \I__12117\ : SRMux
    port map (
            O => \N__51698\,
            I => \N__51269\
        );

    \I__12116\ : SRMux
    port map (
            O => \N__51697\,
            I => \N__51269\
        );

    \I__12115\ : SRMux
    port map (
            O => \N__51696\,
            I => \N__51269\
        );

    \I__12114\ : SRMux
    port map (
            O => \N__51695\,
            I => \N__51269\
        );

    \I__12113\ : SRMux
    port map (
            O => \N__51694\,
            I => \N__51269\
        );

    \I__12112\ : SRMux
    port map (
            O => \N__51693\,
            I => \N__51269\
        );

    \I__12111\ : SRMux
    port map (
            O => \N__51692\,
            I => \N__51269\
        );

    \I__12110\ : SRMux
    port map (
            O => \N__51691\,
            I => \N__51269\
        );

    \I__12109\ : SRMux
    port map (
            O => \N__51690\,
            I => \N__51269\
        );

    \I__12108\ : SRMux
    port map (
            O => \N__51689\,
            I => \N__51269\
        );

    \I__12107\ : SRMux
    port map (
            O => \N__51688\,
            I => \N__51269\
        );

    \I__12106\ : SRMux
    port map (
            O => \N__51687\,
            I => \N__51269\
        );

    \I__12105\ : SRMux
    port map (
            O => \N__51686\,
            I => \N__51269\
        );

    \I__12104\ : SRMux
    port map (
            O => \N__51685\,
            I => \N__51269\
        );

    \I__12103\ : SRMux
    port map (
            O => \N__51684\,
            I => \N__51269\
        );

    \I__12102\ : SRMux
    port map (
            O => \N__51683\,
            I => \N__51269\
        );

    \I__12101\ : SRMux
    port map (
            O => \N__51682\,
            I => \N__51269\
        );

    \I__12100\ : SRMux
    port map (
            O => \N__51681\,
            I => \N__51269\
        );

    \I__12099\ : SRMux
    port map (
            O => \N__51680\,
            I => \N__51269\
        );

    \I__12098\ : SRMux
    port map (
            O => \N__51679\,
            I => \N__51269\
        );

    \I__12097\ : SRMux
    port map (
            O => \N__51678\,
            I => \N__51269\
        );

    \I__12096\ : SRMux
    port map (
            O => \N__51677\,
            I => \N__51269\
        );

    \I__12095\ : SRMux
    port map (
            O => \N__51676\,
            I => \N__51269\
        );

    \I__12094\ : SRMux
    port map (
            O => \N__51675\,
            I => \N__51269\
        );

    \I__12093\ : SRMux
    port map (
            O => \N__51674\,
            I => \N__51269\
        );

    \I__12092\ : SRMux
    port map (
            O => \N__51673\,
            I => \N__51269\
        );

    \I__12091\ : SRMux
    port map (
            O => \N__51672\,
            I => \N__51269\
        );

    \I__12090\ : SRMux
    port map (
            O => \N__51671\,
            I => \N__51269\
        );

    \I__12089\ : SRMux
    port map (
            O => \N__51670\,
            I => \N__51269\
        );

    \I__12088\ : SRMux
    port map (
            O => \N__51669\,
            I => \N__51269\
        );

    \I__12087\ : SRMux
    port map (
            O => \N__51668\,
            I => \N__51269\
        );

    \I__12086\ : SRMux
    port map (
            O => \N__51667\,
            I => \N__51269\
        );

    \I__12085\ : SRMux
    port map (
            O => \N__51666\,
            I => \N__51269\
        );

    \I__12084\ : SRMux
    port map (
            O => \N__51665\,
            I => \N__51269\
        );

    \I__12083\ : SRMux
    port map (
            O => \N__51664\,
            I => \N__51269\
        );

    \I__12082\ : SRMux
    port map (
            O => \N__51663\,
            I => \N__51269\
        );

    \I__12081\ : SRMux
    port map (
            O => \N__51662\,
            I => \N__51269\
        );

    \I__12080\ : SRMux
    port map (
            O => \N__51661\,
            I => \N__51269\
        );

    \I__12079\ : SRMux
    port map (
            O => \N__51660\,
            I => \N__51269\
        );

    \I__12078\ : SRMux
    port map (
            O => \N__51659\,
            I => \N__51269\
        );

    \I__12077\ : SRMux
    port map (
            O => \N__51658\,
            I => \N__51269\
        );

    \I__12076\ : SRMux
    port map (
            O => \N__51657\,
            I => \N__51269\
        );

    \I__12075\ : SRMux
    port map (
            O => \N__51656\,
            I => \N__51269\
        );

    \I__12074\ : SRMux
    port map (
            O => \N__51655\,
            I => \N__51269\
        );

    \I__12073\ : SRMux
    port map (
            O => \N__51654\,
            I => \N__51269\
        );

    \I__12072\ : SRMux
    port map (
            O => \N__51653\,
            I => \N__51269\
        );

    \I__12071\ : SRMux
    port map (
            O => \N__51652\,
            I => \N__51269\
        );

    \I__12070\ : SRMux
    port map (
            O => \N__51651\,
            I => \N__51269\
        );

    \I__12069\ : SRMux
    port map (
            O => \N__51650\,
            I => \N__51269\
        );

    \I__12068\ : SRMux
    port map (
            O => \N__51649\,
            I => \N__51269\
        );

    \I__12067\ : SRMux
    port map (
            O => \N__51648\,
            I => \N__51269\
        );

    \I__12066\ : SRMux
    port map (
            O => \N__51647\,
            I => \N__51269\
        );

    \I__12065\ : SRMux
    port map (
            O => \N__51646\,
            I => \N__51269\
        );

    \I__12064\ : SRMux
    port map (
            O => \N__51645\,
            I => \N__51269\
        );

    \I__12063\ : SRMux
    port map (
            O => \N__51644\,
            I => \N__51269\
        );

    \I__12062\ : SRMux
    port map (
            O => \N__51643\,
            I => \N__51269\
        );

    \I__12061\ : SRMux
    port map (
            O => \N__51642\,
            I => \N__51269\
        );

    \I__12060\ : GlobalMux
    port map (
            O => \N__51269\,
            I => \N__51266\
        );

    \I__12059\ : gio2CtrlBuf
    port map (
            O => \N__51266\,
            I => \LED3_c_i_g\
        );

    \I__12058\ : InMux
    port map (
            O => \N__51263\,
            I => \N__51259\
        );

    \I__12057\ : InMux
    port map (
            O => \N__51262\,
            I => \N__51256\
        );

    \I__12056\ : LocalMux
    port map (
            O => \N__51259\,
            I => \N__51253\
        );

    \I__12055\ : LocalMux
    port map (
            O => \N__51256\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__12054\ : Odrv4
    port map (
            O => \N__51253\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__12053\ : InMux
    port map (
            O => \N__51248\,
            I => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3\
        );

    \I__12052\ : InMux
    port map (
            O => \N__51245\,
            I => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4\
        );

    \I__12051\ : InMux
    port map (
            O => \N__51242\,
            I => \N__51238\
        );

    \I__12050\ : InMux
    port map (
            O => \N__51241\,
            I => \N__51235\
        );

    \I__12049\ : LocalMux
    port map (
            O => \N__51238\,
            I => \N__51232\
        );

    \I__12048\ : LocalMux
    port map (
            O => \N__51235\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__12047\ : Odrv4
    port map (
            O => \N__51232\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__12046\ : InMux
    port map (
            O => \N__51227\,
            I => \N__51224\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__51224\,
            I => \N__51220\
        );

    \I__12044\ : InMux
    port map (
            O => \N__51223\,
            I => \N__51217\
        );

    \I__12043\ : Span4Mux_v
    port map (
            O => \N__51220\,
            I => \N__51208\
        );

    \I__12042\ : LocalMux
    port map (
            O => \N__51217\,
            I => \N__51208\
        );

    \I__12041\ : InMux
    port map (
            O => \N__51216\,
            I => \N__51205\
        );

    \I__12040\ : InMux
    port map (
            O => \N__51215\,
            I => \N__51198\
        );

    \I__12039\ : InMux
    port map (
            O => \N__51214\,
            I => \N__51198\
        );

    \I__12038\ : InMux
    port map (
            O => \N__51213\,
            I => \N__51198\
        );

    \I__12037\ : Span4Mux_v
    port map (
            O => \N__51208\,
            I => \N__51192\
        );

    \I__12036\ : LocalMux
    port map (
            O => \N__51205\,
            I => \N__51192\
        );

    \I__12035\ : LocalMux
    port map (
            O => \N__51198\,
            I => \N__51188\
        );

    \I__12034\ : InMux
    port map (
            O => \N__51197\,
            I => \N__51185\
        );

    \I__12033\ : Span4Mux_h
    port map (
            O => \N__51192\,
            I => \N__51182\
        );

    \I__12032\ : InMux
    port map (
            O => \N__51191\,
            I => \N__51179\
        );

    \I__12031\ : Span4Mux_v
    port map (
            O => \N__51188\,
            I => \N__51175\
        );

    \I__12030\ : LocalMux
    port map (
            O => \N__51185\,
            I => \N__51172\
        );

    \I__12029\ : Span4Mux_h
    port map (
            O => \N__51182\,
            I => \N__51169\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__51179\,
            I => \N__51166\
        );

    \I__12027\ : InMux
    port map (
            O => \N__51178\,
            I => \N__51163\
        );

    \I__12026\ : Span4Mux_v
    port map (
            O => \N__51175\,
            I => \N__51158\
        );

    \I__12025\ : Span4Mux_v
    port map (
            O => \N__51172\,
            I => \N__51158\
        );

    \I__12024\ : Span4Mux_h
    port map (
            O => \N__51169\,
            I => \N__51151\
        );

    \I__12023\ : Span4Mux_v
    port map (
            O => \N__51166\,
            I => \N__51151\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__51163\,
            I => \N__51151\
        );

    \I__12021\ : Odrv4
    port map (
            O => \N__51158\,
            I => \spi_slave_inst.spi_csZ0\
        );

    \I__12020\ : Odrv4
    port map (
            O => \N__51151\,
            I => \spi_slave_inst.spi_csZ0\
        );

    \I__12019\ : InMux
    port map (
            O => \N__51146\,
            I => \N__51138\
        );

    \I__12018\ : InMux
    port map (
            O => \N__51145\,
            I => \N__51138\
        );

    \I__12017\ : InMux
    port map (
            O => \N__51144\,
            I => \N__51133\
        );

    \I__12016\ : InMux
    port map (
            O => \N__51143\,
            I => \N__51133\
        );

    \I__12015\ : LocalMux
    port map (
            O => \N__51138\,
            I => \N__51128\
        );

    \I__12014\ : LocalMux
    port map (
            O => \N__51133\,
            I => \N__51128\
        );

    \I__12013\ : Odrv4
    port map (
            O => \N__51128\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_i6\
        );

    \I__12012\ : InMux
    port map (
            O => \N__51125\,
            I => \N__51121\
        );

    \I__12011\ : InMux
    port map (
            O => \N__51124\,
            I => \N__51118\
        );

    \I__12010\ : LocalMux
    port map (
            O => \N__51121\,
            I => \spi_slave_inst.tx_done_neg_sclk_iZ0\
        );

    \I__12009\ : LocalMux
    port map (
            O => \N__51118\,
            I => \spi_slave_inst.tx_done_neg_sclk_iZ0\
        );

    \I__12008\ : InMux
    port map (
            O => \N__51113\,
            I => \N__51110\
        );

    \I__12007\ : LocalMux
    port map (
            O => \N__51110\,
            I => \spi_slave_inst.tx_done_reg1_iZ0\
        );

    \I__12006\ : InMux
    port map (
            O => \N__51107\,
            I => \N__51104\
        );

    \I__12005\ : LocalMux
    port map (
            O => \N__51104\,
            I => \spi_slave_inst.tx_done_reg3_iZ0\
        );

    \I__12004\ : InMux
    port map (
            O => \N__51101\,
            I => \N__51097\
        );

    \I__12003\ : InMux
    port map (
            O => \N__51100\,
            I => \N__51094\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__51097\,
            I => \spi_slave_inst.tx_done_reg2_iZ0\
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__51094\,
            I => \spi_slave_inst.tx_done_reg2_iZ0\
        );

    \I__12000\ : InMux
    port map (
            O => \N__51089\,
            I => \N__51086\
        );

    \I__11999\ : LocalMux
    port map (
            O => \N__51086\,
            I => \N__51083\
        );

    \I__11998\ : Span4Mux_h
    port map (
            O => \N__51083\,
            I => \N__51080\
        );

    \I__11997\ : Odrv4
    port map (
            O => \N__51080\,
            I => \spi_slave_inst.un4_tx_done_reg2_i\
        );

    \I__11996\ : InMux
    port map (
            O => \N__51077\,
            I => \N__51071\
        );

    \I__11995\ : InMux
    port map (
            O => \N__51076\,
            I => \N__51065\
        );

    \I__11994\ : InMux
    port map (
            O => \N__51075\,
            I => \N__51059\
        );

    \I__11993\ : InMux
    port map (
            O => \N__51074\,
            I => \N__51056\
        );

    \I__11992\ : LocalMux
    port map (
            O => \N__51071\,
            I => \N__51047\
        );

    \I__11991\ : InMux
    port map (
            O => \N__51070\,
            I => \N__51044\
        );

    \I__11990\ : InMux
    port map (
            O => \N__51069\,
            I => \N__51034\
        );

    \I__11989\ : InMux
    port map (
            O => \N__51068\,
            I => \N__51031\
        );

    \I__11988\ : LocalMux
    port map (
            O => \N__51065\,
            I => \N__51026\
        );

    \I__11987\ : InMux
    port map (
            O => \N__51064\,
            I => \N__51023\
        );

    \I__11986\ : InMux
    port map (
            O => \N__51063\,
            I => \N__51020\
        );

    \I__11985\ : InMux
    port map (
            O => \N__51062\,
            I => \N__51014\
        );

    \I__11984\ : LocalMux
    port map (
            O => \N__51059\,
            I => \N__51009\
        );

    \I__11983\ : LocalMux
    port map (
            O => \N__51056\,
            I => \N__51009\
        );

    \I__11982\ : InMux
    port map (
            O => \N__51055\,
            I => \N__51006\
        );

    \I__11981\ : InMux
    port map (
            O => \N__51054\,
            I => \N__51003\
        );

    \I__11980\ : InMux
    port map (
            O => \N__51053\,
            I => \N__51000\
        );

    \I__11979\ : InMux
    port map (
            O => \N__51052\,
            I => \N__50997\
        );

    \I__11978\ : InMux
    port map (
            O => \N__51051\,
            I => \N__50994\
        );

    \I__11977\ : InMux
    port map (
            O => \N__51050\,
            I => \N__50991\
        );

    \I__11976\ : Span4Mux_h
    port map (
            O => \N__51047\,
            I => \N__50986\
        );

    \I__11975\ : LocalMux
    port map (
            O => \N__51044\,
            I => \N__50986\
        );

    \I__11974\ : InMux
    port map (
            O => \N__51043\,
            I => \N__50979\
        );

    \I__11973\ : InMux
    port map (
            O => \N__51042\,
            I => \N__50976\
        );

    \I__11972\ : InMux
    port map (
            O => \N__51041\,
            I => \N__50973\
        );

    \I__11971\ : InMux
    port map (
            O => \N__51040\,
            I => \N__50970\
        );

    \I__11970\ : InMux
    port map (
            O => \N__51039\,
            I => \N__50967\
        );

    \I__11969\ : InMux
    port map (
            O => \N__51038\,
            I => \N__50964\
        );

    \I__11968\ : InMux
    port map (
            O => \N__51037\,
            I => \N__50961\
        );

    \I__11967\ : LocalMux
    port map (
            O => \N__51034\,
            I => \N__50956\
        );

    \I__11966\ : LocalMux
    port map (
            O => \N__51031\,
            I => \N__50956\
        );

    \I__11965\ : InMux
    port map (
            O => \N__51030\,
            I => \N__50953\
        );

    \I__11964\ : InMux
    port map (
            O => \N__51029\,
            I => \N__50950\
        );

    \I__11963\ : Span4Mux_v
    port map (
            O => \N__51026\,
            I => \N__50943\
        );

    \I__11962\ : LocalMux
    port map (
            O => \N__51023\,
            I => \N__50943\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__51020\,
            I => \N__50943\
        );

    \I__11960\ : InMux
    port map (
            O => \N__51019\,
            I => \N__50940\
        );

    \I__11959\ : InMux
    port map (
            O => \N__51018\,
            I => \N__50935\
        );

    \I__11958\ : InMux
    port map (
            O => \N__51017\,
            I => \N__50932\
        );

    \I__11957\ : LocalMux
    port map (
            O => \N__51014\,
            I => \N__50925\
        );

    \I__11956\ : Span4Mux_h
    port map (
            O => \N__51009\,
            I => \N__50914\
        );

    \I__11955\ : LocalMux
    port map (
            O => \N__51006\,
            I => \N__50914\
        );

    \I__11954\ : LocalMux
    port map (
            O => \N__51003\,
            I => \N__50914\
        );

    \I__11953\ : LocalMux
    port map (
            O => \N__51000\,
            I => \N__50914\
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__50997\,
            I => \N__50914\
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__50994\,
            I => \N__50907\
        );

    \I__11950\ : LocalMux
    port map (
            O => \N__50991\,
            I => \N__50907\
        );

    \I__11949\ : Span4Mux_v
    port map (
            O => \N__50986\,
            I => \N__50907\
        );

    \I__11948\ : InMux
    port map (
            O => \N__50985\,
            I => \N__50904\
        );

    \I__11947\ : InMux
    port map (
            O => \N__50984\,
            I => \N__50900\
        );

    \I__11946\ : InMux
    port map (
            O => \N__50983\,
            I => \N__50893\
        );

    \I__11945\ : InMux
    port map (
            O => \N__50982\,
            I => \N__50889\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__50979\,
            I => \N__50884\
        );

    \I__11943\ : LocalMux
    port map (
            O => \N__50976\,
            I => \N__50884\
        );

    \I__11942\ : LocalMux
    port map (
            O => \N__50973\,
            I => \N__50872\
        );

    \I__11941\ : LocalMux
    port map (
            O => \N__50970\,
            I => \N__50872\
        );

    \I__11940\ : LocalMux
    port map (
            O => \N__50967\,
            I => \N__50861\
        );

    \I__11939\ : LocalMux
    port map (
            O => \N__50964\,
            I => \N__50861\
        );

    \I__11938\ : LocalMux
    port map (
            O => \N__50961\,
            I => \N__50861\
        );

    \I__11937\ : Span4Mux_h
    port map (
            O => \N__50956\,
            I => \N__50861\
        );

    \I__11936\ : LocalMux
    port map (
            O => \N__50953\,
            I => \N__50861\
        );

    \I__11935\ : LocalMux
    port map (
            O => \N__50950\,
            I => \N__50858\
        );

    \I__11934\ : Span4Mux_h
    port map (
            O => \N__50943\,
            I => \N__50855\
        );

    \I__11933\ : LocalMux
    port map (
            O => \N__50940\,
            I => \N__50852\
        );

    \I__11932\ : InMux
    port map (
            O => \N__50939\,
            I => \N__50848\
        );

    \I__11931\ : InMux
    port map (
            O => \N__50938\,
            I => \N__50845\
        );

    \I__11930\ : LocalMux
    port map (
            O => \N__50935\,
            I => \N__50840\
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__50932\,
            I => \N__50840\
        );

    \I__11928\ : InMux
    port map (
            O => \N__50931\,
            I => \N__50837\
        );

    \I__11927\ : InMux
    port map (
            O => \N__50930\,
            I => \N__50834\
        );

    \I__11926\ : InMux
    port map (
            O => \N__50929\,
            I => \N__50831\
        );

    \I__11925\ : InMux
    port map (
            O => \N__50928\,
            I => \N__50828\
        );

    \I__11924\ : Span4Mux_v
    port map (
            O => \N__50925\,
            I => \N__50825\
        );

    \I__11923\ : Span4Mux_v
    port map (
            O => \N__50914\,
            I => \N__50820\
        );

    \I__11922\ : Span4Mux_h
    port map (
            O => \N__50907\,
            I => \N__50820\
        );

    \I__11921\ : LocalMux
    port map (
            O => \N__50904\,
            I => \N__50817\
        );

    \I__11920\ : InMux
    port map (
            O => \N__50903\,
            I => \N__50811\
        );

    \I__11919\ : LocalMux
    port map (
            O => \N__50900\,
            I => \N__50808\
        );

    \I__11918\ : InMux
    port map (
            O => \N__50899\,
            I => \N__50805\
        );

    \I__11917\ : InMux
    port map (
            O => \N__50898\,
            I => \N__50802\
        );

    \I__11916\ : InMux
    port map (
            O => \N__50897\,
            I => \N__50799\
        );

    \I__11915\ : InMux
    port map (
            O => \N__50896\,
            I => \N__50796\
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__50893\,
            I => \N__50793\
        );

    \I__11913\ : InMux
    port map (
            O => \N__50892\,
            I => \N__50790\
        );

    \I__11912\ : LocalMux
    port map (
            O => \N__50889\,
            I => \N__50787\
        );

    \I__11911\ : Span4Mux_v
    port map (
            O => \N__50884\,
            I => \N__50784\
        );

    \I__11910\ : InMux
    port map (
            O => \N__50883\,
            I => \N__50781\
        );

    \I__11909\ : InMux
    port map (
            O => \N__50882\,
            I => \N__50778\
        );

    \I__11908\ : InMux
    port map (
            O => \N__50881\,
            I => \N__50775\
        );

    \I__11907\ : InMux
    port map (
            O => \N__50880\,
            I => \N__50772\
        );

    \I__11906\ : InMux
    port map (
            O => \N__50879\,
            I => \N__50769\
        );

    \I__11905\ : InMux
    port map (
            O => \N__50878\,
            I => \N__50766\
        );

    \I__11904\ : InMux
    port map (
            O => \N__50877\,
            I => \N__50763\
        );

    \I__11903\ : Span4Mux_v
    port map (
            O => \N__50872\,
            I => \N__50758\
        );

    \I__11902\ : Span4Mux_v
    port map (
            O => \N__50861\,
            I => \N__50758\
        );

    \I__11901\ : Span4Mux_v
    port map (
            O => \N__50858\,
            I => \N__50755\
        );

    \I__11900\ : Span4Mux_v
    port map (
            O => \N__50855\,
            I => \N__50750\
        );

    \I__11899\ : Span4Mux_v
    port map (
            O => \N__50852\,
            I => \N__50750\
        );

    \I__11898\ : InMux
    port map (
            O => \N__50851\,
            I => \N__50747\
        );

    \I__11897\ : LocalMux
    port map (
            O => \N__50848\,
            I => \N__50742\
        );

    \I__11896\ : LocalMux
    port map (
            O => \N__50845\,
            I => \N__50742\
        );

    \I__11895\ : Span4Mux_v
    port map (
            O => \N__50840\,
            I => \N__50739\
        );

    \I__11894\ : LocalMux
    port map (
            O => \N__50837\,
            I => \N__50724\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__50834\,
            I => \N__50724\
        );

    \I__11892\ : LocalMux
    port map (
            O => \N__50831\,
            I => \N__50724\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__50828\,
            I => \N__50724\
        );

    \I__11890\ : Span4Mux_v
    port map (
            O => \N__50825\,
            I => \N__50724\
        );

    \I__11889\ : Span4Mux_h
    port map (
            O => \N__50820\,
            I => \N__50724\
        );

    \I__11888\ : Span4Mux_h
    port map (
            O => \N__50817\,
            I => \N__50724\
        );

    \I__11887\ : InMux
    port map (
            O => \N__50816\,
            I => \N__50719\
        );

    \I__11886\ : InMux
    port map (
            O => \N__50815\,
            I => \N__50719\
        );

    \I__11885\ : InMux
    port map (
            O => \N__50814\,
            I => \N__50712\
        );

    \I__11884\ : LocalMux
    port map (
            O => \N__50811\,
            I => \N__50707\
        );

    \I__11883\ : Span4Mux_v
    port map (
            O => \N__50808\,
            I => \N__50707\
        );

    \I__11882\ : LocalMux
    port map (
            O => \N__50805\,
            I => \N__50696\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__50802\,
            I => \N__50696\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__50799\,
            I => \N__50696\
        );

    \I__11879\ : LocalMux
    port map (
            O => \N__50796\,
            I => \N__50696\
        );

    \I__11878\ : Span4Mux_v
    port map (
            O => \N__50793\,
            I => \N__50696\
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__50790\,
            I => \N__50689\
        );

    \I__11876\ : Span4Mux_v
    port map (
            O => \N__50787\,
            I => \N__50689\
        );

    \I__11875\ : Span4Mux_h
    port map (
            O => \N__50784\,
            I => \N__50689\
        );

    \I__11874\ : LocalMux
    port map (
            O => \N__50781\,
            I => \N__50682\
        );

    \I__11873\ : LocalMux
    port map (
            O => \N__50778\,
            I => \N__50682\
        );

    \I__11872\ : LocalMux
    port map (
            O => \N__50775\,
            I => \N__50682\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__50772\,
            I => \N__50667\
        );

    \I__11870\ : LocalMux
    port map (
            O => \N__50769\,
            I => \N__50667\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__50766\,
            I => \N__50667\
        );

    \I__11868\ : LocalMux
    port map (
            O => \N__50763\,
            I => \N__50667\
        );

    \I__11867\ : Sp12to4
    port map (
            O => \N__50758\,
            I => \N__50667\
        );

    \I__11866\ : Sp12to4
    port map (
            O => \N__50755\,
            I => \N__50667\
        );

    \I__11865\ : Sp12to4
    port map (
            O => \N__50750\,
            I => \N__50667\
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__50747\,
            I => \N__50664\
        );

    \I__11863\ : Span4Mux_v
    port map (
            O => \N__50742\,
            I => \N__50655\
        );

    \I__11862\ : Span4Mux_v
    port map (
            O => \N__50739\,
            I => \N__50655\
        );

    \I__11861\ : Span4Mux_v
    port map (
            O => \N__50724\,
            I => \N__50655\
        );

    \I__11860\ : LocalMux
    port map (
            O => \N__50719\,
            I => \N__50655\
        );

    \I__11859\ : InMux
    port map (
            O => \N__50718\,
            I => \N__50652\
        );

    \I__11858\ : InMux
    port map (
            O => \N__50717\,
            I => \N__50649\
        );

    \I__11857\ : InMux
    port map (
            O => \N__50716\,
            I => \N__50646\
        );

    \I__11856\ : InMux
    port map (
            O => \N__50715\,
            I => \N__50643\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__50712\,
            I => \N__50634\
        );

    \I__11854\ : Span4Mux_v
    port map (
            O => \N__50707\,
            I => \N__50634\
        );

    \I__11853\ : Span4Mux_v
    port map (
            O => \N__50696\,
            I => \N__50634\
        );

    \I__11852\ : Span4Mux_h
    port map (
            O => \N__50689\,
            I => \N__50634\
        );

    \I__11851\ : Span12Mux_v
    port map (
            O => \N__50682\,
            I => \N__50629\
        );

    \I__11850\ : Span12Mux_h
    port map (
            O => \N__50667\,
            I => \N__50629\
        );

    \I__11849\ : Span4Mux_v
    port map (
            O => \N__50664\,
            I => \N__50624\
        );

    \I__11848\ : Span4Mux_h
    port map (
            O => \N__50655\,
            I => \N__50624\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__50652\,
            I => spi_data_mosi_1
        );

    \I__11846\ : LocalMux
    port map (
            O => \N__50649\,
            I => spi_data_mosi_1
        );

    \I__11845\ : LocalMux
    port map (
            O => \N__50646\,
            I => spi_data_mosi_1
        );

    \I__11844\ : LocalMux
    port map (
            O => \N__50643\,
            I => spi_data_mosi_1
        );

    \I__11843\ : Odrv4
    port map (
            O => \N__50634\,
            I => spi_data_mosi_1
        );

    \I__11842\ : Odrv12
    port map (
            O => \N__50629\,
            I => spi_data_mosi_1
        );

    \I__11841\ : Odrv4
    port map (
            O => \N__50624\,
            I => spi_data_mosi_1
        );

    \I__11840\ : InMux
    port map (
            O => \N__50609\,
            I => \N__50606\
        );

    \I__11839\ : LocalMux
    port map (
            O => \N__50606\,
            I => \N__50603\
        );

    \I__11838\ : Span4Mux_h
    port map (
            O => \N__50603\,
            I => \N__50600\
        );

    \I__11837\ : Span4Mux_h
    port map (
            O => \N__50600\,
            I => \N__50597\
        );

    \I__11836\ : Odrv4
    port map (
            O => \N__50597\,
            I => \sDAC_mem_25Z0Z_1\
        );

    \I__11835\ : CEMux
    port map (
            O => \N__50594\,
            I => \N__50590\
        );

    \I__11834\ : CEMux
    port map (
            O => \N__50593\,
            I => \N__50587\
        );

    \I__11833\ : LocalMux
    port map (
            O => \N__50590\,
            I => \N__50584\
        );

    \I__11832\ : LocalMux
    port map (
            O => \N__50587\,
            I => \N__50581\
        );

    \I__11831\ : Span4Mux_v
    port map (
            O => \N__50584\,
            I => \N__50578\
        );

    \I__11830\ : Span4Mux_v
    port map (
            O => \N__50581\,
            I => \N__50575\
        );

    \I__11829\ : Odrv4
    port map (
            O => \N__50578\,
            I => \sDAC_mem_25_1_sqmuxa\
        );

    \I__11828\ : Odrv4
    port map (
            O => \N__50575\,
            I => \sDAC_mem_25_1_sqmuxa\
        );

    \I__11827\ : InMux
    port map (
            O => \N__50570\,
            I => \N__50567\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__50567\,
            I => \N__50564\
        );

    \I__11825\ : Span4Mux_h
    port map (
            O => \N__50564\,
            I => \N__50561\
        );

    \I__11824\ : Odrv4
    port map (
            O => \N__50561\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_7\
        );

    \I__11823\ : InMux
    port map (
            O => \N__50558\,
            I => \N__50555\
        );

    \I__11822\ : LocalMux
    port map (
            O => \N__50555\,
            I => \N__50552\
        );

    \I__11821\ : Span4Mux_v
    port map (
            O => \N__50552\,
            I => \N__50549\
        );

    \I__11820\ : Odrv4
    port map (
            O => \N__50549\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_7\
        );

    \I__11819\ : InMux
    port map (
            O => \N__50546\,
            I => \N__50538\
        );

    \I__11818\ : InMux
    port map (
            O => \N__50545\,
            I => \N__50535\
        );

    \I__11817\ : InMux
    port map (
            O => \N__50544\,
            I => \N__50532\
        );

    \I__11816\ : InMux
    port map (
            O => \N__50543\,
            I => \N__50523\
        );

    \I__11815\ : InMux
    port map (
            O => \N__50542\,
            I => \N__50520\
        );

    \I__11814\ : InMux
    port map (
            O => \N__50541\,
            I => \N__50517\
        );

    \I__11813\ : LocalMux
    port map (
            O => \N__50538\,
            I => \N__50513\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__50535\,
            I => \N__50508\
        );

    \I__11811\ : LocalMux
    port map (
            O => \N__50532\,
            I => \N__50508\
        );

    \I__11810\ : InMux
    port map (
            O => \N__50531\,
            I => \N__50505\
        );

    \I__11809\ : InMux
    port map (
            O => \N__50530\,
            I => \N__50502\
        );

    \I__11808\ : InMux
    port map (
            O => \N__50529\,
            I => \N__50499\
        );

    \I__11807\ : InMux
    port map (
            O => \N__50528\,
            I => \N__50496\
        );

    \I__11806\ : InMux
    port map (
            O => \N__50527\,
            I => \N__50492\
        );

    \I__11805\ : InMux
    port map (
            O => \N__50526\,
            I => \N__50489\
        );

    \I__11804\ : LocalMux
    port map (
            O => \N__50523\,
            I => \N__50473\
        );

    \I__11803\ : LocalMux
    port map (
            O => \N__50520\,
            I => \N__50473\
        );

    \I__11802\ : LocalMux
    port map (
            O => \N__50517\,
            I => \N__50473\
        );

    \I__11801\ : InMux
    port map (
            O => \N__50516\,
            I => \N__50470\
        );

    \I__11800\ : Span4Mux_h
    port map (
            O => \N__50513\,
            I => \N__50452\
        );

    \I__11799\ : Span4Mux_v
    port map (
            O => \N__50508\,
            I => \N__50452\
        );

    \I__11798\ : LocalMux
    port map (
            O => \N__50505\,
            I => \N__50452\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__50502\,
            I => \N__50452\
        );

    \I__11796\ : LocalMux
    port map (
            O => \N__50499\,
            I => \N__50452\
        );

    \I__11795\ : LocalMux
    port map (
            O => \N__50496\,
            I => \N__50449\
        );

    \I__11794\ : InMux
    port map (
            O => \N__50495\,
            I => \N__50446\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__50492\,
            I => \N__50443\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__50489\,
            I => \N__50440\
        );

    \I__11791\ : InMux
    port map (
            O => \N__50488\,
            I => \N__50437\
        );

    \I__11790\ : InMux
    port map (
            O => \N__50487\,
            I => \N__50434\
        );

    \I__11789\ : InMux
    port map (
            O => \N__50486\,
            I => \N__50431\
        );

    \I__11788\ : InMux
    port map (
            O => \N__50485\,
            I => \N__50427\
        );

    \I__11787\ : InMux
    port map (
            O => \N__50484\,
            I => \N__50424\
        );

    \I__11786\ : InMux
    port map (
            O => \N__50483\,
            I => \N__50421\
        );

    \I__11785\ : InMux
    port map (
            O => \N__50482\,
            I => \N__50417\
        );

    \I__11784\ : InMux
    port map (
            O => \N__50481\,
            I => \N__50414\
        );

    \I__11783\ : InMux
    port map (
            O => \N__50480\,
            I => \N__50410\
        );

    \I__11782\ : Span4Mux_v
    port map (
            O => \N__50473\,
            I => \N__50402\
        );

    \I__11781\ : LocalMux
    port map (
            O => \N__50470\,
            I => \N__50402\
        );

    \I__11780\ : InMux
    port map (
            O => \N__50469\,
            I => \N__50399\
        );

    \I__11779\ : InMux
    port map (
            O => \N__50468\,
            I => \N__50396\
        );

    \I__11778\ : InMux
    port map (
            O => \N__50467\,
            I => \N__50393\
        );

    \I__11777\ : InMux
    port map (
            O => \N__50466\,
            I => \N__50388\
        );

    \I__11776\ : InMux
    port map (
            O => \N__50465\,
            I => \N__50385\
        );

    \I__11775\ : InMux
    port map (
            O => \N__50464\,
            I => \N__50382\
        );

    \I__11774\ : InMux
    port map (
            O => \N__50463\,
            I => \N__50375\
        );

    \I__11773\ : Span4Mux_h
    port map (
            O => \N__50452\,
            I => \N__50367\
        );

    \I__11772\ : Span4Mux_v
    port map (
            O => \N__50449\,
            I => \N__50367\
        );

    \I__11771\ : LocalMux
    port map (
            O => \N__50446\,
            I => \N__50367\
        );

    \I__11770\ : Span4Mux_v
    port map (
            O => \N__50443\,
            I => \N__50356\
        );

    \I__11769\ : Span4Mux_h
    port map (
            O => \N__50440\,
            I => \N__50356\
        );

    \I__11768\ : LocalMux
    port map (
            O => \N__50437\,
            I => \N__50356\
        );

    \I__11767\ : LocalMux
    port map (
            O => \N__50434\,
            I => \N__50356\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__50431\,
            I => \N__50356\
        );

    \I__11765\ : InMux
    port map (
            O => \N__50430\,
            I => \N__50353\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__50427\,
            I => \N__50346\
        );

    \I__11763\ : LocalMux
    port map (
            O => \N__50424\,
            I => \N__50346\
        );

    \I__11762\ : LocalMux
    port map (
            O => \N__50421\,
            I => \N__50346\
        );

    \I__11761\ : InMux
    port map (
            O => \N__50420\,
            I => \N__50343\
        );

    \I__11760\ : LocalMux
    port map (
            O => \N__50417\,
            I => \N__50338\
        );

    \I__11759\ : LocalMux
    port map (
            O => \N__50414\,
            I => \N__50338\
        );

    \I__11758\ : InMux
    port map (
            O => \N__50413\,
            I => \N__50335\
        );

    \I__11757\ : LocalMux
    port map (
            O => \N__50410\,
            I => \N__50331\
        );

    \I__11756\ : InMux
    port map (
            O => \N__50409\,
            I => \N__50324\
        );

    \I__11755\ : InMux
    port map (
            O => \N__50408\,
            I => \N__50321\
        );

    \I__11754\ : InMux
    port map (
            O => \N__50407\,
            I => \N__50318\
        );

    \I__11753\ : Span4Mux_v
    port map (
            O => \N__50402\,
            I => \N__50310\
        );

    \I__11752\ : LocalMux
    port map (
            O => \N__50399\,
            I => \N__50310\
        );

    \I__11751\ : LocalMux
    port map (
            O => \N__50396\,
            I => \N__50310\
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__50393\,
            I => \N__50302\
        );

    \I__11749\ : InMux
    port map (
            O => \N__50392\,
            I => \N__50299\
        );

    \I__11748\ : InMux
    port map (
            O => \N__50391\,
            I => \N__50296\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__50388\,
            I => \N__50289\
        );

    \I__11746\ : LocalMux
    port map (
            O => \N__50385\,
            I => \N__50289\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__50382\,
            I => \N__50289\
        );

    \I__11744\ : InMux
    port map (
            O => \N__50381\,
            I => \N__50286\
        );

    \I__11743\ : InMux
    port map (
            O => \N__50380\,
            I => \N__50283\
        );

    \I__11742\ : InMux
    port map (
            O => \N__50379\,
            I => \N__50280\
        );

    \I__11741\ : InMux
    port map (
            O => \N__50378\,
            I => \N__50277\
        );

    \I__11740\ : LocalMux
    port map (
            O => \N__50375\,
            I => \N__50274\
        );

    \I__11739\ : InMux
    port map (
            O => \N__50374\,
            I => \N__50271\
        );

    \I__11738\ : Span4Mux_v
    port map (
            O => \N__50367\,
            I => \N__50268\
        );

    \I__11737\ : Span4Mux_v
    port map (
            O => \N__50356\,
            I => \N__50261\
        );

    \I__11736\ : LocalMux
    port map (
            O => \N__50353\,
            I => \N__50261\
        );

    \I__11735\ : Span4Mux_v
    port map (
            O => \N__50346\,
            I => \N__50261\
        );

    \I__11734\ : LocalMux
    port map (
            O => \N__50343\,
            I => \N__50254\
        );

    \I__11733\ : Span4Mux_v
    port map (
            O => \N__50338\,
            I => \N__50254\
        );

    \I__11732\ : LocalMux
    port map (
            O => \N__50335\,
            I => \N__50254\
        );

    \I__11731\ : InMux
    port map (
            O => \N__50334\,
            I => \N__50251\
        );

    \I__11730\ : Span12Mux_v
    port map (
            O => \N__50331\,
            I => \N__50248\
        );

    \I__11729\ : InMux
    port map (
            O => \N__50330\,
            I => \N__50245\
        );

    \I__11728\ : InMux
    port map (
            O => \N__50329\,
            I => \N__50242\
        );

    \I__11727\ : InMux
    port map (
            O => \N__50328\,
            I => \N__50239\
        );

    \I__11726\ : InMux
    port map (
            O => \N__50327\,
            I => \N__50236\
        );

    \I__11725\ : LocalMux
    port map (
            O => \N__50324\,
            I => \N__50229\
        );

    \I__11724\ : LocalMux
    port map (
            O => \N__50321\,
            I => \N__50229\
        );

    \I__11723\ : LocalMux
    port map (
            O => \N__50318\,
            I => \N__50229\
        );

    \I__11722\ : InMux
    port map (
            O => \N__50317\,
            I => \N__50226\
        );

    \I__11721\ : Span4Mux_v
    port map (
            O => \N__50310\,
            I => \N__50221\
        );

    \I__11720\ : InMux
    port map (
            O => \N__50309\,
            I => \N__50218\
        );

    \I__11719\ : InMux
    port map (
            O => \N__50308\,
            I => \N__50215\
        );

    \I__11718\ : InMux
    port map (
            O => \N__50307\,
            I => \N__50212\
        );

    \I__11717\ : InMux
    port map (
            O => \N__50306\,
            I => \N__50209\
        );

    \I__11716\ : InMux
    port map (
            O => \N__50305\,
            I => \N__50206\
        );

    \I__11715\ : Span12Mux_s9_v
    port map (
            O => \N__50302\,
            I => \N__50199\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__50299\,
            I => \N__50199\
        );

    \I__11713\ : LocalMux
    port map (
            O => \N__50296\,
            I => \N__50199\
        );

    \I__11712\ : Span4Mux_v
    port map (
            O => \N__50289\,
            I => \N__50196\
        );

    \I__11711\ : LocalMux
    port map (
            O => \N__50286\,
            I => \N__50189\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__50283\,
            I => \N__50189\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__50280\,
            I => \N__50189\
        );

    \I__11708\ : LocalMux
    port map (
            O => \N__50277\,
            I => \N__50186\
        );

    \I__11707\ : Span4Mux_v
    port map (
            O => \N__50274\,
            I => \N__50183\
        );

    \I__11706\ : LocalMux
    port map (
            O => \N__50271\,
            I => \N__50180\
        );

    \I__11705\ : Span4Mux_v
    port map (
            O => \N__50268\,
            I => \N__50171\
        );

    \I__11704\ : Span4Mux_h
    port map (
            O => \N__50261\,
            I => \N__50171\
        );

    \I__11703\ : Span4Mux_v
    port map (
            O => \N__50254\,
            I => \N__50171\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__50251\,
            I => \N__50171\
        );

    \I__11701\ : Span12Mux_h
    port map (
            O => \N__50248\,
            I => \N__50161\
        );

    \I__11700\ : LocalMux
    port map (
            O => \N__50245\,
            I => \N__50161\
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__50242\,
            I => \N__50161\
        );

    \I__11698\ : LocalMux
    port map (
            O => \N__50239\,
            I => \N__50156\
        );

    \I__11697\ : LocalMux
    port map (
            O => \N__50236\,
            I => \N__50156\
        );

    \I__11696\ : Span4Mux_v
    port map (
            O => \N__50229\,
            I => \N__50153\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__50226\,
            I => \N__50150\
        );

    \I__11694\ : InMux
    port map (
            O => \N__50225\,
            I => \N__50147\
        );

    \I__11693\ : InMux
    port map (
            O => \N__50224\,
            I => \N__50144\
        );

    \I__11692\ : Span4Mux_h
    port map (
            O => \N__50221\,
            I => \N__50131\
        );

    \I__11691\ : LocalMux
    port map (
            O => \N__50218\,
            I => \N__50131\
        );

    \I__11690\ : LocalMux
    port map (
            O => \N__50215\,
            I => \N__50131\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__50212\,
            I => \N__50131\
        );

    \I__11688\ : LocalMux
    port map (
            O => \N__50209\,
            I => \N__50131\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__50206\,
            I => \N__50131\
        );

    \I__11686\ : Span12Mux_v
    port map (
            O => \N__50199\,
            I => \N__50128\
        );

    \I__11685\ : Sp12to4
    port map (
            O => \N__50196\,
            I => \N__50117\
        );

    \I__11684\ : Span12Mux_v
    port map (
            O => \N__50189\,
            I => \N__50117\
        );

    \I__11683\ : Span12Mux_v
    port map (
            O => \N__50186\,
            I => \N__50117\
        );

    \I__11682\ : Sp12to4
    port map (
            O => \N__50183\,
            I => \N__50117\
        );

    \I__11681\ : Span12Mux_s10_h
    port map (
            O => \N__50180\,
            I => \N__50117\
        );

    \I__11680\ : Span4Mux_h
    port map (
            O => \N__50171\,
            I => \N__50114\
        );

    \I__11679\ : InMux
    port map (
            O => \N__50170\,
            I => \N__50111\
        );

    \I__11678\ : InMux
    port map (
            O => \N__50169\,
            I => \N__50108\
        );

    \I__11677\ : InMux
    port map (
            O => \N__50168\,
            I => \N__50105\
        );

    \I__11676\ : Span12Mux_v
    port map (
            O => \N__50161\,
            I => \N__50100\
        );

    \I__11675\ : Span12Mux_s11_h
    port map (
            O => \N__50156\,
            I => \N__50100\
        );

    \I__11674\ : Span4Mux_h
    port map (
            O => \N__50153\,
            I => \N__50089\
        );

    \I__11673\ : Span4Mux_v
    port map (
            O => \N__50150\,
            I => \N__50089\
        );

    \I__11672\ : LocalMux
    port map (
            O => \N__50147\,
            I => \N__50089\
        );

    \I__11671\ : LocalMux
    port map (
            O => \N__50144\,
            I => \N__50089\
        );

    \I__11670\ : Span4Mux_v
    port map (
            O => \N__50131\,
            I => \N__50089\
        );

    \I__11669\ : Odrv12
    port map (
            O => \N__50128\,
            I => spi_data_mosi_6
        );

    \I__11668\ : Odrv12
    port map (
            O => \N__50117\,
            I => spi_data_mosi_6
        );

    \I__11667\ : Odrv4
    port map (
            O => \N__50114\,
            I => spi_data_mosi_6
        );

    \I__11666\ : LocalMux
    port map (
            O => \N__50111\,
            I => spi_data_mosi_6
        );

    \I__11665\ : LocalMux
    port map (
            O => \N__50108\,
            I => spi_data_mosi_6
        );

    \I__11664\ : LocalMux
    port map (
            O => \N__50105\,
            I => spi_data_mosi_6
        );

    \I__11663\ : Odrv12
    port map (
            O => \N__50100\,
            I => spi_data_mosi_6
        );

    \I__11662\ : Odrv4
    port map (
            O => \N__50089\,
            I => spi_data_mosi_6
        );

    \I__11661\ : InMux
    port map (
            O => \N__50072\,
            I => \N__50069\
        );

    \I__11660\ : LocalMux
    port map (
            O => \N__50069\,
            I => \N__50066\
        );

    \I__11659\ : Odrv4
    port map (
            O => \N__50066\,
            I => \sEEADC_freqZ0Z_6\
        );

    \I__11658\ : InMux
    port map (
            O => \N__50063\,
            I => \N__50044\
        );

    \I__11657\ : InMux
    port map (
            O => \N__50062\,
            I => \N__50041\
        );

    \I__11656\ : InMux
    port map (
            O => \N__50061\,
            I => \N__50038\
        );

    \I__11655\ : InMux
    port map (
            O => \N__50060\,
            I => \N__50024\
        );

    \I__11654\ : InMux
    port map (
            O => \N__50059\,
            I => \N__50020\
        );

    \I__11653\ : InMux
    port map (
            O => \N__50058\,
            I => \N__50017\
        );

    \I__11652\ : InMux
    port map (
            O => \N__50057\,
            I => \N__50013\
        );

    \I__11651\ : InMux
    port map (
            O => \N__50056\,
            I => \N__50010\
        );

    \I__11650\ : InMux
    port map (
            O => \N__50055\,
            I => \N__50006\
        );

    \I__11649\ : InMux
    port map (
            O => \N__50054\,
            I => \N__50003\
        );

    \I__11648\ : InMux
    port map (
            O => \N__50053\,
            I => \N__50000\
        );

    \I__11647\ : InMux
    port map (
            O => \N__50052\,
            I => \N__49997\
        );

    \I__11646\ : InMux
    port map (
            O => \N__50051\,
            I => \N__49991\
        );

    \I__11645\ : InMux
    port map (
            O => \N__50050\,
            I => \N__49987\
        );

    \I__11644\ : InMux
    port map (
            O => \N__50049\,
            I => \N__49984\
        );

    \I__11643\ : InMux
    port map (
            O => \N__50048\,
            I => \N__49981\
        );

    \I__11642\ : InMux
    port map (
            O => \N__50047\,
            I => \N__49978\
        );

    \I__11641\ : LocalMux
    port map (
            O => \N__50044\,
            I => \N__49973\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__50041\,
            I => \N__49973\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__50038\,
            I => \N__49970\
        );

    \I__11638\ : InMux
    port map (
            O => \N__50037\,
            I => \N__49967\
        );

    \I__11637\ : InMux
    port map (
            O => \N__50036\,
            I => \N__49964\
        );

    \I__11636\ : InMux
    port map (
            O => \N__50035\,
            I => \N__49961\
        );

    \I__11635\ : InMux
    port map (
            O => \N__50034\,
            I => \N__49958\
        );

    \I__11634\ : InMux
    port map (
            O => \N__50033\,
            I => \N__49955\
        );

    \I__11633\ : InMux
    port map (
            O => \N__50032\,
            I => \N__49952\
        );

    \I__11632\ : InMux
    port map (
            O => \N__50031\,
            I => \N__49949\
        );

    \I__11631\ : InMux
    port map (
            O => \N__50030\,
            I => \N__49946\
        );

    \I__11630\ : InMux
    port map (
            O => \N__50029\,
            I => \N__49943\
        );

    \I__11629\ : InMux
    port map (
            O => \N__50028\,
            I => \N__49940\
        );

    \I__11628\ : InMux
    port map (
            O => \N__50027\,
            I => \N__49936\
        );

    \I__11627\ : LocalMux
    port map (
            O => \N__50024\,
            I => \N__49933\
        );

    \I__11626\ : InMux
    port map (
            O => \N__50023\,
            I => \N__49930\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__50020\,
            I => \N__49926\
        );

    \I__11624\ : LocalMux
    port map (
            O => \N__50017\,
            I => \N__49923\
        );

    \I__11623\ : InMux
    port map (
            O => \N__50016\,
            I => \N__49920\
        );

    \I__11622\ : LocalMux
    port map (
            O => \N__50013\,
            I => \N__49915\
        );

    \I__11621\ : LocalMux
    port map (
            O => \N__50010\,
            I => \N__49915\
        );

    \I__11620\ : InMux
    port map (
            O => \N__50009\,
            I => \N__49912\
        );

    \I__11619\ : LocalMux
    port map (
            O => \N__50006\,
            I => \N__49905\
        );

    \I__11618\ : LocalMux
    port map (
            O => \N__50003\,
            I => \N__49905\
        );

    \I__11617\ : LocalMux
    port map (
            O => \N__50000\,
            I => \N__49900\
        );

    \I__11616\ : LocalMux
    port map (
            O => \N__49997\,
            I => \N__49900\
        );

    \I__11615\ : InMux
    port map (
            O => \N__49996\,
            I => \N__49897\
        );

    \I__11614\ : InMux
    port map (
            O => \N__49995\,
            I => \N__49894\
        );

    \I__11613\ : CascadeMux
    port map (
            O => \N__49994\,
            I => \N__49889\
        );

    \I__11612\ : LocalMux
    port map (
            O => \N__49991\,
            I => \N__49886\
        );

    \I__11611\ : InMux
    port map (
            O => \N__49990\,
            I => \N__49883\
        );

    \I__11610\ : LocalMux
    port map (
            O => \N__49987\,
            I => \N__49880\
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__49984\,
            I => \N__49877\
        );

    \I__11608\ : LocalMux
    port map (
            O => \N__49981\,
            I => \N__49871\
        );

    \I__11607\ : LocalMux
    port map (
            O => \N__49978\,
            I => \N__49868\
        );

    \I__11606\ : Span4Mux_v
    port map (
            O => \N__49973\,
            I => \N__49848\
        );

    \I__11605\ : Span4Mux_h
    port map (
            O => \N__49970\,
            I => \N__49848\
        );

    \I__11604\ : LocalMux
    port map (
            O => \N__49967\,
            I => \N__49848\
        );

    \I__11603\ : LocalMux
    port map (
            O => \N__49964\,
            I => \N__49848\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__49961\,
            I => \N__49848\
        );

    \I__11601\ : LocalMux
    port map (
            O => \N__49958\,
            I => \N__49848\
        );

    \I__11600\ : LocalMux
    port map (
            O => \N__49955\,
            I => \N__49848\
        );

    \I__11599\ : LocalMux
    port map (
            O => \N__49952\,
            I => \N__49848\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__49949\,
            I => \N__49838\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__49946\,
            I => \N__49838\
        );

    \I__11596\ : LocalMux
    port map (
            O => \N__49943\,
            I => \N__49838\
        );

    \I__11595\ : LocalMux
    port map (
            O => \N__49940\,
            I => \N__49838\
        );

    \I__11594\ : InMux
    port map (
            O => \N__49939\,
            I => \N__49835\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__49936\,
            I => \N__49828\
        );

    \I__11592\ : Span4Mux_v
    port map (
            O => \N__49933\,
            I => \N__49823\
        );

    \I__11591\ : LocalMux
    port map (
            O => \N__49930\,
            I => \N__49823\
        );

    \I__11590\ : InMux
    port map (
            O => \N__49929\,
            I => \N__49820\
        );

    \I__11589\ : Span4Mux_h
    port map (
            O => \N__49926\,
            I => \N__49813\
        );

    \I__11588\ : Span4Mux_v
    port map (
            O => \N__49923\,
            I => \N__49813\
        );

    \I__11587\ : LocalMux
    port map (
            O => \N__49920\,
            I => \N__49813\
        );

    \I__11586\ : Span4Mux_v
    port map (
            O => \N__49915\,
            I => \N__49808\
        );

    \I__11585\ : LocalMux
    port map (
            O => \N__49912\,
            I => \N__49808\
        );

    \I__11584\ : InMux
    port map (
            O => \N__49911\,
            I => \N__49805\
        );

    \I__11583\ : InMux
    port map (
            O => \N__49910\,
            I => \N__49802\
        );

    \I__11582\ : Span4Mux_h
    port map (
            O => \N__49905\,
            I => \N__49793\
        );

    \I__11581\ : Span4Mux_v
    port map (
            O => \N__49900\,
            I => \N__49793\
        );

    \I__11580\ : LocalMux
    port map (
            O => \N__49897\,
            I => \N__49793\
        );

    \I__11579\ : LocalMux
    port map (
            O => \N__49894\,
            I => \N__49793\
        );

    \I__11578\ : InMux
    port map (
            O => \N__49893\,
            I => \N__49790\
        );

    \I__11577\ : InMux
    port map (
            O => \N__49892\,
            I => \N__49784\
        );

    \I__11576\ : InMux
    port map (
            O => \N__49889\,
            I => \N__49784\
        );

    \I__11575\ : Span4Mux_h
    port map (
            O => \N__49886\,
            I => \N__49779\
        );

    \I__11574\ : LocalMux
    port map (
            O => \N__49883\,
            I => \N__49779\
        );

    \I__11573\ : Span4Mux_h
    port map (
            O => \N__49880\,
            I => \N__49774\
        );

    \I__11572\ : Span4Mux_h
    port map (
            O => \N__49877\,
            I => \N__49774\
        );

    \I__11571\ : InMux
    port map (
            O => \N__49876\,
            I => \N__49771\
        );

    \I__11570\ : InMux
    port map (
            O => \N__49875\,
            I => \N__49768\
        );

    \I__11569\ : InMux
    port map (
            O => \N__49874\,
            I => \N__49765\
        );

    \I__11568\ : Span4Mux_h
    port map (
            O => \N__49871\,
            I => \N__49760\
        );

    \I__11567\ : Span4Mux_h
    port map (
            O => \N__49868\,
            I => \N__49760\
        );

    \I__11566\ : InMux
    port map (
            O => \N__49867\,
            I => \N__49757\
        );

    \I__11565\ : InMux
    port map (
            O => \N__49866\,
            I => \N__49754\
        );

    \I__11564\ : InMux
    port map (
            O => \N__49865\,
            I => \N__49751\
        );

    \I__11563\ : Span4Mux_v
    port map (
            O => \N__49848\,
            I => \N__49748\
        );

    \I__11562\ : InMux
    port map (
            O => \N__49847\,
            I => \N__49745\
        );

    \I__11561\ : Span4Mux_v
    port map (
            O => \N__49838\,
            I => \N__49740\
        );

    \I__11560\ : LocalMux
    port map (
            O => \N__49835\,
            I => \N__49740\
        );

    \I__11559\ : InMux
    port map (
            O => \N__49834\,
            I => \N__49737\
        );

    \I__11558\ : InMux
    port map (
            O => \N__49833\,
            I => \N__49734\
        );

    \I__11557\ : InMux
    port map (
            O => \N__49832\,
            I => \N__49731\
        );

    \I__11556\ : InMux
    port map (
            O => \N__49831\,
            I => \N__49728\
        );

    \I__11555\ : Span4Mux_h
    port map (
            O => \N__49828\,
            I => \N__49719\
        );

    \I__11554\ : Span4Mux_h
    port map (
            O => \N__49823\,
            I => \N__49719\
        );

    \I__11553\ : LocalMux
    port map (
            O => \N__49820\,
            I => \N__49719\
        );

    \I__11552\ : Span4Mux_v
    port map (
            O => \N__49813\,
            I => \N__49710\
        );

    \I__11551\ : Span4Mux_h
    port map (
            O => \N__49808\,
            I => \N__49710\
        );

    \I__11550\ : LocalMux
    port map (
            O => \N__49805\,
            I => \N__49710\
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__49802\,
            I => \N__49710\
        );

    \I__11548\ : Span4Mux_h
    port map (
            O => \N__49793\,
            I => \N__49705\
        );

    \I__11547\ : LocalMux
    port map (
            O => \N__49790\,
            I => \N__49705\
        );

    \I__11546\ : InMux
    port map (
            O => \N__49789\,
            I => \N__49702\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__49784\,
            I => \N__49699\
        );

    \I__11544\ : Sp12to4
    port map (
            O => \N__49779\,
            I => \N__49690\
        );

    \I__11543\ : Sp12to4
    port map (
            O => \N__49774\,
            I => \N__49690\
        );

    \I__11542\ : LocalMux
    port map (
            O => \N__49771\,
            I => \N__49690\
        );

    \I__11541\ : LocalMux
    port map (
            O => \N__49768\,
            I => \N__49690\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__49765\,
            I => \N__49681\
        );

    \I__11539\ : Sp12to4
    port map (
            O => \N__49760\,
            I => \N__49681\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__49757\,
            I => \N__49681\
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__49754\,
            I => \N__49681\
        );

    \I__11536\ : LocalMux
    port map (
            O => \N__49751\,
            I => \N__49678\
        );

    \I__11535\ : Sp12to4
    port map (
            O => \N__49748\,
            I => \N__49673\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__49745\,
            I => \N__49673\
        );

    \I__11533\ : Span4Mux_v
    port map (
            O => \N__49740\,
            I => \N__49662\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__49737\,
            I => \N__49662\
        );

    \I__11531\ : LocalMux
    port map (
            O => \N__49734\,
            I => \N__49662\
        );

    \I__11530\ : LocalMux
    port map (
            O => \N__49731\,
            I => \N__49662\
        );

    \I__11529\ : LocalMux
    port map (
            O => \N__49728\,
            I => \N__49659\
        );

    \I__11528\ : InMux
    port map (
            O => \N__49727\,
            I => \N__49656\
        );

    \I__11527\ : InMux
    port map (
            O => \N__49726\,
            I => \N__49651\
        );

    \I__11526\ : Span4Mux_v
    port map (
            O => \N__49719\,
            I => \N__49648\
        );

    \I__11525\ : Span4Mux_v
    port map (
            O => \N__49710\,
            I => \N__49639\
        );

    \I__11524\ : Span4Mux_v
    port map (
            O => \N__49705\,
            I => \N__49639\
        );

    \I__11523\ : LocalMux
    port map (
            O => \N__49702\,
            I => \N__49639\
        );

    \I__11522\ : Span4Mux_h
    port map (
            O => \N__49699\,
            I => \N__49639\
        );

    \I__11521\ : Span12Mux_v
    port map (
            O => \N__49690\,
            I => \N__49636\
        );

    \I__11520\ : Span12Mux_v
    port map (
            O => \N__49681\,
            I => \N__49629\
        );

    \I__11519\ : Span12Mux_s10_v
    port map (
            O => \N__49678\,
            I => \N__49629\
        );

    \I__11518\ : Span12Mux_s11_h
    port map (
            O => \N__49673\,
            I => \N__49629\
        );

    \I__11517\ : InMux
    port map (
            O => \N__49672\,
            I => \N__49626\
        );

    \I__11516\ : InMux
    port map (
            O => \N__49671\,
            I => \N__49623\
        );

    \I__11515\ : Span4Mux_v
    port map (
            O => \N__49662\,
            I => \N__49616\
        );

    \I__11514\ : Span4Mux_v
    port map (
            O => \N__49659\,
            I => \N__49616\
        );

    \I__11513\ : LocalMux
    port map (
            O => \N__49656\,
            I => \N__49616\
        );

    \I__11512\ : InMux
    port map (
            O => \N__49655\,
            I => \N__49613\
        );

    \I__11511\ : InMux
    port map (
            O => \N__49654\,
            I => \N__49610\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__49651\,
            I => \N__49603\
        );

    \I__11509\ : Span4Mux_h
    port map (
            O => \N__49648\,
            I => \N__49603\
        );

    \I__11508\ : Span4Mux_h
    port map (
            O => \N__49639\,
            I => \N__49603\
        );

    \I__11507\ : Odrv12
    port map (
            O => \N__49636\,
            I => spi_data_mosi_7
        );

    \I__11506\ : Odrv12
    port map (
            O => \N__49629\,
            I => spi_data_mosi_7
        );

    \I__11505\ : LocalMux
    port map (
            O => \N__49626\,
            I => spi_data_mosi_7
        );

    \I__11504\ : LocalMux
    port map (
            O => \N__49623\,
            I => spi_data_mosi_7
        );

    \I__11503\ : Odrv4
    port map (
            O => \N__49616\,
            I => spi_data_mosi_7
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__49613\,
            I => spi_data_mosi_7
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__49610\,
            I => spi_data_mosi_7
        );

    \I__11500\ : Odrv4
    port map (
            O => \N__49603\,
            I => spi_data_mosi_7
        );

    \I__11499\ : InMux
    port map (
            O => \N__49586\,
            I => \N__49583\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__49583\,
            I => \sEEADC_freqZ0Z_7\
        );

    \I__11497\ : CEMux
    port map (
            O => \N__49580\,
            I => \N__49577\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__49577\,
            I => \N__49573\
        );

    \I__11495\ : CEMux
    port map (
            O => \N__49576\,
            I => \N__49570\
        );

    \I__11494\ : Span4Mux_h
    port map (
            O => \N__49573\,
            I => \N__49565\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__49570\,
            I => \N__49565\
        );

    \I__11492\ : Span4Mux_h
    port map (
            O => \N__49565\,
            I => \N__49562\
        );

    \I__11491\ : Span4Mux_h
    port map (
            O => \N__49562\,
            I => \N__49558\
        );

    \I__11490\ : CEMux
    port map (
            O => \N__49561\,
            I => \N__49555\
        );

    \I__11489\ : Span4Mux_h
    port map (
            O => \N__49558\,
            I => \N__49550\
        );

    \I__11488\ : LocalMux
    port map (
            O => \N__49555\,
            I => \N__49550\
        );

    \I__11487\ : Span4Mux_v
    port map (
            O => \N__49550\,
            I => \N__49547\
        );

    \I__11486\ : Span4Mux_v
    port map (
            O => \N__49547\,
            I => \N__49544\
        );

    \I__11485\ : Span4Mux_v
    port map (
            O => \N__49544\,
            I => \N__49541\
        );

    \I__11484\ : Odrv4
    port map (
            O => \N__49541\,
            I => \sEEADC_freq_1_sqmuxa\
        );

    \I__11483\ : InMux
    port map (
            O => \N__49538\,
            I => \N__49519\
        );

    \I__11482\ : InMux
    port map (
            O => \N__49537\,
            I => \N__49519\
        );

    \I__11481\ : InMux
    port map (
            O => \N__49536\,
            I => \N__49519\
        );

    \I__11480\ : InMux
    port map (
            O => \N__49535\,
            I => \N__49510\
        );

    \I__11479\ : InMux
    port map (
            O => \N__49534\,
            I => \N__49510\
        );

    \I__11478\ : InMux
    port map (
            O => \N__49533\,
            I => \N__49510\
        );

    \I__11477\ : InMux
    port map (
            O => \N__49532\,
            I => \N__49510\
        );

    \I__11476\ : InMux
    port map (
            O => \N__49531\,
            I => \N__49505\
        );

    \I__11475\ : InMux
    port map (
            O => \N__49530\,
            I => \N__49505\
        );

    \I__11474\ : InMux
    port map (
            O => \N__49529\,
            I => \N__49496\
        );

    \I__11473\ : InMux
    port map (
            O => \N__49528\,
            I => \N__49496\
        );

    \I__11472\ : InMux
    port map (
            O => \N__49527\,
            I => \N__49496\
        );

    \I__11471\ : InMux
    port map (
            O => \N__49526\,
            I => \N__49496\
        );

    \I__11470\ : LocalMux
    port map (
            O => \N__49519\,
            I => \N__49485\
        );

    \I__11469\ : LocalMux
    port map (
            O => \N__49510\,
            I => \N__49485\
        );

    \I__11468\ : LocalMux
    port map (
            O => \N__49505\,
            I => \N__49485\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__49496\,
            I => \N__49485\
        );

    \I__11466\ : CascadeMux
    port map (
            O => \N__49495\,
            I => \N__49480\
        );

    \I__11465\ : InMux
    port map (
            O => \N__49494\,
            I => \N__49476\
        );

    \I__11464\ : Span4Mux_v
    port map (
            O => \N__49485\,
            I => \N__49473\
        );

    \I__11463\ : InMux
    port map (
            O => \N__49484\,
            I => \N__49470\
        );

    \I__11462\ : InMux
    port map (
            O => \N__49483\,
            I => \N__49463\
        );

    \I__11461\ : InMux
    port map (
            O => \N__49480\,
            I => \N__49463\
        );

    \I__11460\ : InMux
    port map (
            O => \N__49479\,
            I => \N__49463\
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__49476\,
            I => \N__49453\
        );

    \I__11458\ : Sp12to4
    port map (
            O => \N__49473\,
            I => \N__49453\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__49470\,
            I => \N__49453\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__49463\,
            I => \N__49453\
        );

    \I__11455\ : InMux
    port map (
            O => \N__49462\,
            I => \N__49450\
        );

    \I__11454\ : Odrv12
    port map (
            O => \N__49453\,
            I => \N_71\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__49450\,
            I => \N_71\
        );

    \I__11452\ : InMux
    port map (
            O => \N__49445\,
            I => \N__49442\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__49442\,
            I => \N__49423\
        );

    \I__11450\ : CEMux
    port map (
            O => \N__49441\,
            I => \N__49420\
        );

    \I__11449\ : CascadeMux
    port map (
            O => \N__49440\,
            I => \N__49414\
        );

    \I__11448\ : CascadeMux
    port map (
            O => \N__49439\,
            I => \N__49410\
        );

    \I__11447\ : CascadeMux
    port map (
            O => \N__49438\,
            I => \N__49407\
        );

    \I__11446\ : CascadeMux
    port map (
            O => \N__49437\,
            I => \N__49401\
        );

    \I__11445\ : CascadeMux
    port map (
            O => \N__49436\,
            I => \N__49397\
        );

    \I__11444\ : CascadeMux
    port map (
            O => \N__49435\,
            I => \N__49394\
        );

    \I__11443\ : CascadeMux
    port map (
            O => \N__49434\,
            I => \N__49391\
        );

    \I__11442\ : CascadeMux
    port map (
            O => \N__49433\,
            I => \N__49387\
        );

    \I__11441\ : CascadeMux
    port map (
            O => \N__49432\,
            I => \N__49383\
        );

    \I__11440\ : InMux
    port map (
            O => \N__49431\,
            I => \N__49372\
        );

    \I__11439\ : InMux
    port map (
            O => \N__49430\,
            I => \N__49372\
        );

    \I__11438\ : InMux
    port map (
            O => \N__49429\,
            I => \N__49372\
        );

    \I__11437\ : InMux
    port map (
            O => \N__49428\,
            I => \N__49372\
        );

    \I__11436\ : InMux
    port map (
            O => \N__49427\,
            I => \N__49369\
        );

    \I__11435\ : CEMux
    port map (
            O => \N__49426\,
            I => \N__49366\
        );

    \I__11434\ : Span4Mux_v
    port map (
            O => \N__49423\,
            I => \N__49359\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__49420\,
            I => \N__49356\
        );

    \I__11432\ : IoInMux
    port map (
            O => \N__49419\,
            I => \N__49349\
        );

    \I__11431\ : InMux
    port map (
            O => \N__49418\,
            I => \N__49338\
        );

    \I__11430\ : InMux
    port map (
            O => \N__49417\,
            I => \N__49338\
        );

    \I__11429\ : InMux
    port map (
            O => \N__49414\,
            I => \N__49338\
        );

    \I__11428\ : InMux
    port map (
            O => \N__49413\,
            I => \N__49338\
        );

    \I__11427\ : InMux
    port map (
            O => \N__49410\,
            I => \N__49338\
        );

    \I__11426\ : InMux
    port map (
            O => \N__49407\,
            I => \N__49321\
        );

    \I__11425\ : InMux
    port map (
            O => \N__49406\,
            I => \N__49321\
        );

    \I__11424\ : InMux
    port map (
            O => \N__49405\,
            I => \N__49321\
        );

    \I__11423\ : InMux
    port map (
            O => \N__49404\,
            I => \N__49321\
        );

    \I__11422\ : InMux
    port map (
            O => \N__49401\,
            I => \N__49321\
        );

    \I__11421\ : InMux
    port map (
            O => \N__49400\,
            I => \N__49321\
        );

    \I__11420\ : InMux
    port map (
            O => \N__49397\,
            I => \N__49321\
        );

    \I__11419\ : InMux
    port map (
            O => \N__49394\,
            I => \N__49321\
        );

    \I__11418\ : InMux
    port map (
            O => \N__49391\,
            I => \N__49318\
        );

    \I__11417\ : CascadeMux
    port map (
            O => \N__49390\,
            I => \N__49315\
        );

    \I__11416\ : InMux
    port map (
            O => \N__49387\,
            I => \N__49308\
        );

    \I__11415\ : InMux
    port map (
            O => \N__49386\,
            I => \N__49308\
        );

    \I__11414\ : InMux
    port map (
            O => \N__49383\,
            I => \N__49308\
        );

    \I__11413\ : InMux
    port map (
            O => \N__49382\,
            I => \N__49299\
        );

    \I__11412\ : InMux
    port map (
            O => \N__49381\,
            I => \N__49296\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__49372\,
            I => \N__49283\
        );

    \I__11410\ : LocalMux
    port map (
            O => \N__49369\,
            I => \N__49283\
        );

    \I__11409\ : LocalMux
    port map (
            O => \N__49366\,
            I => \N__49280\
        );

    \I__11408\ : InMux
    port map (
            O => \N__49365\,
            I => \N__49275\
        );

    \I__11407\ : InMux
    port map (
            O => \N__49364\,
            I => \N__49275\
        );

    \I__11406\ : CascadeMux
    port map (
            O => \N__49363\,
            I => \N__49272\
        );

    \I__11405\ : CascadeMux
    port map (
            O => \N__49362\,
            I => \N__49269\
        );

    \I__11404\ : Span4Mux_h
    port map (
            O => \N__49359\,
            I => \N__49264\
        );

    \I__11403\ : Span4Mux_v
    port map (
            O => \N__49356\,
            I => \N__49264\
        );

    \I__11402\ : CascadeMux
    port map (
            O => \N__49355\,
            I => \N__49261\
        );

    \I__11401\ : InMux
    port map (
            O => \N__49354\,
            I => \N__49257\
        );

    \I__11400\ : CascadeMux
    port map (
            O => \N__49353\,
            I => \N__49254\
        );

    \I__11399\ : CascadeMux
    port map (
            O => \N__49352\,
            I => \N__49250\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__49349\,
            I => \N__49247\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__49338\,
            I => \N__49241\
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__49321\,
            I => \N__49241\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__49318\,
            I => \N__49237\
        );

    \I__11394\ : InMux
    port map (
            O => \N__49315\,
            I => \N__49234\
        );

    \I__11393\ : LocalMux
    port map (
            O => \N__49308\,
            I => \N__49231\
        );

    \I__11392\ : InMux
    port map (
            O => \N__49307\,
            I => \N__49224\
        );

    \I__11391\ : InMux
    port map (
            O => \N__49306\,
            I => \N__49224\
        );

    \I__11390\ : InMux
    port map (
            O => \N__49305\,
            I => \N__49224\
        );

    \I__11389\ : InMux
    port map (
            O => \N__49304\,
            I => \N__49217\
        );

    \I__11388\ : InMux
    port map (
            O => \N__49303\,
            I => \N__49217\
        );

    \I__11387\ : InMux
    port map (
            O => \N__49302\,
            I => \N__49217\
        );

    \I__11386\ : LocalMux
    port map (
            O => \N__49299\,
            I => \N__49212\
        );

    \I__11385\ : LocalMux
    port map (
            O => \N__49296\,
            I => \N__49212\
        );

    \I__11384\ : InMux
    port map (
            O => \N__49295\,
            I => \N__49203\
        );

    \I__11383\ : InMux
    port map (
            O => \N__49294\,
            I => \N__49203\
        );

    \I__11382\ : InMux
    port map (
            O => \N__49293\,
            I => \N__49203\
        );

    \I__11381\ : InMux
    port map (
            O => \N__49292\,
            I => \N__49203\
        );

    \I__11380\ : InMux
    port map (
            O => \N__49291\,
            I => \N__49194\
        );

    \I__11379\ : InMux
    port map (
            O => \N__49290\,
            I => \N__49194\
        );

    \I__11378\ : InMux
    port map (
            O => \N__49289\,
            I => \N__49194\
        );

    \I__11377\ : InMux
    port map (
            O => \N__49288\,
            I => \N__49194\
        );

    \I__11376\ : Span4Mux_v
    port map (
            O => \N__49283\,
            I => \N__49188\
        );

    \I__11375\ : Span4Mux_h
    port map (
            O => \N__49280\,
            I => \N__49185\
        );

    \I__11374\ : LocalMux
    port map (
            O => \N__49275\,
            I => \N__49182\
        );

    \I__11373\ : InMux
    port map (
            O => \N__49272\,
            I => \N__49179\
        );

    \I__11372\ : InMux
    port map (
            O => \N__49269\,
            I => \N__49176\
        );

    \I__11371\ : Span4Mux_v
    port map (
            O => \N__49264\,
            I => \N__49173\
        );

    \I__11370\ : InMux
    port map (
            O => \N__49261\,
            I => \N__49170\
        );

    \I__11369\ : CascadeMux
    port map (
            O => \N__49260\,
            I => \N__49167\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__49257\,
            I => \N__49164\
        );

    \I__11367\ : InMux
    port map (
            O => \N__49254\,
            I => \N__49161\
        );

    \I__11366\ : InMux
    port map (
            O => \N__49253\,
            I => \N__49158\
        );

    \I__11365\ : InMux
    port map (
            O => \N__49250\,
            I => \N__49155\
        );

    \I__11364\ : Span4Mux_s2_h
    port map (
            O => \N__49247\,
            I => \N__49152\
        );

    \I__11363\ : InMux
    port map (
            O => \N__49246\,
            I => \N__49149\
        );

    \I__11362\ : Span4Mux_v
    port map (
            O => \N__49241\,
            I => \N__49146\
        );

    \I__11361\ : InMux
    port map (
            O => \N__49240\,
            I => \N__49142\
        );

    \I__11360\ : Span4Mux_v
    port map (
            O => \N__49237\,
            I => \N__49137\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__49234\,
            I => \N__49137\
        );

    \I__11358\ : Span4Mux_h
    port map (
            O => \N__49231\,
            I => \N__49124\
        );

    \I__11357\ : LocalMux
    port map (
            O => \N__49224\,
            I => \N__49124\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__49217\,
            I => \N__49124\
        );

    \I__11355\ : Span4Mux_h
    port map (
            O => \N__49212\,
            I => \N__49124\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__49203\,
            I => \N__49124\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__49194\,
            I => \N__49124\
        );

    \I__11352\ : InMux
    port map (
            O => \N__49193\,
            I => \N__49117\
        );

    \I__11351\ : InMux
    port map (
            O => \N__49192\,
            I => \N__49117\
        );

    \I__11350\ : InMux
    port map (
            O => \N__49191\,
            I => \N__49117\
        );

    \I__11349\ : Span4Mux_h
    port map (
            O => \N__49188\,
            I => \N__49105\
        );

    \I__11348\ : Span4Mux_h
    port map (
            O => \N__49185\,
            I => \N__49105\
        );

    \I__11347\ : Span4Mux_h
    port map (
            O => \N__49182\,
            I => \N__49105\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__49179\,
            I => \N__49105\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__49176\,
            I => \N__49105\
        );

    \I__11344\ : Span4Mux_h
    port map (
            O => \N__49173\,
            I => \N__49102\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__49170\,
            I => \N__49099\
        );

    \I__11342\ : InMux
    port map (
            O => \N__49167\,
            I => \N__49096\
        );

    \I__11341\ : Span4Mux_v
    port map (
            O => \N__49164\,
            I => \N__49088\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__49161\,
            I => \N__49088\
        );

    \I__11339\ : LocalMux
    port map (
            O => \N__49158\,
            I => \N__49088\
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__49155\,
            I => \N__49085\
        );

    \I__11337\ : Sp12to4
    port map (
            O => \N__49152\,
            I => \N__49082\
        );

    \I__11336\ : LocalMux
    port map (
            O => \N__49149\,
            I => \N__49079\
        );

    \I__11335\ : Span4Mux_v
    port map (
            O => \N__49146\,
            I => \N__49076\
        );

    \I__11334\ : InMux
    port map (
            O => \N__49145\,
            I => \N__49073\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__49142\,
            I => \N__49064\
        );

    \I__11332\ : Span4Mux_v
    port map (
            O => \N__49137\,
            I => \N__49064\
        );

    \I__11331\ : Span4Mux_v
    port map (
            O => \N__49124\,
            I => \N__49064\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__49117\,
            I => \N__49064\
        );

    \I__11329\ : InMux
    port map (
            O => \N__49116\,
            I => \N__49061\
        );

    \I__11328\ : Span4Mux_v
    port map (
            O => \N__49105\,
            I => \N__49058\
        );

    \I__11327\ : Span4Mux_v
    port map (
            O => \N__49102\,
            I => \N__49053\
        );

    \I__11326\ : Span4Mux_v
    port map (
            O => \N__49099\,
            I => \N__49053\
        );

    \I__11325\ : LocalMux
    port map (
            O => \N__49096\,
            I => \N__49050\
        );

    \I__11324\ : InMux
    port map (
            O => \N__49095\,
            I => \N__49046\
        );

    \I__11323\ : Span4Mux_h
    port map (
            O => \N__49088\,
            I => \N__49043\
        );

    \I__11322\ : Span4Mux_v
    port map (
            O => \N__49085\,
            I => \N__49040\
        );

    \I__11321\ : Span12Mux_v
    port map (
            O => \N__49082\,
            I => \N__49037\
        );

    \I__11320\ : Sp12to4
    port map (
            O => \N__49079\,
            I => \N__49034\
        );

    \I__11319\ : Sp12to4
    port map (
            O => \N__49076\,
            I => \N__49027\
        );

    \I__11318\ : LocalMux
    port map (
            O => \N__49073\,
            I => \N__49027\
        );

    \I__11317\ : Sp12to4
    port map (
            O => \N__49064\,
            I => \N__49027\
        );

    \I__11316\ : LocalMux
    port map (
            O => \N__49061\,
            I => \N__49024\
        );

    \I__11315\ : Span4Mux_v
    port map (
            O => \N__49058\,
            I => \N__49021\
        );

    \I__11314\ : Span4Mux_v
    port map (
            O => \N__49053\,
            I => \N__49018\
        );

    \I__11313\ : Span4Mux_v
    port map (
            O => \N__49050\,
            I => \N__49015\
        );

    \I__11312\ : IoInMux
    port map (
            O => \N__49049\,
            I => \N__49012\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__49046\,
            I => \N__49007\
        );

    \I__11310\ : Sp12to4
    port map (
            O => \N__49043\,
            I => \N__49007\
        );

    \I__11309\ : Span4Mux_h
    port map (
            O => \N__49040\,
            I => \N__49004\
        );

    \I__11308\ : Span12Mux_v
    port map (
            O => \N__49037\,
            I => \N__49001\
        );

    \I__11307\ : Span12Mux_v
    port map (
            O => \N__49034\,
            I => \N__48994\
        );

    \I__11306\ : Span12Mux_h
    port map (
            O => \N__49027\,
            I => \N__48994\
        );

    \I__11305\ : Span12Mux_h
    port map (
            O => \N__49024\,
            I => \N__48994\
        );

    \I__11304\ : Sp12to4
    port map (
            O => \N__49021\,
            I => \N__48987\
        );

    \I__11303\ : Sp12to4
    port map (
            O => \N__49018\,
            I => \N__48987\
        );

    \I__11302\ : Sp12to4
    port map (
            O => \N__49015\,
            I => \N__48987\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__49012\,
            I => \N__48984\
        );

    \I__11300\ : Span12Mux_v
    port map (
            O => \N__49007\,
            I => \N__48979\
        );

    \I__11299\ : Sp12to4
    port map (
            O => \N__49004\,
            I => \N__48979\
        );

    \I__11298\ : Span12Mux_h
    port map (
            O => \N__49001\,
            I => \N__48972\
        );

    \I__11297\ : Span12Mux_v
    port map (
            O => \N__48994\,
            I => \N__48972\
        );

    \I__11296\ : Span12Mux_h
    port map (
            O => \N__48987\,
            I => \N__48972\
        );

    \I__11295\ : IoSpan4Mux
    port map (
            O => \N__48984\,
            I => \N__48969\
        );

    \I__11294\ : Odrv12
    port map (
            O => \N__48979\,
            I => \LED3_c\
        );

    \I__11293\ : Odrv12
    port map (
            O => \N__48972\,
            I => \LED3_c\
        );

    \I__11292\ : Odrv4
    port map (
            O => \N__48969\,
            I => \LED3_c\
        );

    \I__11291\ : InMux
    port map (
            O => \N__48962\,
            I => \N__48957\
        );

    \I__11290\ : InMux
    port map (
            O => \N__48961\,
            I => \N__48953\
        );

    \I__11289\ : CEMux
    port map (
            O => \N__48960\,
            I => \N__48943\
        );

    \I__11288\ : LocalMux
    port map (
            O => \N__48957\,
            I => \N__48940\
        );

    \I__11287\ : InMux
    port map (
            O => \N__48956\,
            I => \N__48937\
        );

    \I__11286\ : LocalMux
    port map (
            O => \N__48953\,
            I => \N__48926\
        );

    \I__11285\ : InMux
    port map (
            O => \N__48952\,
            I => \N__48923\
        );

    \I__11284\ : InMux
    port map (
            O => \N__48951\,
            I => \N__48912\
        );

    \I__11283\ : InMux
    port map (
            O => \N__48950\,
            I => \N__48912\
        );

    \I__11282\ : InMux
    port map (
            O => \N__48949\,
            I => \N__48912\
        );

    \I__11281\ : InMux
    port map (
            O => \N__48948\,
            I => \N__48912\
        );

    \I__11280\ : InMux
    port map (
            O => \N__48947\,
            I => \N__48912\
        );

    \I__11279\ : InMux
    port map (
            O => \N__48946\,
            I => \N__48904\
        );

    \I__11278\ : LocalMux
    port map (
            O => \N__48943\,
            I => \N__48894\
        );

    \I__11277\ : Span4Mux_h
    port map (
            O => \N__48940\,
            I => \N__48889\
        );

    \I__11276\ : LocalMux
    port map (
            O => \N__48937\,
            I => \N__48889\
        );

    \I__11275\ : InMux
    port map (
            O => \N__48936\,
            I => \N__48872\
        );

    \I__11274\ : InMux
    port map (
            O => \N__48935\,
            I => \N__48872\
        );

    \I__11273\ : InMux
    port map (
            O => \N__48934\,
            I => \N__48872\
        );

    \I__11272\ : InMux
    port map (
            O => \N__48933\,
            I => \N__48872\
        );

    \I__11271\ : InMux
    port map (
            O => \N__48932\,
            I => \N__48872\
        );

    \I__11270\ : InMux
    port map (
            O => \N__48931\,
            I => \N__48872\
        );

    \I__11269\ : InMux
    port map (
            O => \N__48930\,
            I => \N__48872\
        );

    \I__11268\ : InMux
    port map (
            O => \N__48929\,
            I => \N__48872\
        );

    \I__11267\ : Span4Mux_v
    port map (
            O => \N__48926\,
            I => \N__48867\
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__48923\,
            I => \N__48867\
        );

    \I__11265\ : LocalMux
    port map (
            O => \N__48912\,
            I => \N__48864\
        );

    \I__11264\ : InMux
    port map (
            O => \N__48911\,
            I => \N__48853\
        );

    \I__11263\ : InMux
    port map (
            O => \N__48910\,
            I => \N__48853\
        );

    \I__11262\ : InMux
    port map (
            O => \N__48909\,
            I => \N__48853\
        );

    \I__11261\ : InMux
    port map (
            O => \N__48908\,
            I => \N__48853\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48907\,
            I => \N__48853\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__48904\,
            I => \N__48850\
        );

    \I__11258\ : InMux
    port map (
            O => \N__48903\,
            I => \N__48845\
        );

    \I__11257\ : InMux
    port map (
            O => \N__48902\,
            I => \N__48845\
        );

    \I__11256\ : InMux
    port map (
            O => \N__48901\,
            I => \N__48834\
        );

    \I__11255\ : InMux
    port map (
            O => \N__48900\,
            I => \N__48834\
        );

    \I__11254\ : InMux
    port map (
            O => \N__48899\,
            I => \N__48834\
        );

    \I__11253\ : InMux
    port map (
            O => \N__48898\,
            I => \N__48834\
        );

    \I__11252\ : InMux
    port map (
            O => \N__48897\,
            I => \N__48834\
        );

    \I__11251\ : Odrv4
    port map (
            O => \N__48894\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__11250\ : Odrv4
    port map (
            O => \N__48889\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__48872\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__11248\ : Odrv4
    port map (
            O => \N__48867\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__11247\ : Odrv4
    port map (
            O => \N__48864\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__11246\ : LocalMux
    port map (
            O => \N__48853\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__11245\ : Odrv4
    port map (
            O => \N__48850\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__11244\ : LocalMux
    port map (
            O => \N__48845\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__48834\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__11242\ : IoInMux
    port map (
            O => \N__48815\,
            I => \N__48812\
        );

    \I__11241\ : LocalMux
    port map (
            O => \N__48812\,
            I => \N__48809\
        );

    \I__11240\ : Span4Mux_s3_h
    port map (
            O => \N__48809\,
            I => \N__48806\
        );

    \I__11239\ : Span4Mux_v
    port map (
            O => \N__48806\,
            I => \N__48803\
        );

    \I__11238\ : Span4Mux_h
    port map (
            O => \N__48803\,
            I => \N__48799\
        );

    \I__11237\ : InMux
    port map (
            O => \N__48802\,
            I => \N__48796\
        );

    \I__11236\ : Odrv4
    port map (
            O => \N__48799\,
            I => \RAM_DATA_cl_5Z0Z_15\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__48796\,
            I => \RAM_DATA_cl_5Z0Z_15\
        );

    \I__11234\ : CascadeMux
    port map (
            O => \N__48791\,
            I => \N__48787\
        );

    \I__11233\ : InMux
    port map (
            O => \N__48790\,
            I => \N__48784\
        );

    \I__11232\ : InMux
    port map (
            O => \N__48787\,
            I => \N__48781\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__48784\,
            I => \N__48776\
        );

    \I__11230\ : LocalMux
    port map (
            O => \N__48781\,
            I => \N__48776\
        );

    \I__11229\ : Odrv4
    port map (
            O => \N__48776\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1\
        );

    \I__11228\ : InMux
    port map (
            O => \N__48773\,
            I => \N__48766\
        );

    \I__11227\ : InMux
    port map (
            O => \N__48772\,
            I => \N__48766\
        );

    \I__11226\ : InMux
    port map (
            O => \N__48771\,
            I => \N__48763\
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__48766\,
            I => \N__48760\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__48763\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__11223\ : Odrv4
    port map (
            O => \N__48760\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__11222\ : InMux
    port map (
            O => \N__48755\,
            I => \N__48745\
        );

    \I__11221\ : InMux
    port map (
            O => \N__48754\,
            I => \N__48745\
        );

    \I__11220\ : InMux
    port map (
            O => \N__48753\,
            I => \N__48745\
        );

    \I__11219\ : InMux
    port map (
            O => \N__48752\,
            I => \N__48742\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__48745\,
            I => \N__48739\
        );

    \I__11217\ : LocalMux
    port map (
            O => \N__48742\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__11216\ : Odrv4
    port map (
            O => \N__48739\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__11215\ : InMux
    port map (
            O => \N__48734\,
            I => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0\
        );

    \I__11214\ : InMux
    port map (
            O => \N__48731\,
            I => \N__48722\
        );

    \I__11213\ : InMux
    port map (
            O => \N__48730\,
            I => \N__48722\
        );

    \I__11212\ : InMux
    port map (
            O => \N__48729\,
            I => \N__48722\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__48722\,
            I => \N__48719\
        );

    \I__11210\ : Span4Mux_v
    port map (
            O => \N__48719\,
            I => \N__48714\
        );

    \I__11209\ : InMux
    port map (
            O => \N__48718\,
            I => \N__48708\
        );

    \I__11208\ : InMux
    port map (
            O => \N__48717\,
            I => \N__48708\
        );

    \I__11207\ : Span4Mux_h
    port map (
            O => \N__48714\,
            I => \N__48705\
        );

    \I__11206\ : InMux
    port map (
            O => \N__48713\,
            I => \N__48702\
        );

    \I__11205\ : LocalMux
    port map (
            O => \N__48708\,
            I => \N__48699\
        );

    \I__11204\ : Odrv4
    port map (
            O => \N__48705\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__11203\ : LocalMux
    port map (
            O => \N__48702\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__11202\ : Odrv4
    port map (
            O => \N__48699\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__11201\ : InMux
    port map (
            O => \N__48692\,
            I => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1\
        );

    \I__11200\ : CascadeMux
    port map (
            O => \N__48689\,
            I => \N__48686\
        );

    \I__11199\ : InMux
    port map (
            O => \N__48686\,
            I => \N__48682\
        );

    \I__11198\ : InMux
    port map (
            O => \N__48685\,
            I => \N__48679\
        );

    \I__11197\ : LocalMux
    port map (
            O => \N__48682\,
            I => \N__48676\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__48679\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__11195\ : Odrv4
    port map (
            O => \N__48676\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__11194\ : InMux
    port map (
            O => \N__48671\,
            I => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2\
        );

    \I__11193\ : InMux
    port map (
            O => \N__48668\,
            I => \N__48662\
        );

    \I__11192\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48659\
        );

    \I__11191\ : InMux
    port map (
            O => \N__48666\,
            I => \N__48656\
        );

    \I__11190\ : InMux
    port map (
            O => \N__48665\,
            I => \N__48653\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__48662\,
            I => \N__48650\
        );

    \I__11188\ : LocalMux
    port map (
            O => \N__48659\,
            I => \sCounterDACZ0Z_3\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__48656\,
            I => \sCounterDACZ0Z_3\
        );

    \I__11186\ : LocalMux
    port map (
            O => \N__48653\,
            I => \sCounterDACZ0Z_3\
        );

    \I__11185\ : Odrv4
    port map (
            O => \N__48650\,
            I => \sCounterDACZ0Z_3\
        );

    \I__11184\ : InMux
    port map (
            O => \N__48641\,
            I => un2_scounterdac_cry_2
        );

    \I__11183\ : InMux
    port map (
            O => \N__48638\,
            I => \N__48633\
        );

    \I__11182\ : InMux
    port map (
            O => \N__48637\,
            I => \N__48628\
        );

    \I__11181\ : InMux
    port map (
            O => \N__48636\,
            I => \N__48628\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__48633\,
            I => \sCounterDACZ0Z_4\
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__48628\,
            I => \sCounterDACZ0Z_4\
        );

    \I__11178\ : InMux
    port map (
            O => \N__48623\,
            I => un2_scounterdac_cry_3
        );

    \I__11177\ : CascadeMux
    port map (
            O => \N__48620\,
            I => \N__48615\
        );

    \I__11176\ : CascadeMux
    port map (
            O => \N__48619\,
            I => \N__48612\
        );

    \I__11175\ : InMux
    port map (
            O => \N__48618\,
            I => \N__48608\
        );

    \I__11174\ : InMux
    port map (
            O => \N__48615\,
            I => \N__48601\
        );

    \I__11173\ : InMux
    port map (
            O => \N__48612\,
            I => \N__48601\
        );

    \I__11172\ : InMux
    port map (
            O => \N__48611\,
            I => \N__48601\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__48608\,
            I => \sCounterDACZ0Z_5\
        );

    \I__11170\ : LocalMux
    port map (
            O => \N__48601\,
            I => \sCounterDACZ0Z_5\
        );

    \I__11169\ : InMux
    port map (
            O => \N__48596\,
            I => un2_scounterdac_cry_4
        );

    \I__11168\ : InMux
    port map (
            O => \N__48593\,
            I => \N__48588\
        );

    \I__11167\ : InMux
    port map (
            O => \N__48592\,
            I => \N__48583\
        );

    \I__11166\ : InMux
    port map (
            O => \N__48591\,
            I => \N__48583\
        );

    \I__11165\ : LocalMux
    port map (
            O => \N__48588\,
            I => \sCounterDACZ0Z_6\
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__48583\,
            I => \sCounterDACZ0Z_6\
        );

    \I__11163\ : InMux
    port map (
            O => \N__48578\,
            I => \N__48575\
        );

    \I__11162\ : LocalMux
    port map (
            O => \N__48575\,
            I => \un2_scounterdac_cry_5_THRU_CO\
        );

    \I__11161\ : InMux
    port map (
            O => \N__48572\,
            I => un2_scounterdac_cry_5
        );

    \I__11160\ : InMux
    port map (
            O => \N__48569\,
            I => \N__48565\
        );

    \I__11159\ : InMux
    port map (
            O => \N__48568\,
            I => \N__48562\
        );

    \I__11158\ : LocalMux
    port map (
            O => \N__48565\,
            I => \sCounterDACZ0Z_7\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__48562\,
            I => \sCounterDACZ0Z_7\
        );

    \I__11156\ : InMux
    port map (
            O => \N__48557\,
            I => un2_scounterdac_cry_6
        );

    \I__11155\ : InMux
    port map (
            O => \N__48554\,
            I => \N__48550\
        );

    \I__11154\ : InMux
    port map (
            O => \N__48553\,
            I => \N__48547\
        );

    \I__11153\ : LocalMux
    port map (
            O => \N__48550\,
            I => \N__48544\
        );

    \I__11152\ : LocalMux
    port map (
            O => \N__48547\,
            I => \N_30_mux\
        );

    \I__11151\ : Odrv4
    port map (
            O => \N__48544\,
            I => \N_30_mux\
        );

    \I__11150\ : InMux
    port map (
            O => \N__48539\,
            I => \N__48536\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__48536\,
            I => \N__48530\
        );

    \I__11148\ : InMux
    port map (
            O => \N__48535\,
            I => \N__48527\
        );

    \I__11147\ : InMux
    port map (
            O => \N__48534\,
            I => \N__48522\
        );

    \I__11146\ : InMux
    port map (
            O => \N__48533\,
            I => \N__48522\
        );

    \I__11145\ : Odrv12
    port map (
            O => \N__48530\,
            I => \sCounterDACZ0Z_8\
        );

    \I__11144\ : LocalMux
    port map (
            O => \N__48527\,
            I => \sCounterDACZ0Z_8\
        );

    \I__11143\ : LocalMux
    port map (
            O => \N__48522\,
            I => \sCounterDACZ0Z_8\
        );

    \I__11142\ : InMux
    port map (
            O => \N__48515\,
            I => un2_scounterdac_cry_7
        );

    \I__11141\ : InMux
    port map (
            O => \N__48512\,
            I => \bfn_20_11_0_\
        );

    \I__11140\ : CascadeMux
    port map (
            O => \N__48509\,
            I => \N__48506\
        );

    \I__11139\ : InMux
    port map (
            O => \N__48506\,
            I => \N__48502\
        );

    \I__11138\ : InMux
    port map (
            O => \N__48505\,
            I => \N__48499\
        );

    \I__11137\ : LocalMux
    port map (
            O => \N__48502\,
            I => \N__48496\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__48499\,
            I => \sCounterDACZ0Z_9\
        );

    \I__11135\ : Odrv4
    port map (
            O => \N__48496\,
            I => \sCounterDACZ0Z_9\
        );

    \I__11134\ : ClkMux
    port map (
            O => \N__48491\,
            I => \N__48347\
        );

    \I__11133\ : ClkMux
    port map (
            O => \N__48490\,
            I => \N__48347\
        );

    \I__11132\ : ClkMux
    port map (
            O => \N__48489\,
            I => \N__48347\
        );

    \I__11131\ : ClkMux
    port map (
            O => \N__48488\,
            I => \N__48347\
        );

    \I__11130\ : ClkMux
    port map (
            O => \N__48487\,
            I => \N__48347\
        );

    \I__11129\ : ClkMux
    port map (
            O => \N__48486\,
            I => \N__48347\
        );

    \I__11128\ : ClkMux
    port map (
            O => \N__48485\,
            I => \N__48347\
        );

    \I__11127\ : ClkMux
    port map (
            O => \N__48484\,
            I => \N__48347\
        );

    \I__11126\ : ClkMux
    port map (
            O => \N__48483\,
            I => \N__48347\
        );

    \I__11125\ : ClkMux
    port map (
            O => \N__48482\,
            I => \N__48347\
        );

    \I__11124\ : ClkMux
    port map (
            O => \N__48481\,
            I => \N__48347\
        );

    \I__11123\ : ClkMux
    port map (
            O => \N__48480\,
            I => \N__48347\
        );

    \I__11122\ : ClkMux
    port map (
            O => \N__48479\,
            I => \N__48347\
        );

    \I__11121\ : ClkMux
    port map (
            O => \N__48478\,
            I => \N__48347\
        );

    \I__11120\ : ClkMux
    port map (
            O => \N__48477\,
            I => \N__48347\
        );

    \I__11119\ : ClkMux
    port map (
            O => \N__48476\,
            I => \N__48347\
        );

    \I__11118\ : ClkMux
    port map (
            O => \N__48475\,
            I => \N__48347\
        );

    \I__11117\ : ClkMux
    port map (
            O => \N__48474\,
            I => \N__48347\
        );

    \I__11116\ : ClkMux
    port map (
            O => \N__48473\,
            I => \N__48347\
        );

    \I__11115\ : ClkMux
    port map (
            O => \N__48472\,
            I => \N__48347\
        );

    \I__11114\ : ClkMux
    port map (
            O => \N__48471\,
            I => \N__48347\
        );

    \I__11113\ : ClkMux
    port map (
            O => \N__48470\,
            I => \N__48347\
        );

    \I__11112\ : ClkMux
    port map (
            O => \N__48469\,
            I => \N__48347\
        );

    \I__11111\ : ClkMux
    port map (
            O => \N__48468\,
            I => \N__48347\
        );

    \I__11110\ : ClkMux
    port map (
            O => \N__48467\,
            I => \N__48347\
        );

    \I__11109\ : ClkMux
    port map (
            O => \N__48466\,
            I => \N__48347\
        );

    \I__11108\ : ClkMux
    port map (
            O => \N__48465\,
            I => \N__48347\
        );

    \I__11107\ : ClkMux
    port map (
            O => \N__48464\,
            I => \N__48347\
        );

    \I__11106\ : ClkMux
    port map (
            O => \N__48463\,
            I => \N__48347\
        );

    \I__11105\ : ClkMux
    port map (
            O => \N__48462\,
            I => \N__48347\
        );

    \I__11104\ : ClkMux
    port map (
            O => \N__48461\,
            I => \N__48347\
        );

    \I__11103\ : ClkMux
    port map (
            O => \N__48460\,
            I => \N__48347\
        );

    \I__11102\ : ClkMux
    port map (
            O => \N__48459\,
            I => \N__48347\
        );

    \I__11101\ : ClkMux
    port map (
            O => \N__48458\,
            I => \N__48347\
        );

    \I__11100\ : ClkMux
    port map (
            O => \N__48457\,
            I => \N__48347\
        );

    \I__11099\ : ClkMux
    port map (
            O => \N__48456\,
            I => \N__48347\
        );

    \I__11098\ : ClkMux
    port map (
            O => \N__48455\,
            I => \N__48347\
        );

    \I__11097\ : ClkMux
    port map (
            O => \N__48454\,
            I => \N__48347\
        );

    \I__11096\ : ClkMux
    port map (
            O => \N__48453\,
            I => \N__48347\
        );

    \I__11095\ : ClkMux
    port map (
            O => \N__48452\,
            I => \N__48347\
        );

    \I__11094\ : ClkMux
    port map (
            O => \N__48451\,
            I => \N__48347\
        );

    \I__11093\ : ClkMux
    port map (
            O => \N__48450\,
            I => \N__48347\
        );

    \I__11092\ : ClkMux
    port map (
            O => \N__48449\,
            I => \N__48347\
        );

    \I__11091\ : ClkMux
    port map (
            O => \N__48448\,
            I => \N__48347\
        );

    \I__11090\ : ClkMux
    port map (
            O => \N__48447\,
            I => \N__48347\
        );

    \I__11089\ : ClkMux
    port map (
            O => \N__48446\,
            I => \N__48347\
        );

    \I__11088\ : ClkMux
    port map (
            O => \N__48445\,
            I => \N__48347\
        );

    \I__11087\ : ClkMux
    port map (
            O => \N__48444\,
            I => \N__48347\
        );

    \I__11086\ : GlobalMux
    port map (
            O => \N__48347\,
            I => \N__48344\
        );

    \I__11085\ : gio2CtrlBuf
    port map (
            O => \N__48344\,
            I => pll_clk64_0_g
        );

    \I__11084\ : InMux
    port map (
            O => \N__48341\,
            I => \N__48338\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__48338\,
            I => \N__48335\
        );

    \I__11082\ : Span12Mux_h
    port map (
            O => \N__48335\,
            I => \N__48332\
        );

    \I__11081\ : Odrv12
    port map (
            O => \N__48332\,
            I => \spi_slave_inst.un23_i_ssn_3\
        );

    \I__11080\ : InMux
    port map (
            O => \N__48329\,
            I => \N__48325\
        );

    \I__11079\ : InMux
    port map (
            O => \N__48328\,
            I => \N__48321\
        );

    \I__11078\ : LocalMux
    port map (
            O => \N__48325\,
            I => \N__48318\
        );

    \I__11077\ : InMux
    port map (
            O => \N__48324\,
            I => \N__48315\
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__48321\,
            I => \N__48310\
        );

    \I__11075\ : Span12Mux_h
    port map (
            O => \N__48318\,
            I => \N__48310\
        );

    \I__11074\ : LocalMux
    port map (
            O => \N__48315\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4\
        );

    \I__11073\ : Odrv12
    port map (
            O => \N__48310\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4\
        );

    \I__11072\ : InMux
    port map (
            O => \N__48305\,
            I => \N__48300\
        );

    \I__11071\ : InMux
    port map (
            O => \N__48304\,
            I => \N__48297\
        );

    \I__11070\ : InMux
    port map (
            O => \N__48303\,
            I => \N__48294\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__48300\,
            I => \N__48289\
        );

    \I__11068\ : LocalMux
    port map (
            O => \N__48297\,
            I => \N__48289\
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__48294\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3\
        );

    \I__11066\ : Odrv12
    port map (
            O => \N__48289\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3\
        );

    \I__11065\ : InMux
    port map (
            O => \N__48284\,
            I => \N__48281\
        );

    \I__11064\ : LocalMux
    port map (
            O => \N__48281\,
            I => \N__48278\
        );

    \I__11063\ : Span12Mux_v
    port map (
            O => \N__48278\,
            I => \N__48275\
        );

    \I__11062\ : Span12Mux_h
    port map (
            O => \N__48275\,
            I => \N__48272\
        );

    \I__11061\ : Span12Mux_v
    port map (
            O => \N__48272\,
            I => \N__48269\
        );

    \I__11060\ : Odrv12
    port map (
            O => \N__48269\,
            I => \spi_slave_inst.rx_done_pos_sclk_iZ0\
        );

    \I__11059\ : ClkMux
    port map (
            O => \N__48266\,
            I => \N__48242\
        );

    \I__11058\ : ClkMux
    port map (
            O => \N__48265\,
            I => \N__48242\
        );

    \I__11057\ : ClkMux
    port map (
            O => \N__48264\,
            I => \N__48242\
        );

    \I__11056\ : ClkMux
    port map (
            O => \N__48263\,
            I => \N__48242\
        );

    \I__11055\ : ClkMux
    port map (
            O => \N__48262\,
            I => \N__48242\
        );

    \I__11054\ : ClkMux
    port map (
            O => \N__48261\,
            I => \N__48242\
        );

    \I__11053\ : ClkMux
    port map (
            O => \N__48260\,
            I => \N__48242\
        );

    \I__11052\ : ClkMux
    port map (
            O => \N__48259\,
            I => \N__48242\
        );

    \I__11051\ : GlobalMux
    port map (
            O => \N__48242\,
            I => \N__48239\
        );

    \I__11050\ : gio2CtrlBuf
    port map (
            O => \N__48239\,
            I => spi_sclk_g
        );

    \I__11049\ : CEMux
    port map (
            O => \N__48236\,
            I => \N__48233\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__48233\,
            I => \N__48228\
        );

    \I__11047\ : CEMux
    port map (
            O => \N__48232\,
            I => \N__48225\
        );

    \I__11046\ : CEMux
    port map (
            O => \N__48231\,
            I => \N__48222\
        );

    \I__11045\ : Span4Mux_h
    port map (
            O => \N__48228\,
            I => \N__48219\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__48225\,
            I => \N__48216\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__48222\,
            I => \N__48213\
        );

    \I__11042\ : Span4Mux_v
    port map (
            O => \N__48219\,
            I => \N__48210\
        );

    \I__11041\ : Span4Mux_v
    port map (
            O => \N__48216\,
            I => \N__48207\
        );

    \I__11040\ : Span12Mux_h
    port map (
            O => \N__48213\,
            I => \N__48204\
        );

    \I__11039\ : Span4Mux_v
    port map (
            O => \N__48210\,
            I => \N__48201\
        );

    \I__11038\ : Span4Mux_h
    port map (
            O => \N__48207\,
            I => \N__48198\
        );

    \I__11037\ : Odrv12
    port map (
            O => \N__48204\,
            I => \spi_slave_inst.spi_cs_iZ0\
        );

    \I__11036\ : Odrv4
    port map (
            O => \N__48201\,
            I => \spi_slave_inst.spi_cs_iZ0\
        );

    \I__11035\ : Odrv4
    port map (
            O => \N__48198\,
            I => \spi_slave_inst.spi_cs_iZ0\
        );

    \I__11034\ : CascadeMux
    port map (
            O => \N__48191\,
            I => \N_23_mux_cascade_\
        );

    \I__11033\ : CascadeMux
    port map (
            O => \N__48188\,
            I => \N_25_mux_cascade_\
        );

    \I__11032\ : InMux
    port map (
            O => \N__48185\,
            I => \N__48182\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__48182\,
            I => m15_1
        );

    \I__11030\ : IoInMux
    port map (
            O => \N__48179\,
            I => \N__48176\
        );

    \I__11029\ : LocalMux
    port map (
            O => \N__48176\,
            I => \N__48173\
        );

    \I__11028\ : IoSpan4Mux
    port map (
            O => \N__48173\,
            I => \N__48170\
        );

    \I__11027\ : Span4Mux_s0_h
    port map (
            O => \N__48170\,
            I => \N__48167\
        );

    \I__11026\ : Span4Mux_h
    port map (
            O => \N__48167\,
            I => \N__48164\
        );

    \I__11025\ : Odrv4
    port map (
            O => \N__48164\,
            I => op_eq_scounterdac10
        );

    \I__11024\ : InMux
    port map (
            O => \N__48161\,
            I => \N__48158\
        );

    \I__11023\ : LocalMux
    port map (
            O => \N__48158\,
            I => m8_2
        );

    \I__11022\ : InMux
    port map (
            O => \N__48155\,
            I => \N__48152\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__48152\,
            I => \N_23_mux\
        );

    \I__11020\ : CascadeMux
    port map (
            O => \N__48149\,
            I => \N_30_mux_cascade_\
        );

    \I__11019\ : InMux
    port map (
            O => \N__48146\,
            I => \N__48143\
        );

    \I__11018\ : LocalMux
    port map (
            O => \N__48143\,
            I => \N_25_mux\
        );

    \I__11017\ : InMux
    port map (
            O => \N__48140\,
            I => \N__48137\
        );

    \I__11016\ : LocalMux
    port map (
            O => \N__48137\,
            I => \N__48134\
        );

    \I__11015\ : Odrv12
    port map (
            O => \N__48134\,
            I => \N_32_mux\
        );

    \I__11014\ : InMux
    port map (
            O => \N__48131\,
            I => \N__48119\
        );

    \I__11013\ : InMux
    port map (
            O => \N__48130\,
            I => \N__48119\
        );

    \I__11012\ : InMux
    port map (
            O => \N__48129\,
            I => \N__48119\
        );

    \I__11011\ : InMux
    port map (
            O => \N__48128\,
            I => \N__48116\
        );

    \I__11010\ : InMux
    port map (
            O => \N__48127\,
            I => \N__48113\
        );

    \I__11009\ : InMux
    port map (
            O => \N__48126\,
            I => \N__48110\
        );

    \I__11008\ : LocalMux
    port map (
            O => \N__48119\,
            I => \N__48103\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__48116\,
            I => \N__48103\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__48113\,
            I => \N__48103\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__48110\,
            I => \sCounterDACZ0Z_0\
        );

    \I__11004\ : Odrv12
    port map (
            O => \N__48103\,
            I => \sCounterDACZ0Z_0\
        );

    \I__11003\ : CascadeMux
    port map (
            O => \N__48098\,
            I => \N__48094\
        );

    \I__11002\ : CascadeMux
    port map (
            O => \N__48097\,
            I => \N__48091\
        );

    \I__11001\ : InMux
    port map (
            O => \N__48094\,
            I => \N__48086\
        );

    \I__11000\ : InMux
    port map (
            O => \N__48091\,
            I => \N__48079\
        );

    \I__10999\ : InMux
    port map (
            O => \N__48090\,
            I => \N__48079\
        );

    \I__10998\ : InMux
    port map (
            O => \N__48089\,
            I => \N__48079\
        );

    \I__10997\ : LocalMux
    port map (
            O => \N__48086\,
            I => \sCounterDACZ0Z_1\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__48079\,
            I => \sCounterDACZ0Z_1\
        );

    \I__10995\ : InMux
    port map (
            O => \N__48074\,
            I => \N__48070\
        );

    \I__10994\ : InMux
    port map (
            O => \N__48073\,
            I => \N__48067\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__48070\,
            I => \sCounterDACZ0Z_2\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__48067\,
            I => \sCounterDACZ0Z_2\
        );

    \I__10991\ : InMux
    port map (
            O => \N__48062\,
            I => un2_scounterdac_cry_1
        );

    \I__10990\ : CascadeMux
    port map (
            O => \N__48059\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_\
        );

    \I__10989\ : InMux
    port map (
            O => \N__48056\,
            I => \N__48053\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__48053\,
            I => \N__48048\
        );

    \I__10987\ : InMux
    port map (
            O => \N__48052\,
            I => \N__48045\
        );

    \I__10986\ : InMux
    port map (
            O => \N__48051\,
            I => \N__48042\
        );

    \I__10985\ : Span4Mux_v
    port map (
            O => \N__48048\,
            I => \N__48038\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__48045\,
            I => \N__48033\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__48042\,
            I => \N__48033\
        );

    \I__10982\ : InMux
    port map (
            O => \N__48041\,
            I => \N__48029\
        );

    \I__10981\ : Span4Mux_v
    port map (
            O => \N__48038\,
            I => \N__48024\
        );

    \I__10980\ : Span4Mux_v
    port map (
            O => \N__48033\,
            I => \N__48024\
        );

    \I__10979\ : InMux
    port map (
            O => \N__48032\,
            I => \N__48021\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__48029\,
            I => \N__48018\
        );

    \I__10977\ : Span4Mux_h
    port map (
            O => \N__48024\,
            I => \N__48015\
        );

    \I__10976\ : LocalMux
    port map (
            O => \N__48021\,
            I => \N__48012\
        );

    \I__10975\ : Span4Mux_h
    port map (
            O => \N__48018\,
            I => \N__48008\
        );

    \I__10974\ : Span4Mux_h
    port map (
            O => \N__48015\,
            I => \N__48001\
        );

    \I__10973\ : Span4Mux_v
    port map (
            O => \N__48012\,
            I => \N__48001\
        );

    \I__10972\ : InMux
    port map (
            O => \N__48011\,
            I => \N__47998\
        );

    \I__10971\ : Span4Mux_h
    port map (
            O => \N__48008\,
            I => \N__47995\
        );

    \I__10970\ : InMux
    port map (
            O => \N__48007\,
            I => \N__47992\
        );

    \I__10969\ : InMux
    port map (
            O => \N__48006\,
            I => \N__47989\
        );

    \I__10968\ : Span4Mux_h
    port map (
            O => \N__48001\,
            I => \N__47984\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__47998\,
            I => \N__47984\
        );

    \I__10966\ : Sp12to4
    port map (
            O => \N__47995\,
            I => \N__47977\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__47992\,
            I => \N__47977\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__47989\,
            I => \N__47977\
        );

    \I__10963\ : Span4Mux_h
    port map (
            O => \N__47984\,
            I => \N__47974\
        );

    \I__10962\ : Span12Mux_v
    port map (
            O => \N__47977\,
            I => \N__47971\
        );

    \I__10961\ : Span4Mux_v
    port map (
            O => \N__47974\,
            I => \N__47968\
        );

    \I__10960\ : Span12Mux_h
    port map (
            O => \N__47971\,
            I => \N__47965\
        );

    \I__10959\ : Sp12to4
    port map (
            O => \N__47968\,
            I => \N__47962\
        );

    \I__10958\ : Odrv12
    port map (
            O => \N__47965\,
            I => spi_select_c
        );

    \I__10957\ : Odrv12
    port map (
            O => \N__47962\,
            I => spi_select_c
        );

    \I__10956\ : InMux
    port map (
            O => \N__47957\,
            I => \N__47951\
        );

    \I__10955\ : InMux
    port map (
            O => \N__47956\,
            I => \N__47951\
        );

    \I__10954\ : LocalMux
    port map (
            O => \N__47951\,
            I => \N__47948\
        );

    \I__10953\ : Span4Mux_h
    port map (
            O => \N__47948\,
            I => \N__47944\
        );

    \I__10952\ : InMux
    port map (
            O => \N__47947\,
            I => \N__47941\
        );

    \I__10951\ : Span4Mux_h
    port map (
            O => \N__47944\,
            I => \N__47936\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__47941\,
            I => \N__47936\
        );

    \I__10949\ : Span4Mux_v
    port map (
            O => \N__47936\,
            I => \N__47933\
        );

    \I__10948\ : Span4Mux_h
    port map (
            O => \N__47933\,
            I => \N__47930\
        );

    \I__10947\ : Span4Mux_v
    port map (
            O => \N__47930\,
            I => \N__47925\
        );

    \I__10946\ : InMux
    port map (
            O => \N__47929\,
            I => \N__47922\
        );

    \I__10945\ : InMux
    port map (
            O => \N__47928\,
            I => \N__47919\
        );

    \I__10944\ : Sp12to4
    port map (
            O => \N__47925\,
            I => \N__47912\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__47922\,
            I => \N__47912\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__47919\,
            I => \N__47912\
        );

    \I__10941\ : Span12Mux_v
    port map (
            O => \N__47912\,
            I => \N__47909\
        );

    \I__10940\ : Odrv12
    port map (
            O => \N__47909\,
            I => spi_cs_ft_c
        );

    \I__10939\ : CascadeMux
    port map (
            O => \N__47906\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_\
        );

    \I__10938\ : InMux
    port map (
            O => \N__47903\,
            I => \N__47900\
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__47900\,
            I => \N__47897\
        );

    \I__10936\ : Span4Mux_v
    port map (
            O => \N__47897\,
            I => \N__47894\
        );

    \I__10935\ : Span4Mux_h
    port map (
            O => \N__47894\,
            I => \N__47889\
        );

    \I__10934\ : InMux
    port map (
            O => \N__47893\,
            I => \N__47882\
        );

    \I__10933\ : InMux
    port map (
            O => \N__47892\,
            I => \N__47882\
        );

    \I__10932\ : Span4Mux_h
    port map (
            O => \N__47889\,
            I => \N__47879\
        );

    \I__10931\ : InMux
    port map (
            O => \N__47888\,
            I => \N__47876\
        );

    \I__10930\ : InMux
    port map (
            O => \N__47887\,
            I => \N__47873\
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__47882\,
            I => \N__47870\
        );

    \I__10928\ : Span4Mux_v
    port map (
            O => \N__47879\,
            I => \N__47867\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__47876\,
            I => \N__47864\
        );

    \I__10926\ : LocalMux
    port map (
            O => \N__47873\,
            I => \N__47861\
        );

    \I__10925\ : Span12Mux_v
    port map (
            O => \N__47870\,
            I => \N__47858\
        );

    \I__10924\ : Sp12to4
    port map (
            O => \N__47867\,
            I => \N__47855\
        );

    \I__10923\ : Span4Mux_h
    port map (
            O => \N__47864\,
            I => \N__47852\
        );

    \I__10922\ : Span4Mux_h
    port map (
            O => \N__47861\,
            I => \N__47849\
        );

    \I__10921\ : Span12Mux_v
    port map (
            O => \N__47858\,
            I => \N__47846\
        );

    \I__10920\ : Span12Mux_s6_h
    port map (
            O => \N__47855\,
            I => \N__47839\
        );

    \I__10919\ : Sp12to4
    port map (
            O => \N__47852\,
            I => \N__47839\
        );

    \I__10918\ : Sp12to4
    port map (
            O => \N__47849\,
            I => \N__47839\
        );

    \I__10917\ : Span12Mux_h
    port map (
            O => \N__47846\,
            I => \N__47834\
        );

    \I__10916\ : Span12Mux_v
    port map (
            O => \N__47839\,
            I => \N__47834\
        );

    \I__10915\ : Odrv12
    port map (
            O => \N__47834\,
            I => spi_cs_rpi_c
        );

    \I__10914\ : InMux
    port map (
            O => \N__47831\,
            I => \N__47828\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__47828\,
            I => \N__47825\
        );

    \I__10912\ : Span4Mux_v
    port map (
            O => \N__47825\,
            I => \N__47822\
        );

    \I__10911\ : Span4Mux_v
    port map (
            O => \N__47822\,
            I => \N__47819\
        );

    \I__10910\ : Odrv4
    port map (
            O => \N__47819\,
            I => \spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1\
        );

    \I__10909\ : InMux
    port map (
            O => \N__47816\,
            I => \N__47813\
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__47813\,
            I => \N__47810\
        );

    \I__10907\ : Span4Mux_v
    port map (
            O => \N__47810\,
            I => \N__47807\
        );

    \I__10906\ : Span4Mux_v
    port map (
            O => \N__47807\,
            I => \N__47804\
        );

    \I__10905\ : Odrv4
    port map (
            O => \N__47804\,
            I => \spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3\
        );

    \I__10904\ : CascadeMux
    port map (
            O => \N__47801\,
            I => \spi_slave_inst.N_1393_cascade_\
        );

    \I__10903\ : IoInMux
    port map (
            O => \N__47798\,
            I => \N__47795\
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__47795\,
            I => \N__47792\
        );

    \I__10901\ : IoSpan4Mux
    port map (
            O => \N__47792\,
            I => \N__47789\
        );

    \I__10900\ : Span4Mux_s2_h
    port map (
            O => \N__47789\,
            I => \N__47786\
        );

    \I__10899\ : Span4Mux_v
    port map (
            O => \N__47786\,
            I => \N__47783\
        );

    \I__10898\ : Sp12to4
    port map (
            O => \N__47783\,
            I => \N__47779\
        );

    \I__10897\ : InMux
    port map (
            O => \N__47782\,
            I => \N__47776\
        );

    \I__10896\ : Span12Mux_h
    port map (
            O => \N__47779\,
            I => \N__47773\
        );

    \I__10895\ : LocalMux
    port map (
            O => \N__47776\,
            I => \N__47770\
        );

    \I__10894\ : Odrv12
    port map (
            O => \N__47773\,
            I => spi_miso
        );

    \I__10893\ : Odrv12
    port map (
            O => \N__47770\,
            I => spi_miso
        );

    \I__10892\ : InMux
    port map (
            O => \N__47765\,
            I => \N__47762\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__47762\,
            I => \N__47759\
        );

    \I__10890\ : Span4Mux_v
    port map (
            O => \N__47759\,
            I => \N__47756\
        );

    \I__10889\ : Odrv4
    port map (
            O => \N__47756\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_0\
        );

    \I__10888\ : InMux
    port map (
            O => \N__47753\,
            I => \N__47750\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__47750\,
            I => \N__47747\
        );

    \I__10886\ : Span4Mux_v
    port map (
            O => \N__47747\,
            I => \N__47744\
        );

    \I__10885\ : Odrv4
    port map (
            O => \N__47744\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_4\
        );

    \I__10884\ : CascadeMux
    port map (
            O => \N__47741\,
            I => \spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0_cascade_\
        );

    \I__10883\ : InMux
    port map (
            O => \N__47738\,
            I => \N__47735\
        );

    \I__10882\ : LocalMux
    port map (
            O => \N__47735\,
            I => \N__47732\
        );

    \I__10881\ : Span4Mux_v
    port map (
            O => \N__47732\,
            I => \N__47729\
        );

    \I__10880\ : Span4Mux_v
    port map (
            O => \N__47729\,
            I => \N__47726\
        );

    \I__10879\ : Odrv4
    port map (
            O => \N__47726\,
            I => \spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2\
        );

    \I__10878\ : InMux
    port map (
            O => \N__47723\,
            I => \N__47720\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__47720\,
            I => \spi_slave_inst.N_1396\
        );

    \I__10876\ : InMux
    port map (
            O => \N__47717\,
            I => \N__47714\
        );

    \I__10875\ : LocalMux
    port map (
            O => \N__47714\,
            I => \N__47711\
        );

    \I__10874\ : Span12Mux_h
    port map (
            O => \N__47711\,
            I => \N__47708\
        );

    \I__10873\ : Span12Mux_h
    port map (
            O => \N__47708\,
            I => \N__47705\
        );

    \I__10872\ : Odrv12
    port map (
            O => \N__47705\,
            I => \ADC7_c\
        );

    \I__10871\ : IoInMux
    port map (
            O => \N__47702\,
            I => \N__47699\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__47699\,
            I => \N__47696\
        );

    \I__10869\ : IoSpan4Mux
    port map (
            O => \N__47696\,
            I => \N__47693\
        );

    \I__10868\ : Span4Mux_s2_h
    port map (
            O => \N__47693\,
            I => \N__47690\
        );

    \I__10867\ : Sp12to4
    port map (
            O => \N__47690\,
            I => \N__47687\
        );

    \I__10866\ : Span12Mux_s9_h
    port map (
            O => \N__47687\,
            I => \N__47684\
        );

    \I__10865\ : Span12Mux_v
    port map (
            O => \N__47684\,
            I => \N__47681\
        );

    \I__10864\ : Odrv12
    port map (
            O => \N__47681\,
            I => \RAM_DATA_1Z0Z_8\
        );

    \I__10863\ : InMux
    port map (
            O => \N__47678\,
            I => \N__47675\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__47675\,
            I => \N__47672\
        );

    \I__10861\ : Span4Mux_v
    port map (
            O => \N__47672\,
            I => \N__47669\
        );

    \I__10860\ : Sp12to4
    port map (
            O => \N__47669\,
            I => \N__47666\
        );

    \I__10859\ : Span12Mux_h
    port map (
            O => \N__47666\,
            I => \N__47663\
        );

    \I__10858\ : Span12Mux_h
    port map (
            O => \N__47663\,
            I => \N__47660\
        );

    \I__10857\ : Odrv12
    port map (
            O => \N__47660\,
            I => \ADC8_c\
        );

    \I__10856\ : IoInMux
    port map (
            O => \N__47657\,
            I => \N__47654\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__47654\,
            I => \N__47651\
        );

    \I__10854\ : IoSpan4Mux
    port map (
            O => \N__47651\,
            I => \N__47648\
        );

    \I__10853\ : IoSpan4Mux
    port map (
            O => \N__47648\,
            I => \N__47645\
        );

    \I__10852\ : Sp12to4
    port map (
            O => \N__47645\,
            I => \N__47642\
        );

    \I__10851\ : Span12Mux_s9_h
    port map (
            O => \N__47642\,
            I => \N__47639\
        );

    \I__10850\ : Odrv12
    port map (
            O => \N__47639\,
            I => \RAM_DATA_1Z0Z_9\
        );

    \I__10849\ : InMux
    port map (
            O => \N__47636\,
            I => \N__47633\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__47633\,
            I => \N__47630\
        );

    \I__10847\ : Span12Mux_h
    port map (
            O => \N__47630\,
            I => \N__47627\
        );

    \I__10846\ : Span12Mux_h
    port map (
            O => \N__47627\,
            I => \N__47624\
        );

    \I__10845\ : Span12Mux_v
    port map (
            O => \N__47624\,
            I => \N__47621\
        );

    \I__10844\ : Odrv12
    port map (
            O => \N__47621\,
            I => top_tour2_c
        );

    \I__10843\ : IoInMux
    port map (
            O => \N__47618\,
            I => \N__47615\
        );

    \I__10842\ : LocalMux
    port map (
            O => \N__47615\,
            I => \N__47612\
        );

    \I__10841\ : IoSpan4Mux
    port map (
            O => \N__47612\,
            I => \N__47609\
        );

    \I__10840\ : Sp12to4
    port map (
            O => \N__47609\,
            I => \N__47606\
        );

    \I__10839\ : Span12Mux_s9_h
    port map (
            O => \N__47606\,
            I => \N__47603\
        );

    \I__10838\ : Odrv12
    port map (
            O => \N__47603\,
            I => \RAM_DATA_1Z0Z_12\
        );

    \I__10837\ : IoInMux
    port map (
            O => \N__47600\,
            I => \N__47597\
        );

    \I__10836\ : LocalMux
    port map (
            O => \N__47597\,
            I => \N__47594\
        );

    \I__10835\ : Span4Mux_s0_v
    port map (
            O => \N__47594\,
            I => \N__47591\
        );

    \I__10834\ : Span4Mux_v
    port map (
            O => \N__47591\,
            I => \N__47588\
        );

    \I__10833\ : Span4Mux_v
    port map (
            O => \N__47588\,
            I => \N__47585\
        );

    \I__10832\ : Odrv4
    port map (
            O => \N__47585\,
            I => spi_miso_ft_c
        );

    \I__10831\ : InMux
    port map (
            O => \N__47582\,
            I => \N__47579\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__47579\,
            I => \N__47576\
        );

    \I__10829\ : Span4Mux_h
    port map (
            O => \N__47576\,
            I => \N__47573\
        );

    \I__10828\ : Span4Mux_h
    port map (
            O => \N__47573\,
            I => \N__47570\
        );

    \I__10827\ : Odrv4
    port map (
            O => \N__47570\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_8\
        );

    \I__10826\ : InMux
    port map (
            O => \N__47567\,
            I => \N__47564\
        );

    \I__10825\ : LocalMux
    port map (
            O => \N__47564\,
            I => \N__47561\
        );

    \I__10824\ : Span12Mux_h
    port map (
            O => \N__47561\,
            I => \N__47558\
        );

    \I__10823\ : Odrv12
    port map (
            O => \N__47558\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8\
        );

    \I__10822\ : InMux
    port map (
            O => \N__47555\,
            I => \N__47549\
        );

    \I__10821\ : InMux
    port map (
            O => \N__47554\,
            I => \N__47549\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__47549\,
            I => \N__47546\
        );

    \I__10819\ : Span4Mux_v
    port map (
            O => \N__47546\,
            I => \N__47542\
        );

    \I__10818\ : CascadeMux
    port map (
            O => \N__47545\,
            I => \N__47539\
        );

    \I__10817\ : Sp12to4
    port map (
            O => \N__47542\,
            I => \N__47536\
        );

    \I__10816\ : InMux
    port map (
            O => \N__47539\,
            I => \N__47533\
        );

    \I__10815\ : Span12Mux_h
    port map (
            O => \N__47536\,
            I => \N__47530\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__47533\,
            I => \sDAC_spi_startZ0\
        );

    \I__10813\ : Odrv12
    port map (
            O => \N__47530\,
            I => \sDAC_spi_startZ0\
        );

    \I__10812\ : InMux
    port map (
            O => \N__47525\,
            I => \N__47522\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__47522\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_5\
        );

    \I__10810\ : InMux
    port map (
            O => \N__47519\,
            I => \N__47516\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__47516\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_5\
        );

    \I__10808\ : InMux
    port map (
            O => \N__47513\,
            I => \N__47508\
        );

    \I__10807\ : InMux
    port map (
            O => \N__47512\,
            I => \N__47503\
        );

    \I__10806\ : InMux
    port map (
            O => \N__47511\,
            I => \N__47493\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__47508\,
            I => \N__47489\
        );

    \I__10804\ : InMux
    port map (
            O => \N__47507\,
            I => \N__47486\
        );

    \I__10803\ : InMux
    port map (
            O => \N__47506\,
            I => \N__47477\
        );

    \I__10802\ : LocalMux
    port map (
            O => \N__47503\,
            I => \N__47474\
        );

    \I__10801\ : InMux
    port map (
            O => \N__47502\,
            I => \N__47471\
        );

    \I__10800\ : InMux
    port map (
            O => \N__47501\,
            I => \N__47468\
        );

    \I__10799\ : InMux
    port map (
            O => \N__47500\,
            I => \N__47465\
        );

    \I__10798\ : InMux
    port map (
            O => \N__47499\,
            I => \N__47462\
        );

    \I__10797\ : InMux
    port map (
            O => \N__47498\,
            I => \N__47454\
        );

    \I__10796\ : InMux
    port map (
            O => \N__47497\,
            I => \N__47451\
        );

    \I__10795\ : InMux
    port map (
            O => \N__47496\,
            I => \N__47448\
        );

    \I__10794\ : LocalMux
    port map (
            O => \N__47493\,
            I => \N__47443\
        );

    \I__10793\ : InMux
    port map (
            O => \N__47492\,
            I => \N__47440\
        );

    \I__10792\ : Span4Mux_v
    port map (
            O => \N__47489\,
            I => \N__47432\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__47486\,
            I => \N__47432\
        );

    \I__10790\ : InMux
    port map (
            O => \N__47485\,
            I => \N__47429\
        );

    \I__10789\ : InMux
    port map (
            O => \N__47484\,
            I => \N__47426\
        );

    \I__10788\ : InMux
    port map (
            O => \N__47483\,
            I => \N__47423\
        );

    \I__10787\ : InMux
    port map (
            O => \N__47482\,
            I => \N__47420\
        );

    \I__10786\ : InMux
    port map (
            O => \N__47481\,
            I => \N__47417\
        );

    \I__10785\ : InMux
    port map (
            O => \N__47480\,
            I => \N__47414\
        );

    \I__10784\ : LocalMux
    port map (
            O => \N__47477\,
            I => \N__47410\
        );

    \I__10783\ : Span4Mux_v
    port map (
            O => \N__47474\,
            I => \N__47399\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__47471\,
            I => \N__47399\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__47468\,
            I => \N__47399\
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__47465\,
            I => \N__47399\
        );

    \I__10779\ : LocalMux
    port map (
            O => \N__47462\,
            I => \N__47399\
        );

    \I__10778\ : InMux
    port map (
            O => \N__47461\,
            I => \N__47396\
        );

    \I__10777\ : InMux
    port map (
            O => \N__47460\,
            I => \N__47390\
        );

    \I__10776\ : InMux
    port map (
            O => \N__47459\,
            I => \N__47387\
        );

    \I__10775\ : InMux
    port map (
            O => \N__47458\,
            I => \N__47384\
        );

    \I__10774\ : InMux
    port map (
            O => \N__47457\,
            I => \N__47381\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__47454\,
            I => \N__47374\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__47451\,
            I => \N__47374\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__47448\,
            I => \N__47371\
        );

    \I__10770\ : InMux
    port map (
            O => \N__47447\,
            I => \N__47368\
        );

    \I__10769\ : InMux
    port map (
            O => \N__47446\,
            I => \N__47365\
        );

    \I__10768\ : Span4Mux_v
    port map (
            O => \N__47443\,
            I => \N__47358\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__47440\,
            I => \N__47358\
        );

    \I__10766\ : InMux
    port map (
            O => \N__47439\,
            I => \N__47355\
        );

    \I__10765\ : InMux
    port map (
            O => \N__47438\,
            I => \N__47352\
        );

    \I__10764\ : InMux
    port map (
            O => \N__47437\,
            I => \N__47349\
        );

    \I__10763\ : Span4Mux_v
    port map (
            O => \N__47432\,
            I => \N__47330\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__47429\,
            I => \N__47330\
        );

    \I__10761\ : LocalMux
    port map (
            O => \N__47426\,
            I => \N__47330\
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__47423\,
            I => \N__47330\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__47420\,
            I => \N__47330\
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__47417\,
            I => \N__47330\
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__47414\,
            I => \N__47325\
        );

    \I__10756\ : InMux
    port map (
            O => \N__47413\,
            I => \N__47322\
        );

    \I__10755\ : Span4Mux_h
    port map (
            O => \N__47410\,
            I => \N__47315\
        );

    \I__10754\ : Span4Mux_v
    port map (
            O => \N__47399\,
            I => \N__47315\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__47396\,
            I => \N__47315\
        );

    \I__10752\ : InMux
    port map (
            O => \N__47395\,
            I => \N__47312\
        );

    \I__10751\ : InMux
    port map (
            O => \N__47394\,
            I => \N__47309\
        );

    \I__10750\ : InMux
    port map (
            O => \N__47393\,
            I => \N__47306\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__47390\,
            I => \N__47301\
        );

    \I__10748\ : LocalMux
    port map (
            O => \N__47387\,
            I => \N__47301\
        );

    \I__10747\ : LocalMux
    port map (
            O => \N__47384\,
            I => \N__47298\
        );

    \I__10746\ : LocalMux
    port map (
            O => \N__47381\,
            I => \N__47295\
        );

    \I__10745\ : InMux
    port map (
            O => \N__47380\,
            I => \N__47292\
        );

    \I__10744\ : InMux
    port map (
            O => \N__47379\,
            I => \N__47289\
        );

    \I__10743\ : Span4Mux_h
    port map (
            O => \N__47374\,
            I => \N__47282\
        );

    \I__10742\ : Span4Mux_v
    port map (
            O => \N__47371\,
            I => \N__47282\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__47368\,
            I => \N__47282\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__47365\,
            I => \N__47279\
        );

    \I__10739\ : InMux
    port map (
            O => \N__47364\,
            I => \N__47276\
        );

    \I__10738\ : InMux
    port map (
            O => \N__47363\,
            I => \N__47272\
        );

    \I__10737\ : Span4Mux_v
    port map (
            O => \N__47358\,
            I => \N__47267\
        );

    \I__10736\ : LocalMux
    port map (
            O => \N__47355\,
            I => \N__47267\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__47352\,
            I => \N__47264\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__47349\,
            I => \N__47261\
        );

    \I__10733\ : InMux
    port map (
            O => \N__47348\,
            I => \N__47258\
        );

    \I__10732\ : InMux
    port map (
            O => \N__47347\,
            I => \N__47255\
        );

    \I__10731\ : InMux
    port map (
            O => \N__47346\,
            I => \N__47252\
        );

    \I__10730\ : InMux
    port map (
            O => \N__47345\,
            I => \N__47248\
        );

    \I__10729\ : InMux
    port map (
            O => \N__47344\,
            I => \N__47241\
        );

    \I__10728\ : InMux
    port map (
            O => \N__47343\,
            I => \N__47238\
        );

    \I__10727\ : Span4Mux_v
    port map (
            O => \N__47330\,
            I => \N__47235\
        );

    \I__10726\ : InMux
    port map (
            O => \N__47329\,
            I => \N__47232\
        );

    \I__10725\ : InMux
    port map (
            O => \N__47328\,
            I => \N__47229\
        );

    \I__10724\ : Span4Mux_v
    port map (
            O => \N__47325\,
            I => \N__47224\
        );

    \I__10723\ : LocalMux
    port map (
            O => \N__47322\,
            I => \N__47224\
        );

    \I__10722\ : Span4Mux_v
    port map (
            O => \N__47315\,
            I => \N__47215\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__47312\,
            I => \N__47215\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__47309\,
            I => \N__47215\
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__47306\,
            I => \N__47215\
        );

    \I__10718\ : Span4Mux_v
    port map (
            O => \N__47301\,
            I => \N__47210\
        );

    \I__10717\ : Span4Mux_v
    port map (
            O => \N__47298\,
            I => \N__47210\
        );

    \I__10716\ : Span4Mux_v
    port map (
            O => \N__47295\,
            I => \N__47203\
        );

    \I__10715\ : LocalMux
    port map (
            O => \N__47292\,
            I => \N__47203\
        );

    \I__10714\ : LocalMux
    port map (
            O => \N__47289\,
            I => \N__47203\
        );

    \I__10713\ : Span4Mux_v
    port map (
            O => \N__47282\,
            I => \N__47195\
        );

    \I__10712\ : Span4Mux_h
    port map (
            O => \N__47279\,
            I => \N__47195\
        );

    \I__10711\ : LocalMux
    port map (
            O => \N__47276\,
            I => \N__47195\
        );

    \I__10710\ : InMux
    port map (
            O => \N__47275\,
            I => \N__47192\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__47272\,
            I => \N__47189\
        );

    \I__10708\ : Span4Mux_v
    port map (
            O => \N__47267\,
            I => \N__47178\
        );

    \I__10707\ : Span4Mux_v
    port map (
            O => \N__47264\,
            I => \N__47178\
        );

    \I__10706\ : Span4Mux_h
    port map (
            O => \N__47261\,
            I => \N__47178\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__47258\,
            I => \N__47178\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__47255\,
            I => \N__47178\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__47252\,
            I => \N__47175\
        );

    \I__10702\ : InMux
    port map (
            O => \N__47251\,
            I => \N__47171\
        );

    \I__10701\ : LocalMux
    port map (
            O => \N__47248\,
            I => \N__47166\
        );

    \I__10700\ : InMux
    port map (
            O => \N__47247\,
            I => \N__47163\
        );

    \I__10699\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47160\
        );

    \I__10698\ : InMux
    port map (
            O => \N__47245\,
            I => \N__47157\
        );

    \I__10697\ : InMux
    port map (
            O => \N__47244\,
            I => \N__47154\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__47241\,
            I => \N__47149\
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__47238\,
            I => \N__47149\
        );

    \I__10694\ : Sp12to4
    port map (
            O => \N__47235\,
            I => \N__47144\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__47232\,
            I => \N__47144\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__47229\,
            I => \N__47141\
        );

    \I__10691\ : Span4Mux_v
    port map (
            O => \N__47224\,
            I => \N__47138\
        );

    \I__10690\ : Span4Mux_v
    port map (
            O => \N__47215\,
            I => \N__47135\
        );

    \I__10689\ : Span4Mux_h
    port map (
            O => \N__47210\,
            I => \N__47130\
        );

    \I__10688\ : Span4Mux_v
    port map (
            O => \N__47203\,
            I => \N__47130\
        );

    \I__10687\ : InMux
    port map (
            O => \N__47202\,
            I => \N__47127\
        );

    \I__10686\ : Span4Mux_h
    port map (
            O => \N__47195\,
            I => \N__47122\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__47192\,
            I => \N__47122\
        );

    \I__10684\ : Span4Mux_v
    port map (
            O => \N__47189\,
            I => \N__47115\
        );

    \I__10683\ : Span4Mux_h
    port map (
            O => \N__47178\,
            I => \N__47110\
        );

    \I__10682\ : Span4Mux_v
    port map (
            O => \N__47175\,
            I => \N__47110\
        );

    \I__10681\ : InMux
    port map (
            O => \N__47174\,
            I => \N__47107\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__47171\,
            I => \N__47104\
        );

    \I__10679\ : InMux
    port map (
            O => \N__47170\,
            I => \N__47101\
        );

    \I__10678\ : InMux
    port map (
            O => \N__47169\,
            I => \N__47098\
        );

    \I__10677\ : Span4Mux_h
    port map (
            O => \N__47166\,
            I => \N__47087\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__47163\,
            I => \N__47087\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__47160\,
            I => \N__47087\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__47157\,
            I => \N__47087\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__47154\,
            I => \N__47087\
        );

    \I__10672\ : Span12Mux_v
    port map (
            O => \N__47149\,
            I => \N__47080\
        );

    \I__10671\ : Span12Mux_h
    port map (
            O => \N__47144\,
            I => \N__47080\
        );

    \I__10670\ : Span12Mux_s10_v
    port map (
            O => \N__47141\,
            I => \N__47080\
        );

    \I__10669\ : Span4Mux_v
    port map (
            O => \N__47138\,
            I => \N__47075\
        );

    \I__10668\ : Span4Mux_v
    port map (
            O => \N__47135\,
            I => \N__47075\
        );

    \I__10667\ : Span4Mux_v
    port map (
            O => \N__47130\,
            I => \N__47070\
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__47127\,
            I => \N__47070\
        );

    \I__10665\ : Span4Mux_h
    port map (
            O => \N__47122\,
            I => \N__47067\
        );

    \I__10664\ : InMux
    port map (
            O => \N__47121\,
            I => \N__47064\
        );

    \I__10663\ : InMux
    port map (
            O => \N__47120\,
            I => \N__47061\
        );

    \I__10662\ : InMux
    port map (
            O => \N__47119\,
            I => \N__47058\
        );

    \I__10661\ : InMux
    port map (
            O => \N__47118\,
            I => \N__47055\
        );

    \I__10660\ : Span4Mux_v
    port map (
            O => \N__47115\,
            I => \N__47048\
        );

    \I__10659\ : Span4Mux_h
    port map (
            O => \N__47110\,
            I => \N__47048\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__47107\,
            I => \N__47048\
        );

    \I__10657\ : Span4Mux_v
    port map (
            O => \N__47104\,
            I => \N__47039\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__47101\,
            I => \N__47039\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__47098\,
            I => \N__47039\
        );

    \I__10654\ : Span4Mux_v
    port map (
            O => \N__47087\,
            I => \N__47039\
        );

    \I__10653\ : Odrv12
    port map (
            O => \N__47080\,
            I => spi_data_mosi_2
        );

    \I__10652\ : Odrv4
    port map (
            O => \N__47075\,
            I => spi_data_mosi_2
        );

    \I__10651\ : Odrv4
    port map (
            O => \N__47070\,
            I => spi_data_mosi_2
        );

    \I__10650\ : Odrv4
    port map (
            O => \N__47067\,
            I => spi_data_mosi_2
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__47064\,
            I => spi_data_mosi_2
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__47061\,
            I => spi_data_mosi_2
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__47058\,
            I => spi_data_mosi_2
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__47055\,
            I => spi_data_mosi_2
        );

    \I__10645\ : Odrv4
    port map (
            O => \N__47048\,
            I => spi_data_mosi_2
        );

    \I__10644\ : Odrv4
    port map (
            O => \N__47039\,
            I => spi_data_mosi_2
        );

    \I__10643\ : InMux
    port map (
            O => \N__47018\,
            I => \N__47014\
        );

    \I__10642\ : InMux
    port map (
            O => \N__47017\,
            I => \N__47011\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__47014\,
            I => \sCounterADCZ0Z_2\
        );

    \I__10640\ : LocalMux
    port map (
            O => \N__47011\,
            I => \sCounterADCZ0Z_2\
        );

    \I__10639\ : InMux
    port map (
            O => \N__47006\,
            I => \N__47003\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__47003\,
            I => \sEEADC_freqZ0Z_2\
        );

    \I__10637\ : InMux
    port map (
            O => \N__47000\,
            I => \N__46996\
        );

    \I__10636\ : InMux
    port map (
            O => \N__46999\,
            I => \N__46993\
        );

    \I__10635\ : LocalMux
    port map (
            O => \N__46996\,
            I => \sCounterADCZ0Z_3\
        );

    \I__10634\ : LocalMux
    port map (
            O => \N__46993\,
            I => \sCounterADCZ0Z_3\
        );

    \I__10633\ : InMux
    port map (
            O => \N__46988\,
            I => \N__46985\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__46985\,
            I => \N__46982\
        );

    \I__10631\ : Span12Mux_v
    port map (
            O => \N__46982\,
            I => \N__46979\
        );

    \I__10630\ : Span12Mux_h
    port map (
            O => \N__46979\,
            I => \N__46976\
        );

    \I__10629\ : Odrv12
    port map (
            O => \N__46976\,
            I => \un11_sacqtime_NE_3\
        );

    \I__10628\ : CascadeMux
    port map (
            O => \N__46973\,
            I => \un11_sacqtime_NE_0_0_cascade_\
        );

    \I__10627\ : CascadeMux
    port map (
            O => \N__46970\,
            I => \N__46967\
        );

    \I__10626\ : InMux
    port map (
            O => \N__46967\,
            I => \N__46964\
        );

    \I__10625\ : LocalMux
    port map (
            O => \N__46964\,
            I => \N__46953\
        );

    \I__10624\ : InMux
    port map (
            O => \N__46963\,
            I => \N__46944\
        );

    \I__10623\ : InMux
    port map (
            O => \N__46962\,
            I => \N__46944\
        );

    \I__10622\ : InMux
    port map (
            O => \N__46961\,
            I => \N__46944\
        );

    \I__10621\ : InMux
    port map (
            O => \N__46960\,
            I => \N__46944\
        );

    \I__10620\ : InMux
    port map (
            O => \N__46959\,
            I => \N__46935\
        );

    \I__10619\ : InMux
    port map (
            O => \N__46958\,
            I => \N__46935\
        );

    \I__10618\ : InMux
    port map (
            O => \N__46957\,
            I => \N__46935\
        );

    \I__10617\ : InMux
    port map (
            O => \N__46956\,
            I => \N__46935\
        );

    \I__10616\ : Span4Mux_h
    port map (
            O => \N__46953\,
            I => \N__46932\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__46944\,
            I => \un11_sacqtime_NE_0\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__46935\,
            I => \un11_sacqtime_NE_0\
        );

    \I__10613\ : Odrv4
    port map (
            O => \N__46932\,
            I => \un11_sacqtime_NE_0\
        );

    \I__10612\ : InMux
    port map (
            O => \N__46925\,
            I => \N__46916\
        );

    \I__10611\ : InMux
    port map (
            O => \N__46924\,
            I => \N__46910\
        );

    \I__10610\ : InMux
    port map (
            O => \N__46923\,
            I => \N__46902\
        );

    \I__10609\ : InMux
    port map (
            O => \N__46922\,
            I => \N__46898\
        );

    \I__10608\ : InMux
    port map (
            O => \N__46921\,
            I => \N__46895\
        );

    \I__10607\ : InMux
    port map (
            O => \N__46920\,
            I => \N__46892\
        );

    \I__10606\ : InMux
    port map (
            O => \N__46919\,
            I => \N__46888\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__46916\,
            I => \N__46885\
        );

    \I__10604\ : InMux
    port map (
            O => \N__46915\,
            I => \N__46882\
        );

    \I__10603\ : InMux
    port map (
            O => \N__46914\,
            I => \N__46879\
        );

    \I__10602\ : InMux
    port map (
            O => \N__46913\,
            I => \N__46876\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__46910\,
            I => \N__46873\
        );

    \I__10600\ : InMux
    port map (
            O => \N__46909\,
            I => \N__46870\
        );

    \I__10599\ : InMux
    port map (
            O => \N__46908\,
            I => \N__46867\
        );

    \I__10598\ : InMux
    port map (
            O => \N__46907\,
            I => \N__46863\
        );

    \I__10597\ : InMux
    port map (
            O => \N__46906\,
            I => \N__46860\
        );

    \I__10596\ : InMux
    port map (
            O => \N__46905\,
            I => \N__46848\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__46902\,
            I => \N__46844\
        );

    \I__10594\ : InMux
    port map (
            O => \N__46901\,
            I => \N__46841\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__46898\,
            I => \N__46833\
        );

    \I__10592\ : LocalMux
    port map (
            O => \N__46895\,
            I => \N__46833\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__46892\,
            I => \N__46833\
        );

    \I__10590\ : InMux
    port map (
            O => \N__46891\,
            I => \N__46830\
        );

    \I__10589\ : LocalMux
    port map (
            O => \N__46888\,
            I => \N__46826\
        );

    \I__10588\ : Span4Mux_v
    port map (
            O => \N__46885\,
            I => \N__46817\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__46882\,
            I => \N__46817\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__46879\,
            I => \N__46817\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__46876\,
            I => \N__46817\
        );

    \I__10584\ : Span4Mux_h
    port map (
            O => \N__46873\,
            I => \N__46810\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__46870\,
            I => \N__46810\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__46867\,
            I => \N__46810\
        );

    \I__10581\ : InMux
    port map (
            O => \N__46866\,
            I => \N__46807\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__46863\,
            I => \N__46804\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__46860\,
            I => \N__46801\
        );

    \I__10578\ : InMux
    port map (
            O => \N__46859\,
            I => \N__46798\
        );

    \I__10577\ : InMux
    port map (
            O => \N__46858\,
            I => \N__46795\
        );

    \I__10576\ : InMux
    port map (
            O => \N__46857\,
            I => \N__46790\
        );

    \I__10575\ : InMux
    port map (
            O => \N__46856\,
            I => \N__46786\
        );

    \I__10574\ : InMux
    port map (
            O => \N__46855\,
            I => \N__46783\
        );

    \I__10573\ : InMux
    port map (
            O => \N__46854\,
            I => \N__46780\
        );

    \I__10572\ : InMux
    port map (
            O => \N__46853\,
            I => \N__46776\
        );

    \I__10571\ : InMux
    port map (
            O => \N__46852\,
            I => \N__46771\
        );

    \I__10570\ : InMux
    port map (
            O => \N__46851\,
            I => \N__46766\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__46848\,
            I => \N__46759\
        );

    \I__10568\ : InMux
    port map (
            O => \N__46847\,
            I => \N__46756\
        );

    \I__10567\ : Span4Mux_v
    port map (
            O => \N__46844\,
            I => \N__46753\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__46841\,
            I => \N__46747\
        );

    \I__10565\ : InMux
    port map (
            O => \N__46840\,
            I => \N__46743\
        );

    \I__10564\ : Span4Mux_h
    port map (
            O => \N__46833\,
            I => \N__46738\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__46830\,
            I => \N__46738\
        );

    \I__10562\ : InMux
    port map (
            O => \N__46829\,
            I => \N__46735\
        );

    \I__10561\ : Span4Mux_h
    port map (
            O => \N__46826\,
            I => \N__46726\
        );

    \I__10560\ : Span4Mux_h
    port map (
            O => \N__46817\,
            I => \N__46726\
        );

    \I__10559\ : Span4Mux_v
    port map (
            O => \N__46810\,
            I => \N__46726\
        );

    \I__10558\ : LocalMux
    port map (
            O => \N__46807\,
            I => \N__46726\
        );

    \I__10557\ : Span4Mux_v
    port map (
            O => \N__46804\,
            I => \N__46719\
        );

    \I__10556\ : Span4Mux_h
    port map (
            O => \N__46801\,
            I => \N__46719\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__46798\,
            I => \N__46719\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__46795\,
            I => \N__46716\
        );

    \I__10553\ : InMux
    port map (
            O => \N__46794\,
            I => \N__46713\
        );

    \I__10552\ : InMux
    port map (
            O => \N__46793\,
            I => \N__46710\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__46790\,
            I => \N__46704\
        );

    \I__10550\ : InMux
    port map (
            O => \N__46789\,
            I => \N__46701\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__46786\,
            I => \N__46696\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__46783\,
            I => \N__46696\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__46780\,
            I => \N__46693\
        );

    \I__10546\ : InMux
    port map (
            O => \N__46779\,
            I => \N__46690\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__46776\,
            I => \N__46686\
        );

    \I__10544\ : InMux
    port map (
            O => \N__46775\,
            I => \N__46683\
        );

    \I__10543\ : InMux
    port map (
            O => \N__46774\,
            I => \N__46680\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__46771\,
            I => \N__46677\
        );

    \I__10541\ : InMux
    port map (
            O => \N__46770\,
            I => \N__46674\
        );

    \I__10540\ : InMux
    port map (
            O => \N__46769\,
            I => \N__46671\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__46766\,
            I => \N__46668\
        );

    \I__10538\ : InMux
    port map (
            O => \N__46765\,
            I => \N__46665\
        );

    \I__10537\ : InMux
    port map (
            O => \N__46764\,
            I => \N__46662\
        );

    \I__10536\ : InMux
    port map (
            O => \N__46763\,
            I => \N__46659\
        );

    \I__10535\ : InMux
    port map (
            O => \N__46762\,
            I => \N__46656\
        );

    \I__10534\ : Span4Mux_h
    port map (
            O => \N__46759\,
            I => \N__46651\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__46756\,
            I => \N__46651\
        );

    \I__10532\ : Span4Mux_v
    port map (
            O => \N__46753\,
            I => \N__46647\
        );

    \I__10531\ : InMux
    port map (
            O => \N__46752\,
            I => \N__46644\
        );

    \I__10530\ : InMux
    port map (
            O => \N__46751\,
            I => \N__46641\
        );

    \I__10529\ : InMux
    port map (
            O => \N__46750\,
            I => \N__46638\
        );

    \I__10528\ : Span4Mux_v
    port map (
            O => \N__46747\,
            I => \N__46635\
        );

    \I__10527\ : InMux
    port map (
            O => \N__46746\,
            I => \N__46632\
        );

    \I__10526\ : LocalMux
    port map (
            O => \N__46743\,
            I => \N__46629\
        );

    \I__10525\ : Span4Mux_h
    port map (
            O => \N__46738\,
            I => \N__46624\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__46735\,
            I => \N__46624\
        );

    \I__10523\ : Span4Mux_v
    port map (
            O => \N__46726\,
            I => \N__46621\
        );

    \I__10522\ : Span4Mux_v
    port map (
            O => \N__46719\,
            I => \N__46614\
        );

    \I__10521\ : Span4Mux_h
    port map (
            O => \N__46716\,
            I => \N__46614\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__46713\,
            I => \N__46614\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__46710\,
            I => \N__46611\
        );

    \I__10518\ : InMux
    port map (
            O => \N__46709\,
            I => \N__46608\
        );

    \I__10517\ : InMux
    port map (
            O => \N__46708\,
            I => \N__46605\
        );

    \I__10516\ : InMux
    port map (
            O => \N__46707\,
            I => \N__46600\
        );

    \I__10515\ : Span4Mux_v
    port map (
            O => \N__46704\,
            I => \N__46593\
        );

    \I__10514\ : LocalMux
    port map (
            O => \N__46701\,
            I => \N__46593\
        );

    \I__10513\ : Span4Mux_h
    port map (
            O => \N__46696\,
            I => \N__46586\
        );

    \I__10512\ : Span4Mux_v
    port map (
            O => \N__46693\,
            I => \N__46586\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__46690\,
            I => \N__46586\
        );

    \I__10510\ : InMux
    port map (
            O => \N__46689\,
            I => \N__46583\
        );

    \I__10509\ : Span4Mux_h
    port map (
            O => \N__46686\,
            I => \N__46572\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__46683\,
            I => \N__46572\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__46680\,
            I => \N__46572\
        );

    \I__10506\ : Span4Mux_h
    port map (
            O => \N__46677\,
            I => \N__46572\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__46674\,
            I => \N__46572\
        );

    \I__10504\ : LocalMux
    port map (
            O => \N__46671\,
            I => \N__46569\
        );

    \I__10503\ : Span4Mux_h
    port map (
            O => \N__46668\,
            I => \N__46566\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__46665\,
            I => \N__46557\
        );

    \I__10501\ : LocalMux
    port map (
            O => \N__46662\,
            I => \N__46557\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__46659\,
            I => \N__46557\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__46656\,
            I => \N__46557\
        );

    \I__10498\ : Span4Mux_h
    port map (
            O => \N__46651\,
            I => \N__46554\
        );

    \I__10497\ : InMux
    port map (
            O => \N__46650\,
            I => \N__46551\
        );

    \I__10496\ : Sp12to4
    port map (
            O => \N__46647\,
            I => \N__46538\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__46644\,
            I => \N__46538\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__46641\,
            I => \N__46538\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__46638\,
            I => \N__46538\
        );

    \I__10492\ : Sp12to4
    port map (
            O => \N__46635\,
            I => \N__46538\
        );

    \I__10491\ : LocalMux
    port map (
            O => \N__46632\,
            I => \N__46538\
        );

    \I__10490\ : Span4Mux_h
    port map (
            O => \N__46629\,
            I => \N__46533\
        );

    \I__10489\ : Span4Mux_h
    port map (
            O => \N__46624\,
            I => \N__46533\
        );

    \I__10488\ : Span4Mux_v
    port map (
            O => \N__46621\,
            I => \N__46522\
        );

    \I__10487\ : Span4Mux_h
    port map (
            O => \N__46614\,
            I => \N__46522\
        );

    \I__10486\ : Span4Mux_v
    port map (
            O => \N__46611\,
            I => \N__46522\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__46608\,
            I => \N__46522\
        );

    \I__10484\ : LocalMux
    port map (
            O => \N__46605\,
            I => \N__46522\
        );

    \I__10483\ : InMux
    port map (
            O => \N__46604\,
            I => \N__46515\
        );

    \I__10482\ : InMux
    port map (
            O => \N__46603\,
            I => \N__46512\
        );

    \I__10481\ : LocalMux
    port map (
            O => \N__46600\,
            I => \N__46509\
        );

    \I__10480\ : InMux
    port map (
            O => \N__46599\,
            I => \N__46506\
        );

    \I__10479\ : InMux
    port map (
            O => \N__46598\,
            I => \N__46503\
        );

    \I__10478\ : Span4Mux_h
    port map (
            O => \N__46593\,
            I => \N__46494\
        );

    \I__10477\ : Span4Mux_v
    port map (
            O => \N__46586\,
            I => \N__46494\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__46583\,
            I => \N__46494\
        );

    \I__10475\ : Span4Mux_v
    port map (
            O => \N__46572\,
            I => \N__46494\
        );

    \I__10474\ : Span4Mux_h
    port map (
            O => \N__46569\,
            I => \N__46491\
        );

    \I__10473\ : Sp12to4
    port map (
            O => \N__46566\,
            I => \N__46478\
        );

    \I__10472\ : Span12Mux_h
    port map (
            O => \N__46557\,
            I => \N__46478\
        );

    \I__10471\ : Sp12to4
    port map (
            O => \N__46554\,
            I => \N__46478\
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__46551\,
            I => \N__46478\
        );

    \I__10469\ : Span12Mux_h
    port map (
            O => \N__46538\,
            I => \N__46478\
        );

    \I__10468\ : Sp12to4
    port map (
            O => \N__46533\,
            I => \N__46478\
        );

    \I__10467\ : Span4Mux_h
    port map (
            O => \N__46522\,
            I => \N__46475\
        );

    \I__10466\ : InMux
    port map (
            O => \N__46521\,
            I => \N__46472\
        );

    \I__10465\ : InMux
    port map (
            O => \N__46520\,
            I => \N__46469\
        );

    \I__10464\ : InMux
    port map (
            O => \N__46519\,
            I => \N__46466\
        );

    \I__10463\ : InMux
    port map (
            O => \N__46518\,
            I => \N__46463\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__46515\,
            I => \N__46458\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__46512\,
            I => \N__46458\
        );

    \I__10460\ : Span4Mux_v
    port map (
            O => \N__46509\,
            I => \N__46449\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__46506\,
            I => \N__46449\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__46503\,
            I => \N__46449\
        );

    \I__10457\ : Span4Mux_h
    port map (
            O => \N__46494\,
            I => \N__46449\
        );

    \I__10456\ : Odrv4
    port map (
            O => \N__46491\,
            I => spi_data_mosi_3
        );

    \I__10455\ : Odrv12
    port map (
            O => \N__46478\,
            I => spi_data_mosi_3
        );

    \I__10454\ : Odrv4
    port map (
            O => \N__46475\,
            I => spi_data_mosi_3
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__46472\,
            I => spi_data_mosi_3
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__46469\,
            I => spi_data_mosi_3
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__46466\,
            I => spi_data_mosi_3
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__46463\,
            I => spi_data_mosi_3
        );

    \I__10449\ : Odrv4
    port map (
            O => \N__46458\,
            I => spi_data_mosi_3
        );

    \I__10448\ : Odrv4
    port map (
            O => \N__46449\,
            I => spi_data_mosi_3
        );

    \I__10447\ : CascadeMux
    port map (
            O => \N__46430\,
            I => \N__46427\
        );

    \I__10446\ : InMux
    port map (
            O => \N__46427\,
            I => \N__46424\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__46424\,
            I => \sEEADC_freqZ0Z_3\
        );

    \I__10444\ : InMux
    port map (
            O => \N__46421\,
            I => \N__46417\
        );

    \I__10443\ : InMux
    port map (
            O => \N__46420\,
            I => \N__46414\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__46417\,
            I => \sCounterADCZ0Z_1\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__46414\,
            I => \sCounterADCZ0Z_1\
        );

    \I__10440\ : InMux
    port map (
            O => \N__46409\,
            I => \N__46405\
        );

    \I__10439\ : InMux
    port map (
            O => \N__46408\,
            I => \N__46402\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__46405\,
            I => \sCounterADCZ0Z_0\
        );

    \I__10437\ : LocalMux
    port map (
            O => \N__46402\,
            I => \sCounterADCZ0Z_0\
        );

    \I__10436\ : InMux
    port map (
            O => \N__46397\,
            I => \N__46394\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__46394\,
            I => \un11_sacqtime_NE_1\
        );

    \I__10434\ : InMux
    port map (
            O => \N__46391\,
            I => \N__46376\
        );

    \I__10433\ : InMux
    port map (
            O => \N__46390\,
            I => \N__46371\
        );

    \I__10432\ : InMux
    port map (
            O => \N__46389\,
            I => \N__46368\
        );

    \I__10431\ : InMux
    port map (
            O => \N__46388\,
            I => \N__46365\
        );

    \I__10430\ : InMux
    port map (
            O => \N__46387\,
            I => \N__46362\
        );

    \I__10429\ : InMux
    port map (
            O => \N__46386\,
            I => \N__46359\
        );

    \I__10428\ : InMux
    port map (
            O => \N__46385\,
            I => \N__46356\
        );

    \I__10427\ : InMux
    port map (
            O => \N__46384\,
            I => \N__46353\
        );

    \I__10426\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46349\
        );

    \I__10425\ : InMux
    port map (
            O => \N__46382\,
            I => \N__46346\
        );

    \I__10424\ : InMux
    port map (
            O => \N__46381\,
            I => \N__46339\
        );

    \I__10423\ : InMux
    port map (
            O => \N__46380\,
            I => \N__46335\
        );

    \I__10422\ : InMux
    port map (
            O => \N__46379\,
            I => \N__46332\
        );

    \I__10421\ : LocalMux
    port map (
            O => \N__46376\,
            I => \N__46328\
        );

    \I__10420\ : InMux
    port map (
            O => \N__46375\,
            I => \N__46325\
        );

    \I__10419\ : InMux
    port map (
            O => \N__46374\,
            I => \N__46318\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__46371\,
            I => \N__46309\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__46368\,
            I => \N__46309\
        );

    \I__10416\ : LocalMux
    port map (
            O => \N__46365\,
            I => \N__46300\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__46362\,
            I => \N__46300\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__46359\,
            I => \N__46300\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__46356\,
            I => \N__46300\
        );

    \I__10412\ : LocalMux
    port map (
            O => \N__46353\,
            I => \N__46297\
        );

    \I__10411\ : InMux
    port map (
            O => \N__46352\,
            I => \N__46294\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__46349\,
            I => \N__46288\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__46346\,
            I => \N__46288\
        );

    \I__10408\ : InMux
    port map (
            O => \N__46345\,
            I => \N__46285\
        );

    \I__10407\ : InMux
    port map (
            O => \N__46344\,
            I => \N__46282\
        );

    \I__10406\ : InMux
    port map (
            O => \N__46343\,
            I => \N__46276\
        );

    \I__10405\ : InMux
    port map (
            O => \N__46342\,
            I => \N__46273\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__46339\,
            I => \N__46270\
        );

    \I__10403\ : InMux
    port map (
            O => \N__46338\,
            I => \N__46267\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__46335\,
            I => \N__46262\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__46332\,
            I => \N__46262\
        );

    \I__10400\ : InMux
    port map (
            O => \N__46331\,
            I => \N__46259\
        );

    \I__10399\ : Span4Mux_v
    port map (
            O => \N__46328\,
            I => \N__46254\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__46325\,
            I => \N__46254\
        );

    \I__10397\ : InMux
    port map (
            O => \N__46324\,
            I => \N__46251\
        );

    \I__10396\ : InMux
    port map (
            O => \N__46323\,
            I => \N__46248\
        );

    \I__10395\ : InMux
    port map (
            O => \N__46322\,
            I => \N__46245\
        );

    \I__10394\ : InMux
    port map (
            O => \N__46321\,
            I => \N__46242\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__46318\,
            I => \N__46239\
        );

    \I__10392\ : InMux
    port map (
            O => \N__46317\,
            I => \N__46236\
        );

    \I__10391\ : InMux
    port map (
            O => \N__46316\,
            I => \N__46230\
        );

    \I__10390\ : InMux
    port map (
            O => \N__46315\,
            I => \N__46227\
        );

    \I__10389\ : InMux
    port map (
            O => \N__46314\,
            I => \N__46224\
        );

    \I__10388\ : Span4Mux_h
    port map (
            O => \N__46309\,
            I => \N__46215\
        );

    \I__10387\ : Span4Mux_v
    port map (
            O => \N__46300\,
            I => \N__46215\
        );

    \I__10386\ : Span4Mux_h
    port map (
            O => \N__46297\,
            I => \N__46215\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__46294\,
            I => \N__46215\
        );

    \I__10384\ : InMux
    port map (
            O => \N__46293\,
            I => \N__46212\
        );

    \I__10383\ : Span4Mux_v
    port map (
            O => \N__46288\,
            I => \N__46202\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__46285\,
            I => \N__46202\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__46282\,
            I => \N__46202\
        );

    \I__10380\ : InMux
    port map (
            O => \N__46281\,
            I => \N__46199\
        );

    \I__10379\ : InMux
    port map (
            O => \N__46280\,
            I => \N__46196\
        );

    \I__10378\ : InMux
    port map (
            O => \N__46279\,
            I => \N__46193\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__46276\,
            I => \N__46184\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__46273\,
            I => \N__46184\
        );

    \I__10375\ : Span4Mux_h
    port map (
            O => \N__46270\,
            I => \N__46184\
        );

    \I__10374\ : LocalMux
    port map (
            O => \N__46267\,
            I => \N__46184\
        );

    \I__10373\ : Span4Mux_v
    port map (
            O => \N__46262\,
            I => \N__46179\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__46259\,
            I => \N__46179\
        );

    \I__10371\ : Span4Mux_h
    port map (
            O => \N__46254\,
            I => \N__46174\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__46251\,
            I => \N__46174\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__46248\,
            I => \N__46167\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__46245\,
            I => \N__46167\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__46242\,
            I => \N__46167\
        );

    \I__10366\ : Span4Mux_h
    port map (
            O => \N__46239\,
            I => \N__46162\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__46236\,
            I => \N__46162\
        );

    \I__10364\ : InMux
    port map (
            O => \N__46235\,
            I => \N__46159\
        );

    \I__10363\ : InMux
    port map (
            O => \N__46234\,
            I => \N__46156\
        );

    \I__10362\ : InMux
    port map (
            O => \N__46233\,
            I => \N__46153\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__46230\,
            I => \N__46150\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__46227\,
            I => \N__46136\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__46224\,
            I => \N__46136\
        );

    \I__10358\ : Span4Mux_v
    port map (
            O => \N__46215\,
            I => \N__46131\
        );

    \I__10357\ : LocalMux
    port map (
            O => \N__46212\,
            I => \N__46131\
        );

    \I__10356\ : CascadeMux
    port map (
            O => \N__46211\,
            I => \N__46127\
        );

    \I__10355\ : InMux
    port map (
            O => \N__46210\,
            I => \N__46124\
        );

    \I__10354\ : InMux
    port map (
            O => \N__46209\,
            I => \N__46121\
        );

    \I__10353\ : Span4Mux_h
    port map (
            O => \N__46202\,
            I => \N__46118\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__46199\,
            I => \N__46115\
        );

    \I__10351\ : LocalMux
    port map (
            O => \N__46196\,
            I => \N__46106\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__46193\,
            I => \N__46106\
        );

    \I__10349\ : Span4Mux_h
    port map (
            O => \N__46184\,
            I => \N__46106\
        );

    \I__10348\ : Span4Mux_h
    port map (
            O => \N__46179\,
            I => \N__46106\
        );

    \I__10347\ : Span4Mux_v
    port map (
            O => \N__46174\,
            I => \N__46101\
        );

    \I__10346\ : Span4Mux_v
    port map (
            O => \N__46167\,
            I => \N__46101\
        );

    \I__10345\ : Span4Mux_v
    port map (
            O => \N__46162\,
            I => \N__46098\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__46159\,
            I => \N__46093\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__46156\,
            I => \N__46093\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__46153\,
            I => \N__46090\
        );

    \I__10341\ : Span4Mux_v
    port map (
            O => \N__46150\,
            I => \N__46087\
        );

    \I__10340\ : InMux
    port map (
            O => \N__46149\,
            I => \N__46084\
        );

    \I__10339\ : InMux
    port map (
            O => \N__46148\,
            I => \N__46081\
        );

    \I__10338\ : InMux
    port map (
            O => \N__46147\,
            I => \N__46078\
        );

    \I__10337\ : InMux
    port map (
            O => \N__46146\,
            I => \N__46075\
        );

    \I__10336\ : InMux
    port map (
            O => \N__46145\,
            I => \N__46072\
        );

    \I__10335\ : InMux
    port map (
            O => \N__46144\,
            I => \N__46069\
        );

    \I__10334\ : InMux
    port map (
            O => \N__46143\,
            I => \N__46066\
        );

    \I__10333\ : InMux
    port map (
            O => \N__46142\,
            I => \N__46063\
        );

    \I__10332\ : InMux
    port map (
            O => \N__46141\,
            I => \N__46060\
        );

    \I__10331\ : Span4Mux_v
    port map (
            O => \N__46136\,
            I => \N__46055\
        );

    \I__10330\ : Span4Mux_v
    port map (
            O => \N__46131\,
            I => \N__46055\
        );

    \I__10329\ : InMux
    port map (
            O => \N__46130\,
            I => \N__46047\
        );

    \I__10328\ : InMux
    port map (
            O => \N__46127\,
            I => \N__46044\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__46124\,
            I => \N__46039\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__46121\,
            I => \N__46034\
        );

    \I__10325\ : Span4Mux_h
    port map (
            O => \N__46118\,
            I => \N__46034\
        );

    \I__10324\ : Span4Mux_h
    port map (
            O => \N__46115\,
            I => \N__46029\
        );

    \I__10323\ : Span4Mux_v
    port map (
            O => \N__46106\,
            I => \N__46029\
        );

    \I__10322\ : Span4Mux_h
    port map (
            O => \N__46101\,
            I => \N__46022\
        );

    \I__10321\ : Span4Mux_h
    port map (
            O => \N__46098\,
            I => \N__46022\
        );

    \I__10320\ : Span4Mux_v
    port map (
            O => \N__46093\,
            I => \N__46022\
        );

    \I__10319\ : Span4Mux_v
    port map (
            O => \N__46090\,
            I => \N__46019\
        );

    \I__10318\ : Sp12to4
    port map (
            O => \N__46087\,
            I => \N__46016\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__46084\,
            I => \N__46010\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__46081\,
            I => \N__46010\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__46078\,
            I => \N__46005\
        );

    \I__10314\ : LocalMux
    port map (
            O => \N__46075\,
            I => \N__46005\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__46072\,
            I => \N__46002\
        );

    \I__10312\ : LocalMux
    port map (
            O => \N__46069\,
            I => \N__45999\
        );

    \I__10311\ : LocalMux
    port map (
            O => \N__46066\,
            I => \N__45990\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__46063\,
            I => \N__45990\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__46060\,
            I => \N__45990\
        );

    \I__10308\ : Span4Mux_h
    port map (
            O => \N__46055\,
            I => \N__45990\
        );

    \I__10307\ : InMux
    port map (
            O => \N__46054\,
            I => \N__45987\
        );

    \I__10306\ : InMux
    port map (
            O => \N__46053\,
            I => \N__45980\
        );

    \I__10305\ : InMux
    port map (
            O => \N__46052\,
            I => \N__45980\
        );

    \I__10304\ : InMux
    port map (
            O => \N__46051\,
            I => \N__45980\
        );

    \I__10303\ : InMux
    port map (
            O => \N__46050\,
            I => \N__45974\
        );

    \I__10302\ : LocalMux
    port map (
            O => \N__46047\,
            I => \N__45969\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__46044\,
            I => \N__45969\
        );

    \I__10300\ : InMux
    port map (
            O => \N__46043\,
            I => \N__45966\
        );

    \I__10299\ : InMux
    port map (
            O => \N__46042\,
            I => \N__45963\
        );

    \I__10298\ : Span4Mux_h
    port map (
            O => \N__46039\,
            I => \N__45956\
        );

    \I__10297\ : Span4Mux_h
    port map (
            O => \N__46034\,
            I => \N__45956\
        );

    \I__10296\ : Span4Mux_v
    port map (
            O => \N__46029\,
            I => \N__45956\
        );

    \I__10295\ : Sp12to4
    port map (
            O => \N__46022\,
            I => \N__45953\
        );

    \I__10294\ : Sp12to4
    port map (
            O => \N__46019\,
            I => \N__45948\
        );

    \I__10293\ : Span12Mux_v
    port map (
            O => \N__46016\,
            I => \N__45948\
        );

    \I__10292\ : InMux
    port map (
            O => \N__46015\,
            I => \N__45945\
        );

    \I__10291\ : Span4Mux_v
    port map (
            O => \N__46010\,
            I => \N__45942\
        );

    \I__10290\ : Span4Mux_v
    port map (
            O => \N__46005\,
            I => \N__45935\
        );

    \I__10289\ : Span4Mux_h
    port map (
            O => \N__46002\,
            I => \N__45935\
        );

    \I__10288\ : Span4Mux_v
    port map (
            O => \N__45999\,
            I => \N__45935\
        );

    \I__10287\ : Span4Mux_v
    port map (
            O => \N__45990\,
            I => \N__45932\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__45987\,
            I => \N__45927\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__45980\,
            I => \N__45927\
        );

    \I__10284\ : InMux
    port map (
            O => \N__45979\,
            I => \N__45924\
        );

    \I__10283\ : InMux
    port map (
            O => \N__45978\,
            I => \N__45921\
        );

    \I__10282\ : InMux
    port map (
            O => \N__45977\,
            I => \N__45918\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__45974\,
            I => \N__45911\
        );

    \I__10280\ : Span4Mux_v
    port map (
            O => \N__45969\,
            I => \N__45911\
        );

    \I__10279\ : LocalMux
    port map (
            O => \N__45966\,
            I => \N__45911\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__45963\,
            I => \N__45908\
        );

    \I__10277\ : Span4Mux_v
    port map (
            O => \N__45956\,
            I => \N__45905\
        );

    \I__10276\ : Span12Mux_h
    port map (
            O => \N__45953\,
            I => \N__45900\
        );

    \I__10275\ : Span12Mux_h
    port map (
            O => \N__45948\,
            I => \N__45900\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__45945\,
            I => \N__45889\
        );

    \I__10273\ : Span4Mux_v
    port map (
            O => \N__45942\,
            I => \N__45889\
        );

    \I__10272\ : Span4Mux_h
    port map (
            O => \N__45935\,
            I => \N__45889\
        );

    \I__10271\ : Span4Mux_h
    port map (
            O => \N__45932\,
            I => \N__45889\
        );

    \I__10270\ : Span4Mux_h
    port map (
            O => \N__45927\,
            I => \N__45889\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__45924\,
            I => spi_data_mosi_0
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__45921\,
            I => spi_data_mosi_0
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__45918\,
            I => spi_data_mosi_0
        );

    \I__10266\ : Odrv4
    port map (
            O => \N__45911\,
            I => spi_data_mosi_0
        );

    \I__10265\ : Odrv4
    port map (
            O => \N__45908\,
            I => spi_data_mosi_0
        );

    \I__10264\ : Odrv4
    port map (
            O => \N__45905\,
            I => spi_data_mosi_0
        );

    \I__10263\ : Odrv12
    port map (
            O => \N__45900\,
            I => spi_data_mosi_0
        );

    \I__10262\ : Odrv4
    port map (
            O => \N__45889\,
            I => spi_data_mosi_0
        );

    \I__10261\ : InMux
    port map (
            O => \N__45872\,
            I => \N__45869\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__45869\,
            I => \sEEADC_freqZ0Z_0\
        );

    \I__10259\ : CascadeMux
    port map (
            O => \N__45866\,
            I => \N__45863\
        );

    \I__10258\ : InMux
    port map (
            O => \N__45863\,
            I => \N__45860\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__45860\,
            I => \sEEADC_freqZ0Z_1\
        );

    \I__10256\ : InMux
    port map (
            O => \N__45857\,
            I => \N__45853\
        );

    \I__10255\ : InMux
    port map (
            O => \N__45856\,
            I => \N__45850\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__45853\,
            I => \sCounterADCZ0Z_7\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__45850\,
            I => \sCounterADCZ0Z_7\
        );

    \I__10252\ : CascadeMux
    port map (
            O => \N__45845\,
            I => \N__45841\
        );

    \I__10251\ : InMux
    port map (
            O => \N__45844\,
            I => \N__45838\
        );

    \I__10250\ : InMux
    port map (
            O => \N__45841\,
            I => \N__45835\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__45838\,
            I => \sCounterADCZ0Z_6\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__45835\,
            I => \sCounterADCZ0Z_6\
        );

    \I__10247\ : InMux
    port map (
            O => \N__45830\,
            I => \N__45827\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__45827\,
            I => \un11_sacqtime_NE_2\
        );

    \I__10245\ : InMux
    port map (
            O => \N__45824\,
            I => \N__45821\
        );

    \I__10244\ : LocalMux
    port map (
            O => \N__45821\,
            I => \N__45818\
        );

    \I__10243\ : Odrv4
    port map (
            O => \N__45818\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_4\
        );

    \I__10242\ : InMux
    port map (
            O => \N__45815\,
            I => \N__45812\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__45812\,
            I => \N__45809\
        );

    \I__10240\ : Odrv4
    port map (
            O => \N__45809\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_0\
        );

    \I__10239\ : InMux
    port map (
            O => \N__45806\,
            I => \N__45803\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__45803\,
            I => \N__45800\
        );

    \I__10237\ : Odrv4
    port map (
            O => \N__45800\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_2\
        );

    \I__10236\ : InMux
    port map (
            O => \N__45797\,
            I => \N__45794\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__45794\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_2\
        );

    \I__10234\ : InMux
    port map (
            O => \N__45791\,
            I => \N__45788\
        );

    \I__10233\ : LocalMux
    port map (
            O => \N__45788\,
            I => \N__45785\
        );

    \I__10232\ : Odrv4
    port map (
            O => \N__45785\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_1\
        );

    \I__10231\ : InMux
    port map (
            O => \N__45782\,
            I => \N__45779\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__45779\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_1\
        );

    \I__10229\ : InMux
    port map (
            O => \N__45776\,
            I => \N__45773\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__45773\,
            I => \N__45768\
        );

    \I__10227\ : InMux
    port map (
            O => \N__45772\,
            I => \N__45765\
        );

    \I__10226\ : InMux
    port map (
            O => \N__45771\,
            I => \N__45762\
        );

    \I__10225\ : Span12Mux_h
    port map (
            O => \N__45768\,
            I => \N__45757\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45757\
        );

    \I__10223\ : LocalMux
    port map (
            O => \N__45762\,
            I => \button_debounce_counterZ0Z_1\
        );

    \I__10222\ : Odrv12
    port map (
            O => \N__45757\,
            I => \button_debounce_counterZ0Z_1\
        );

    \I__10221\ : InMux
    port map (
            O => \N__45752\,
            I => \N__45748\
        );

    \I__10220\ : CascadeMux
    port map (
            O => \N__45751\,
            I => \N__45745\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__45748\,
            I => \N__45740\
        );

    \I__10218\ : InMux
    port map (
            O => \N__45745\,
            I => \N__45737\
        );

    \I__10217\ : InMux
    port map (
            O => \N__45744\,
            I => \N__45732\
        );

    \I__10216\ : InMux
    port map (
            O => \N__45743\,
            I => \N__45732\
        );

    \I__10215\ : Span12Mux_h
    port map (
            O => \N__45740\,
            I => \N__45727\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__45737\,
            I => \N__45727\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__45732\,
            I => \button_debounce_counterZ0Z_0\
        );

    \I__10212\ : Odrv12
    port map (
            O => \N__45727\,
            I => \button_debounce_counterZ0Z_0\
        );

    \I__10211\ : InMux
    port map (
            O => \N__45722\,
            I => \N__45719\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__45719\,
            I => \N__45711\
        );

    \I__10209\ : SRMux
    port map (
            O => \N__45718\,
            I => \N__45698\
        );

    \I__10208\ : SRMux
    port map (
            O => \N__45717\,
            I => \N__45698\
        );

    \I__10207\ : SRMux
    port map (
            O => \N__45716\,
            I => \N__45698\
        );

    \I__10206\ : SRMux
    port map (
            O => \N__45715\,
            I => \N__45698\
        );

    \I__10205\ : SRMux
    port map (
            O => \N__45714\,
            I => \N__45698\
        );

    \I__10204\ : Glb2LocalMux
    port map (
            O => \N__45711\,
            I => \N__45698\
        );

    \I__10203\ : GlobalMux
    port map (
            O => \N__45698\,
            I => \N__45695\
        );

    \I__10202\ : gio2CtrlBuf
    port map (
            O => \N__45695\,
            I => \N_3154_g\
        );

    \I__10201\ : InMux
    port map (
            O => \N__45692\,
            I => \N__45689\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__45689\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_3\
        );

    \I__10199\ : InMux
    port map (
            O => \N__45686\,
            I => \N__45683\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__45683\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_3\
        );

    \I__10197\ : InMux
    port map (
            O => \N__45680\,
            I => \N__45677\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__45677\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_6\
        );

    \I__10195\ : InMux
    port map (
            O => \N__45674\,
            I => \N__45671\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__45671\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_6\
        );

    \I__10193\ : InMux
    port map (
            O => \N__45668\,
            I => \N__45665\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__45665\,
            I => \N__45662\
        );

    \I__10191\ : Span4Mux_v
    port map (
            O => \N__45662\,
            I => \N__45659\
        );

    \I__10190\ : Span4Mux_h
    port map (
            O => \N__45659\,
            I => \N__45656\
        );

    \I__10189\ : Odrv4
    port map (
            O => \N__45656\,
            I => \sDAC_mem_13Z0Z_0\
        );

    \I__10188\ : InMux
    port map (
            O => \N__45653\,
            I => \N__45650\
        );

    \I__10187\ : LocalMux
    port map (
            O => \N__45650\,
            I => \N__45647\
        );

    \I__10186\ : Span4Mux_v
    port map (
            O => \N__45647\,
            I => \N__45644\
        );

    \I__10185\ : Span4Mux_h
    port map (
            O => \N__45644\,
            I => \N__45641\
        );

    \I__10184\ : Odrv4
    port map (
            O => \N__45641\,
            I => \sDAC_mem_13Z0Z_1\
        );

    \I__10183\ : InMux
    port map (
            O => \N__45638\,
            I => \N__45635\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__45635\,
            I => \N__45632\
        );

    \I__10181\ : Span4Mux_h
    port map (
            O => \N__45632\,
            I => \N__45629\
        );

    \I__10180\ : Span4Mux_h
    port map (
            O => \N__45629\,
            I => \N__45626\
        );

    \I__10179\ : Odrv4
    port map (
            O => \N__45626\,
            I => \sDAC_mem_13Z0Z_2\
        );

    \I__10178\ : InMux
    port map (
            O => \N__45623\,
            I => \N__45620\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__45620\,
            I => \N__45617\
        );

    \I__10176\ : Span12Mux_h
    port map (
            O => \N__45617\,
            I => \N__45614\
        );

    \I__10175\ : Odrv12
    port map (
            O => \N__45614\,
            I => \sDAC_mem_13Z0Z_3\
        );

    \I__10174\ : InMux
    port map (
            O => \N__45611\,
            I => \N__45608\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__45608\,
            I => \N__45597\
        );

    \I__10172\ : InMux
    port map (
            O => \N__45607\,
            I => \N__45594\
        );

    \I__10171\ : InMux
    port map (
            O => \N__45606\,
            I => \N__45589\
        );

    \I__10170\ : InMux
    port map (
            O => \N__45605\,
            I => \N__45586\
        );

    \I__10169\ : InMux
    port map (
            O => \N__45604\,
            I => \N__45582\
        );

    \I__10168\ : InMux
    port map (
            O => \N__45603\,
            I => \N__45571\
        );

    \I__10167\ : InMux
    port map (
            O => \N__45602\,
            I => \N__45564\
        );

    \I__10166\ : InMux
    port map (
            O => \N__45601\,
            I => \N__45555\
        );

    \I__10165\ : InMux
    port map (
            O => \N__45600\,
            I => \N__45551\
        );

    \I__10164\ : Span4Mux_v
    port map (
            O => \N__45597\,
            I => \N__45546\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__45594\,
            I => \N__45546\
        );

    \I__10162\ : InMux
    port map (
            O => \N__45593\,
            I => \N__45543\
        );

    \I__10161\ : InMux
    port map (
            O => \N__45592\,
            I => \N__45540\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__45589\,
            I => \N__45535\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__45586\,
            I => \N__45535\
        );

    \I__10158\ : InMux
    port map (
            O => \N__45585\,
            I => \N__45532\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__45582\,
            I => \N__45525\
        );

    \I__10156\ : InMux
    port map (
            O => \N__45581\,
            I => \N__45522\
        );

    \I__10155\ : InMux
    port map (
            O => \N__45580\,
            I => \N__45519\
        );

    \I__10154\ : InMux
    port map (
            O => \N__45579\,
            I => \N__45516\
        );

    \I__10153\ : InMux
    port map (
            O => \N__45578\,
            I => \N__45513\
        );

    \I__10152\ : InMux
    port map (
            O => \N__45577\,
            I => \N__45510\
        );

    \I__10151\ : InMux
    port map (
            O => \N__45576\,
            I => \N__45503\
        );

    \I__10150\ : InMux
    port map (
            O => \N__45575\,
            I => \N__45500\
        );

    \I__10149\ : InMux
    port map (
            O => \N__45574\,
            I => \N__45497\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__45571\,
            I => \N__45494\
        );

    \I__10147\ : InMux
    port map (
            O => \N__45570\,
            I => \N__45491\
        );

    \I__10146\ : InMux
    port map (
            O => \N__45569\,
            I => \N__45488\
        );

    \I__10145\ : InMux
    port map (
            O => \N__45568\,
            I => \N__45485\
        );

    \I__10144\ : InMux
    port map (
            O => \N__45567\,
            I => \N__45482\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__45564\,
            I => \N__45478\
        );

    \I__10142\ : InMux
    port map (
            O => \N__45563\,
            I => \N__45475\
        );

    \I__10141\ : InMux
    port map (
            O => \N__45562\,
            I => \N__45472\
        );

    \I__10140\ : InMux
    port map (
            O => \N__45561\,
            I => \N__45469\
        );

    \I__10139\ : InMux
    port map (
            O => \N__45560\,
            I => \N__45466\
        );

    \I__10138\ : InMux
    port map (
            O => \N__45559\,
            I => \N__45463\
        );

    \I__10137\ : InMux
    port map (
            O => \N__45558\,
            I => \N__45460\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__45555\,
            I => \N__45457\
        );

    \I__10135\ : InMux
    port map (
            O => \N__45554\,
            I => \N__45454\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__45551\,
            I => \N__45451\
        );

    \I__10133\ : Span4Mux_v
    port map (
            O => \N__45546\,
            I => \N__45444\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__45543\,
            I => \N__45444\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__45540\,
            I => \N__45444\
        );

    \I__10130\ : Span4Mux_v
    port map (
            O => \N__45535\,
            I => \N__45439\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__45532\,
            I => \N__45439\
        );

    \I__10128\ : InMux
    port map (
            O => \N__45531\,
            I => \N__45436\
        );

    \I__10127\ : InMux
    port map (
            O => \N__45530\,
            I => \N__45433\
        );

    \I__10126\ : InMux
    port map (
            O => \N__45529\,
            I => \N__45430\
        );

    \I__10125\ : InMux
    port map (
            O => \N__45528\,
            I => \N__45427\
        );

    \I__10124\ : Span4Mux_v
    port map (
            O => \N__45525\,
            I => \N__45414\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__45522\,
            I => \N__45414\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__45519\,
            I => \N__45414\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__45516\,
            I => \N__45414\
        );

    \I__10120\ : LocalMux
    port map (
            O => \N__45513\,
            I => \N__45414\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__45510\,
            I => \N__45414\
        );

    \I__10118\ : InMux
    port map (
            O => \N__45509\,
            I => \N__45407\
        );

    \I__10117\ : InMux
    port map (
            O => \N__45508\,
            I => \N__45404\
        );

    \I__10116\ : InMux
    port map (
            O => \N__45507\,
            I => \N__45401\
        );

    \I__10115\ : InMux
    port map (
            O => \N__45506\,
            I => \N__45398\
        );

    \I__10114\ : LocalMux
    port map (
            O => \N__45503\,
            I => \N__45394\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__45500\,
            I => \N__45389\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__45497\,
            I => \N__45389\
        );

    \I__10111\ : Span4Mux_v
    port map (
            O => \N__45494\,
            I => \N__45384\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__45491\,
            I => \N__45375\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__45488\,
            I => \N__45375\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__45485\,
            I => \N__45375\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__45482\,
            I => \N__45375\
        );

    \I__10106\ : CascadeMux
    port map (
            O => \N__45481\,
            I => \N__45369\
        );

    \I__10105\ : Span4Mux_v
    port map (
            O => \N__45478\,
            I => \N__45360\
        );

    \I__10104\ : LocalMux
    port map (
            O => \N__45475\,
            I => \N__45360\
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__45472\,
            I => \N__45360\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__45469\,
            I => \N__45360\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__45466\,
            I => \N__45354\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__45463\,
            I => \N__45354\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__45460\,
            I => \N__45351\
        );

    \I__10098\ : Span4Mux_v
    port map (
            O => \N__45457\,
            I => \N__45343\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__45454\,
            I => \N__45343\
        );

    \I__10096\ : Span4Mux_v
    port map (
            O => \N__45451\,
            I => \N__45338\
        );

    \I__10095\ : Span4Mux_v
    port map (
            O => \N__45444\,
            I => \N__45338\
        );

    \I__10094\ : Span4Mux_v
    port map (
            O => \N__45439\,
            I => \N__45333\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__45436\,
            I => \N__45333\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__45433\,
            I => \N__45326\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__45430\,
            I => \N__45326\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__45427\,
            I => \N__45326\
        );

    \I__10089\ : Span4Mux_v
    port map (
            O => \N__45414\,
            I => \N__45323\
        );

    \I__10088\ : InMux
    port map (
            O => \N__45413\,
            I => \N__45320\
        );

    \I__10087\ : InMux
    port map (
            O => \N__45412\,
            I => \N__45317\
        );

    \I__10086\ : InMux
    port map (
            O => \N__45411\,
            I => \N__45314\
        );

    \I__10085\ : InMux
    port map (
            O => \N__45410\,
            I => \N__45311\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__45407\,
            I => \N__45308\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__45404\,
            I => \N__45301\
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__45401\,
            I => \N__45301\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__45398\,
            I => \N__45301\
        );

    \I__10080\ : InMux
    port map (
            O => \N__45397\,
            I => \N__45298\
        );

    \I__10079\ : Span4Mux_v
    port map (
            O => \N__45394\,
            I => \N__45291\
        );

    \I__10078\ : Span4Mux_v
    port map (
            O => \N__45389\,
            I => \N__45291\
        );

    \I__10077\ : InMux
    port map (
            O => \N__45388\,
            I => \N__45288\
        );

    \I__10076\ : InMux
    port map (
            O => \N__45387\,
            I => \N__45285\
        );

    \I__10075\ : Span4Mux_h
    port map (
            O => \N__45384\,
            I => \N__45280\
        );

    \I__10074\ : Span4Mux_v
    port map (
            O => \N__45375\,
            I => \N__45280\
        );

    \I__10073\ : InMux
    port map (
            O => \N__45374\,
            I => \N__45277\
        );

    \I__10072\ : InMux
    port map (
            O => \N__45373\,
            I => \N__45274\
        );

    \I__10071\ : InMux
    port map (
            O => \N__45372\,
            I => \N__45271\
        );

    \I__10070\ : InMux
    port map (
            O => \N__45369\,
            I => \N__45268\
        );

    \I__10069\ : Sp12to4
    port map (
            O => \N__45360\,
            I => \N__45265\
        );

    \I__10068\ : InMux
    port map (
            O => \N__45359\,
            I => \N__45262\
        );

    \I__10067\ : Span4Mux_v
    port map (
            O => \N__45354\,
            I => \N__45257\
        );

    \I__10066\ : Span4Mux_v
    port map (
            O => \N__45351\,
            I => \N__45257\
        );

    \I__10065\ : InMux
    port map (
            O => \N__45350\,
            I => \N__45254\
        );

    \I__10064\ : InMux
    port map (
            O => \N__45349\,
            I => \N__45251\
        );

    \I__10063\ : InMux
    port map (
            O => \N__45348\,
            I => \N__45248\
        );

    \I__10062\ : Span4Mux_v
    port map (
            O => \N__45343\,
            I => \N__45245\
        );

    \I__10061\ : Span4Mux_h
    port map (
            O => \N__45338\,
            I => \N__45238\
        );

    \I__10060\ : Span4Mux_v
    port map (
            O => \N__45333\,
            I => \N__45238\
        );

    \I__10059\ : Span4Mux_v
    port map (
            O => \N__45326\,
            I => \N__45238\
        );

    \I__10058\ : Span4Mux_v
    port map (
            O => \N__45323\,
            I => \N__45227\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__45320\,
            I => \N__45227\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__45317\,
            I => \N__45227\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__45314\,
            I => \N__45227\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__45311\,
            I => \N__45227\
        );

    \I__10053\ : Span4Mux_v
    port map (
            O => \N__45308\,
            I => \N__45221\
        );

    \I__10052\ : Span4Mux_v
    port map (
            O => \N__45301\,
            I => \N__45218\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__45298\,
            I => \N__45215\
        );

    \I__10050\ : InMux
    port map (
            O => \N__45297\,
            I => \N__45212\
        );

    \I__10049\ : InMux
    port map (
            O => \N__45296\,
            I => \N__45209\
        );

    \I__10048\ : Span4Mux_v
    port map (
            O => \N__45291\,
            I => \N__45202\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__45288\,
            I => \N__45202\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__45285\,
            I => \N__45202\
        );

    \I__10045\ : Span4Mux_v
    port map (
            O => \N__45280\,
            I => \N__45191\
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__45277\,
            I => \N__45191\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__45274\,
            I => \N__45191\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__45271\,
            I => \N__45191\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__45268\,
            I => \N__45191\
        );

    \I__10040\ : Span12Mux_v
    port map (
            O => \N__45265\,
            I => \N__45178\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__45262\,
            I => \N__45178\
        );

    \I__10038\ : Sp12to4
    port map (
            O => \N__45257\,
            I => \N__45178\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__45254\,
            I => \N__45178\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__45251\,
            I => \N__45178\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__45248\,
            I => \N__45178\
        );

    \I__10034\ : Span4Mux_v
    port map (
            O => \N__45245\,
            I => \N__45171\
        );

    \I__10033\ : Span4Mux_h
    port map (
            O => \N__45238\,
            I => \N__45171\
        );

    \I__10032\ : Span4Mux_v
    port map (
            O => \N__45227\,
            I => \N__45171\
        );

    \I__10031\ : InMux
    port map (
            O => \N__45226\,
            I => \N__45168\
        );

    \I__10030\ : InMux
    port map (
            O => \N__45225\,
            I => \N__45165\
        );

    \I__10029\ : InMux
    port map (
            O => \N__45224\,
            I => \N__45162\
        );

    \I__10028\ : Span4Mux_h
    port map (
            O => \N__45221\,
            I => \N__45147\
        );

    \I__10027\ : Span4Mux_h
    port map (
            O => \N__45218\,
            I => \N__45147\
        );

    \I__10026\ : Span4Mux_v
    port map (
            O => \N__45215\,
            I => \N__45147\
        );

    \I__10025\ : LocalMux
    port map (
            O => \N__45212\,
            I => \N__45147\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__45209\,
            I => \N__45147\
        );

    \I__10023\ : Span4Mux_v
    port map (
            O => \N__45202\,
            I => \N__45147\
        );

    \I__10022\ : Span4Mux_v
    port map (
            O => \N__45191\,
            I => \N__45147\
        );

    \I__10021\ : Odrv12
    port map (
            O => \N__45178\,
            I => spi_data_mosi_4
        );

    \I__10020\ : Odrv4
    port map (
            O => \N__45171\,
            I => spi_data_mosi_4
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__45168\,
            I => spi_data_mosi_4
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__45165\,
            I => spi_data_mosi_4
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__45162\,
            I => spi_data_mosi_4
        );

    \I__10016\ : Odrv4
    port map (
            O => \N__45147\,
            I => spi_data_mosi_4
        );

    \I__10015\ : InMux
    port map (
            O => \N__45134\,
            I => \N__45131\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__45131\,
            I => \N__45128\
        );

    \I__10013\ : Span4Mux_v
    port map (
            O => \N__45128\,
            I => \N__45125\
        );

    \I__10012\ : Span4Mux_h
    port map (
            O => \N__45125\,
            I => \N__45122\
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__45122\,
            I => \sDAC_mem_13Z0Z_4\
        );

    \I__10010\ : InMux
    port map (
            O => \N__45119\,
            I => \N__45111\
        );

    \I__10009\ : InMux
    port map (
            O => \N__45118\,
            I => \N__45108\
        );

    \I__10008\ : InMux
    port map (
            O => \N__45117\,
            I => \N__45097\
        );

    \I__10007\ : InMux
    port map (
            O => \N__45116\,
            I => \N__45091\
        );

    \I__10006\ : InMux
    port map (
            O => \N__45115\,
            I => \N__45086\
        );

    \I__10005\ : InMux
    port map (
            O => \N__45114\,
            I => \N__45082\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__45111\,
            I => \N__45072\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__45108\,
            I => \N__45072\
        );

    \I__10002\ : InMux
    port map (
            O => \N__45107\,
            I => \N__45069\
        );

    \I__10001\ : InMux
    port map (
            O => \N__45106\,
            I => \N__45061\
        );

    \I__10000\ : InMux
    port map (
            O => \N__45105\,
            I => \N__45058\
        );

    \I__9999\ : InMux
    port map (
            O => \N__45104\,
            I => \N__45050\
        );

    \I__9998\ : InMux
    port map (
            O => \N__45103\,
            I => \N__45047\
        );

    \I__9997\ : InMux
    port map (
            O => \N__45102\,
            I => \N__45044\
        );

    \I__9996\ : InMux
    port map (
            O => \N__45101\,
            I => \N__45041\
        );

    \I__9995\ : InMux
    port map (
            O => \N__45100\,
            I => \N__45038\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__45097\,
            I => \N__45034\
        );

    \I__9993\ : InMux
    port map (
            O => \N__45096\,
            I => \N__45031\
        );

    \I__9992\ : InMux
    port map (
            O => \N__45095\,
            I => \N__45028\
        );

    \I__9991\ : InMux
    port map (
            O => \N__45094\,
            I => \N__45025\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__45091\,
            I => \N__45022\
        );

    \I__9989\ : InMux
    port map (
            O => \N__45090\,
            I => \N__45019\
        );

    \I__9988\ : InMux
    port map (
            O => \N__45089\,
            I => \N__45016\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__45086\,
            I => \N__45013\
        );

    \I__9986\ : InMux
    port map (
            O => \N__45085\,
            I => \N__45010\
        );

    \I__9985\ : LocalMux
    port map (
            O => \N__45082\,
            I => \N__45006\
        );

    \I__9984\ : InMux
    port map (
            O => \N__45081\,
            I => \N__45002\
        );

    \I__9983\ : InMux
    port map (
            O => \N__45080\,
            I => \N__44997\
        );

    \I__9982\ : InMux
    port map (
            O => \N__45079\,
            I => \N__44994\
        );

    \I__9981\ : InMux
    port map (
            O => \N__45078\,
            I => \N__44991\
        );

    \I__9980\ : InMux
    port map (
            O => \N__45077\,
            I => \N__44988\
        );

    \I__9979\ : Span4Mux_h
    port map (
            O => \N__45072\,
            I => \N__44983\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__45069\,
            I => \N__44983\
        );

    \I__9977\ : InMux
    port map (
            O => \N__45068\,
            I => \N__44977\
        );

    \I__9976\ : InMux
    port map (
            O => \N__45067\,
            I => \N__44974\
        );

    \I__9975\ : InMux
    port map (
            O => \N__45066\,
            I => \N__44971\
        );

    \I__9974\ : InMux
    port map (
            O => \N__45065\,
            I => \N__44968\
        );

    \I__9973\ : InMux
    port map (
            O => \N__45064\,
            I => \N__44965\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__45061\,
            I => \N__44962\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__45058\,
            I => \N__44959\
        );

    \I__9970\ : InMux
    port map (
            O => \N__45057\,
            I => \N__44956\
        );

    \I__9969\ : InMux
    port map (
            O => \N__45056\,
            I => \N__44953\
        );

    \I__9968\ : InMux
    port map (
            O => \N__45055\,
            I => \N__44948\
        );

    \I__9967\ : InMux
    port map (
            O => \N__45054\,
            I => \N__44945\
        );

    \I__9966\ : InMux
    port map (
            O => \N__45053\,
            I => \N__44942\
        );

    \I__9965\ : LocalMux
    port map (
            O => \N__45050\,
            I => \N__44939\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__45047\,
            I => \N__44930\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__45044\,
            I => \N__44930\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__45041\,
            I => \N__44930\
        );

    \I__9961\ : LocalMux
    port map (
            O => \N__45038\,
            I => \N__44930\
        );

    \I__9960\ : InMux
    port map (
            O => \N__45037\,
            I => \N__44925\
        );

    \I__9959\ : Span4Mux_v
    port map (
            O => \N__45034\,
            I => \N__44920\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__45031\,
            I => \N__44915\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__45028\,
            I => \N__44915\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__45025\,
            I => \N__44908\
        );

    \I__9955\ : Span4Mux_v
    port map (
            O => \N__45022\,
            I => \N__44908\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__45019\,
            I => \N__44908\
        );

    \I__9953\ : LocalMux
    port map (
            O => \N__45016\,
            I => \N__44905\
        );

    \I__9952\ : Span4Mux_h
    port map (
            O => \N__45013\,
            I => \N__44902\
        );

    \I__9951\ : LocalMux
    port map (
            O => \N__45010\,
            I => \N__44899\
        );

    \I__9950\ : InMux
    port map (
            O => \N__45009\,
            I => \N__44896\
        );

    \I__9949\ : Span4Mux_h
    port map (
            O => \N__45006\,
            I => \N__44893\
        );

    \I__9948\ : InMux
    port map (
            O => \N__45005\,
            I => \N__44890\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__45002\,
            I => \N__44887\
        );

    \I__9946\ : InMux
    port map (
            O => \N__45001\,
            I => \N__44884\
        );

    \I__9945\ : InMux
    port map (
            O => \N__45000\,
            I => \N__44881\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__44997\,
            I => \N__44876\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__44994\,
            I => \N__44876\
        );

    \I__9942\ : LocalMux
    port map (
            O => \N__44991\,
            I => \N__44871\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__44988\,
            I => \N__44871\
        );

    \I__9940\ : Span4Mux_v
    port map (
            O => \N__44983\,
            I => \N__44868\
        );

    \I__9939\ : InMux
    port map (
            O => \N__44982\,
            I => \N__44864\
        );

    \I__9938\ : InMux
    port map (
            O => \N__44981\,
            I => \N__44861\
        );

    \I__9937\ : InMux
    port map (
            O => \N__44980\,
            I => \N__44858\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__44977\,
            I => \N__44853\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__44974\,
            I => \N__44853\
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__44971\,
            I => \N__44842\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__44968\,
            I => \N__44842\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__44965\,
            I => \N__44842\
        );

    \I__9931\ : Span4Mux_h
    port map (
            O => \N__44962\,
            I => \N__44842\
        );

    \I__9930\ : Span4Mux_v
    port map (
            O => \N__44959\,
            I => \N__44842\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__44956\,
            I => \N__44835\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__44953\,
            I => \N__44835\
        );

    \I__9927\ : InMux
    port map (
            O => \N__44952\,
            I => \N__44830\
        );

    \I__9926\ : InMux
    port map (
            O => \N__44951\,
            I => \N__44827\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__44948\,
            I => \N__44820\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__44945\,
            I => \N__44820\
        );

    \I__9923\ : LocalMux
    port map (
            O => \N__44942\,
            I => \N__44820\
        );

    \I__9922\ : Span4Mux_v
    port map (
            O => \N__44939\,
            I => \N__44815\
        );

    \I__9921\ : Span4Mux_v
    port map (
            O => \N__44930\,
            I => \N__44815\
        );

    \I__9920\ : InMux
    port map (
            O => \N__44929\,
            I => \N__44812\
        );

    \I__9919\ : InMux
    port map (
            O => \N__44928\,
            I => \N__44809\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__44925\,
            I => \N__44806\
        );

    \I__9917\ : InMux
    port map (
            O => \N__44924\,
            I => \N__44803\
        );

    \I__9916\ : InMux
    port map (
            O => \N__44923\,
            I => \N__44800\
        );

    \I__9915\ : Span4Mux_h
    port map (
            O => \N__44920\,
            I => \N__44793\
        );

    \I__9914\ : Span4Mux_v
    port map (
            O => \N__44915\,
            I => \N__44793\
        );

    \I__9913\ : Span4Mux_v
    port map (
            O => \N__44908\,
            I => \N__44793\
        );

    \I__9912\ : Span4Mux_v
    port map (
            O => \N__44905\,
            I => \N__44788\
        );

    \I__9911\ : Span4Mux_h
    port map (
            O => \N__44902\,
            I => \N__44788\
        );

    \I__9910\ : Span4Mux_v
    port map (
            O => \N__44899\,
            I => \N__44781\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__44896\,
            I => \N__44781\
        );

    \I__9908\ : Span4Mux_h
    port map (
            O => \N__44893\,
            I => \N__44781\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__44890\,
            I => \N__44774\
        );

    \I__9906\ : Span4Mux_h
    port map (
            O => \N__44887\,
            I => \N__44774\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__44884\,
            I => \N__44774\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__44881\,
            I => \N__44771\
        );

    \I__9903\ : Span4Mux_v
    port map (
            O => \N__44876\,
            I => \N__44764\
        );

    \I__9902\ : Span4Mux_v
    port map (
            O => \N__44871\,
            I => \N__44764\
        );

    \I__9901\ : Span4Mux_h
    port map (
            O => \N__44868\,
            I => \N__44764\
        );

    \I__9900\ : InMux
    port map (
            O => \N__44867\,
            I => \N__44760\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__44864\,
            I => \N__44753\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__44861\,
            I => \N__44753\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__44858\,
            I => \N__44753\
        );

    \I__9896\ : Span4Mux_v
    port map (
            O => \N__44853\,
            I => \N__44748\
        );

    \I__9895\ : Span4Mux_v
    port map (
            O => \N__44842\,
            I => \N__44748\
        );

    \I__9894\ : InMux
    port map (
            O => \N__44841\,
            I => \N__44745\
        );

    \I__9893\ : InMux
    port map (
            O => \N__44840\,
            I => \N__44742\
        );

    \I__9892\ : Span4Mux_v
    port map (
            O => \N__44835\,
            I => \N__44739\
        );

    \I__9891\ : InMux
    port map (
            O => \N__44834\,
            I => \N__44734\
        );

    \I__9890\ : InMux
    port map (
            O => \N__44833\,
            I => \N__44734\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__44830\,
            I => \N__44727\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__44827\,
            I => \N__44720\
        );

    \I__9887\ : Span4Mux_v
    port map (
            O => \N__44820\,
            I => \N__44720\
        );

    \I__9886\ : Span4Mux_h
    port map (
            O => \N__44815\,
            I => \N__44720\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__44812\,
            I => \N__44707\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__44809\,
            I => \N__44707\
        );

    \I__9883\ : Span4Mux_h
    port map (
            O => \N__44806\,
            I => \N__44707\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__44803\,
            I => \N__44707\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__44800\,
            I => \N__44707\
        );

    \I__9880\ : Span4Mux_v
    port map (
            O => \N__44793\,
            I => \N__44707\
        );

    \I__9879\ : Span4Mux_h
    port map (
            O => \N__44788\,
            I => \N__44702\
        );

    \I__9878\ : Span4Mux_v
    port map (
            O => \N__44781\,
            I => \N__44702\
        );

    \I__9877\ : Span4Mux_v
    port map (
            O => \N__44774\,
            I => \N__44699\
        );

    \I__9876\ : Span4Mux_h
    port map (
            O => \N__44771\,
            I => \N__44694\
        );

    \I__9875\ : Span4Mux_h
    port map (
            O => \N__44764\,
            I => \N__44694\
        );

    \I__9874\ : InMux
    port map (
            O => \N__44763\,
            I => \N__44691\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__44760\,
            I => \N__44684\
        );

    \I__9872\ : Span4Mux_v
    port map (
            O => \N__44753\,
            I => \N__44684\
        );

    \I__9871\ : Span4Mux_h
    port map (
            O => \N__44748\,
            I => \N__44684\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__44745\,
            I => \N__44675\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__44742\,
            I => \N__44675\
        );

    \I__9868\ : Span4Mux_v
    port map (
            O => \N__44739\,
            I => \N__44675\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__44734\,
            I => \N__44675\
        );

    \I__9866\ : InMux
    port map (
            O => \N__44733\,
            I => \N__44672\
        );

    \I__9865\ : InMux
    port map (
            O => \N__44732\,
            I => \N__44669\
        );

    \I__9864\ : InMux
    port map (
            O => \N__44731\,
            I => \N__44666\
        );

    \I__9863\ : InMux
    port map (
            O => \N__44730\,
            I => \N__44663\
        );

    \I__9862\ : Span4Mux_v
    port map (
            O => \N__44727\,
            I => \N__44656\
        );

    \I__9861\ : Span4Mux_h
    port map (
            O => \N__44720\,
            I => \N__44656\
        );

    \I__9860\ : Span4Mux_v
    port map (
            O => \N__44707\,
            I => \N__44656\
        );

    \I__9859\ : Span4Mux_v
    port map (
            O => \N__44702\,
            I => \N__44653\
        );

    \I__9858\ : Span4Mux_h
    port map (
            O => \N__44699\,
            I => \N__44648\
        );

    \I__9857\ : Span4Mux_v
    port map (
            O => \N__44694\,
            I => \N__44648\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__44691\,
            I => \N__44641\
        );

    \I__9855\ : Span4Mux_h
    port map (
            O => \N__44684\,
            I => \N__44641\
        );

    \I__9854\ : Span4Mux_v
    port map (
            O => \N__44675\,
            I => \N__44641\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__44672\,
            I => spi_data_mosi_5
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__44669\,
            I => spi_data_mosi_5
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__44666\,
            I => spi_data_mosi_5
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__44663\,
            I => spi_data_mosi_5
        );

    \I__9849\ : Odrv4
    port map (
            O => \N__44656\,
            I => spi_data_mosi_5
        );

    \I__9848\ : Odrv4
    port map (
            O => \N__44653\,
            I => spi_data_mosi_5
        );

    \I__9847\ : Odrv4
    port map (
            O => \N__44648\,
            I => spi_data_mosi_5
        );

    \I__9846\ : Odrv4
    port map (
            O => \N__44641\,
            I => spi_data_mosi_5
        );

    \I__9845\ : InMux
    port map (
            O => \N__44624\,
            I => \N__44621\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__44621\,
            I => \N__44618\
        );

    \I__9843\ : Span4Mux_v
    port map (
            O => \N__44618\,
            I => \N__44615\
        );

    \I__9842\ : Span4Mux_h
    port map (
            O => \N__44615\,
            I => \N__44612\
        );

    \I__9841\ : Odrv4
    port map (
            O => \N__44612\,
            I => \sDAC_mem_13Z0Z_5\
        );

    \I__9840\ : InMux
    port map (
            O => \N__44609\,
            I => \N__44606\
        );

    \I__9839\ : LocalMux
    port map (
            O => \N__44606\,
            I => \N__44603\
        );

    \I__9838\ : Span4Mux_h
    port map (
            O => \N__44603\,
            I => \N__44600\
        );

    \I__9837\ : Odrv4
    port map (
            O => \N__44600\,
            I => \sDAC_mem_13Z0Z_6\
        );

    \I__9836\ : InMux
    port map (
            O => \N__44597\,
            I => \N__44594\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__44594\,
            I => \N__44591\
        );

    \I__9834\ : Span4Mux_v
    port map (
            O => \N__44591\,
            I => \N__44588\
        );

    \I__9833\ : Odrv4
    port map (
            O => \N__44588\,
            I => \sDAC_mem_13Z0Z_7\
        );

    \I__9832\ : CEMux
    port map (
            O => \N__44585\,
            I => \N__44582\
        );

    \I__9831\ : LocalMux
    port map (
            O => \N__44582\,
            I => \N__44579\
        );

    \I__9830\ : Span4Mux_h
    port map (
            O => \N__44579\,
            I => \N__44576\
        );

    \I__9829\ : Span4Mux_h
    port map (
            O => \N__44576\,
            I => \N__44573\
        );

    \I__9828\ : Odrv4
    port map (
            O => \N__44573\,
            I => \sDAC_mem_13_1_sqmuxa\
        );

    \I__9827\ : InMux
    port map (
            O => \N__44570\,
            I => \N__44567\
        );

    \I__9826\ : LocalMux
    port map (
            O => \N__44567\,
            I => \N__44564\
        );

    \I__9825\ : Span4Mux_v
    port map (
            O => \N__44564\,
            I => \N__44561\
        );

    \I__9824\ : Span4Mux_h
    port map (
            O => \N__44561\,
            I => \N__44558\
        );

    \I__9823\ : Span4Mux_v
    port map (
            O => \N__44558\,
            I => \N__44554\
        );

    \I__9822\ : InMux
    port map (
            O => \N__44557\,
            I => \N__44551\
        );

    \I__9821\ : Span4Mux_h
    port map (
            O => \N__44554\,
            I => \N__44548\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__44551\,
            I => \spi_slave_inst.tx_ready_iZ0\
        );

    \I__9819\ : Odrv4
    port map (
            O => \N__44548\,
            I => \spi_slave_inst.tx_ready_iZ0\
        );

    \I__9818\ : InMux
    port map (
            O => \N__44543\,
            I => \N__44540\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__44540\,
            I => \N__44537\
        );

    \I__9816\ : Span4Mux_v
    port map (
            O => \N__44537\,
            I => \N__44534\
        );

    \I__9815\ : Odrv4
    port map (
            O => \N__44534\,
            I => \sDAC_mem_33Z0Z_7\
        );

    \I__9814\ : CEMux
    port map (
            O => \N__44531\,
            I => \N__44528\
        );

    \I__9813\ : LocalMux
    port map (
            O => \N__44528\,
            I => \N__44525\
        );

    \I__9812\ : Odrv4
    port map (
            O => \N__44525\,
            I => \sDAC_mem_33_1_sqmuxa\
        );

    \I__9811\ : InMux
    port map (
            O => \N__44522\,
            I => \N__44519\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__44519\,
            I => \N__44516\
        );

    \I__9809\ : Odrv4
    port map (
            O => \N__44516\,
            I => \sDAC_mem_5Z0Z_0\
        );

    \I__9808\ : InMux
    port map (
            O => \N__44513\,
            I => \N__44510\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__44510\,
            I => \N__44507\
        );

    \I__9806\ : Odrv4
    port map (
            O => \N__44507\,
            I => \sDAC_mem_5Z0Z_1\
        );

    \I__9805\ : InMux
    port map (
            O => \N__44504\,
            I => \N__44501\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__44501\,
            I => \N__44498\
        );

    \I__9803\ : Odrv4
    port map (
            O => \N__44498\,
            I => \sDAC_mem_5Z0Z_2\
        );

    \I__9802\ : InMux
    port map (
            O => \N__44495\,
            I => \N__44492\
        );

    \I__9801\ : LocalMux
    port map (
            O => \N__44492\,
            I => \N__44489\
        );

    \I__9800\ : Span4Mux_h
    port map (
            O => \N__44489\,
            I => \N__44486\
        );

    \I__9799\ : Odrv4
    port map (
            O => \N__44486\,
            I => \sDAC_mem_5Z0Z_3\
        );

    \I__9798\ : InMux
    port map (
            O => \N__44483\,
            I => \N__44480\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__44480\,
            I => \N__44477\
        );

    \I__9796\ : Span4Mux_h
    port map (
            O => \N__44477\,
            I => \N__44474\
        );

    \I__9795\ : Odrv4
    port map (
            O => \N__44474\,
            I => \sDAC_mem_5Z0Z_4\
        );

    \I__9794\ : InMux
    port map (
            O => \N__44471\,
            I => \N__44468\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__44468\,
            I => \N__44465\
        );

    \I__9792\ : Span4Mux_h
    port map (
            O => \N__44465\,
            I => \N__44462\
        );

    \I__9791\ : Odrv4
    port map (
            O => \N__44462\,
            I => \sDAC_mem_5Z0Z_5\
        );

    \I__9790\ : InMux
    port map (
            O => \N__44459\,
            I => \N__44456\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__44456\,
            I => \N__44453\
        );

    \I__9788\ : Span4Mux_v
    port map (
            O => \N__44453\,
            I => \N__44450\
        );

    \I__9787\ : Odrv4
    port map (
            O => \N__44450\,
            I => \sDAC_mem_5Z0Z_6\
        );

    \I__9786\ : InMux
    port map (
            O => \N__44447\,
            I => \N__44444\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__44444\,
            I => \N__44441\
        );

    \I__9784\ : Span4Mux_h
    port map (
            O => \N__44441\,
            I => \N__44438\
        );

    \I__9783\ : Odrv4
    port map (
            O => \N__44438\,
            I => \sDAC_mem_5Z0Z_7\
        );

    \I__9782\ : CEMux
    port map (
            O => \N__44435\,
            I => \N__44432\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__44432\,
            I => \N__44429\
        );

    \I__9780\ : Span12Mux_s10_h
    port map (
            O => \N__44429\,
            I => \N__44426\
        );

    \I__9779\ : Odrv12
    port map (
            O => \N__44426\,
            I => \sDAC_mem_5_1_sqmuxa\
        );

    \I__9778\ : InMux
    port map (
            O => \N__44423\,
            I => \N__44420\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__44420\,
            I => \N__44417\
        );

    \I__9776\ : Odrv4
    port map (
            O => \N__44417\,
            I => \sDAC_mem_1Z0Z_6\
        );

    \I__9775\ : InMux
    port map (
            O => \N__44414\,
            I => \N__44411\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__44411\,
            I => \N__44408\
        );

    \I__9773\ : Span12Mux_v
    port map (
            O => \N__44408\,
            I => \N__44405\
        );

    \I__9772\ : Odrv12
    port map (
            O => \N__44405\,
            I => \sDAC_mem_1Z0Z_7\
        );

    \I__9771\ : CEMux
    port map (
            O => \N__44402\,
            I => \N__44399\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__44399\,
            I => \N__44396\
        );

    \I__9769\ : Span4Mux_v
    port map (
            O => \N__44396\,
            I => \N__44393\
        );

    \I__9768\ : Odrv4
    port map (
            O => \N__44393\,
            I => \sDAC_mem_1_1_sqmuxa\
        );

    \I__9767\ : InMux
    port map (
            O => \N__44390\,
            I => \N__44387\
        );

    \I__9766\ : LocalMux
    port map (
            O => \N__44387\,
            I => \N__44384\
        );

    \I__9765\ : Span4Mux_h
    port map (
            O => \N__44384\,
            I => \N__44381\
        );

    \I__9764\ : Odrv4
    port map (
            O => \N__44381\,
            I => \sDAC_mem_33Z0Z_0\
        );

    \I__9763\ : InMux
    port map (
            O => \N__44378\,
            I => \N__44375\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__44375\,
            I => \N__44372\
        );

    \I__9761\ : Odrv4
    port map (
            O => \N__44372\,
            I => \sDAC_mem_33Z0Z_1\
        );

    \I__9760\ : InMux
    port map (
            O => \N__44369\,
            I => \N__44366\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__44366\,
            I => \N__44363\
        );

    \I__9758\ : Odrv4
    port map (
            O => \N__44363\,
            I => \sDAC_mem_33Z0Z_2\
        );

    \I__9757\ : InMux
    port map (
            O => \N__44360\,
            I => \N__44357\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__44357\,
            I => \N__44354\
        );

    \I__9755\ : Span4Mux_h
    port map (
            O => \N__44354\,
            I => \N__44351\
        );

    \I__9754\ : Odrv4
    port map (
            O => \N__44351\,
            I => \sDAC_mem_33Z0Z_3\
        );

    \I__9753\ : InMux
    port map (
            O => \N__44348\,
            I => \N__44345\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__44345\,
            I => \N__44342\
        );

    \I__9751\ : Span4Mux_h
    port map (
            O => \N__44342\,
            I => \N__44339\
        );

    \I__9750\ : Odrv4
    port map (
            O => \N__44339\,
            I => \sDAC_mem_33Z0Z_4\
        );

    \I__9749\ : InMux
    port map (
            O => \N__44336\,
            I => \N__44333\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__44333\,
            I => \N__44330\
        );

    \I__9747\ : Span4Mux_h
    port map (
            O => \N__44330\,
            I => \N__44327\
        );

    \I__9746\ : Odrv4
    port map (
            O => \N__44327\,
            I => \sDAC_mem_33Z0Z_5\
        );

    \I__9745\ : InMux
    port map (
            O => \N__44324\,
            I => \N__44321\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__44321\,
            I => \N__44318\
        );

    \I__9743\ : Span4Mux_h
    port map (
            O => \N__44318\,
            I => \N__44315\
        );

    \I__9742\ : Odrv4
    port map (
            O => \N__44315\,
            I => \sDAC_mem_33Z0Z_6\
        );

    \I__9741\ : InMux
    port map (
            O => \N__44312\,
            I => \N__44309\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__44309\,
            I => \N__44306\
        );

    \I__9739\ : Span4Mux_h
    port map (
            O => \N__44306\,
            I => \N__44303\
        );

    \I__9738\ : Span4Mux_h
    port map (
            O => \N__44303\,
            I => \N__44300\
        );

    \I__9737\ : Odrv4
    port map (
            O => \N__44300\,
            I => \sDAC_mem_7Z0Z_4\
        );

    \I__9736\ : InMux
    port map (
            O => \N__44297\,
            I => \N__44294\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__44294\,
            I => \N__44291\
        );

    \I__9734\ : Span4Mux_v
    port map (
            O => \N__44291\,
            I => \N__44288\
        );

    \I__9733\ : Odrv4
    port map (
            O => \N__44288\,
            I => \sDAC_mem_7Z0Z_6\
        );

    \I__9732\ : CEMux
    port map (
            O => \N__44285\,
            I => \N__44282\
        );

    \I__9731\ : LocalMux
    port map (
            O => \N__44282\,
            I => \N__44279\
        );

    \I__9730\ : Span4Mux_h
    port map (
            O => \N__44279\,
            I => \N__44275\
        );

    \I__9729\ : CEMux
    port map (
            O => \N__44278\,
            I => \N__44272\
        );

    \I__9728\ : Span4Mux_h
    port map (
            O => \N__44275\,
            I => \N__44267\
        );

    \I__9727\ : LocalMux
    port map (
            O => \N__44272\,
            I => \N__44267\
        );

    \I__9726\ : Span4Mux_v
    port map (
            O => \N__44267\,
            I => \N__44264\
        );

    \I__9725\ : Odrv4
    port map (
            O => \N__44264\,
            I => \sDAC_mem_7_1_sqmuxa\
        );

    \I__9724\ : InMux
    port map (
            O => \N__44261\,
            I => \N__44258\
        );

    \I__9723\ : LocalMux
    port map (
            O => \N__44258\,
            I => \N__44255\
        );

    \I__9722\ : Span4Mux_h
    port map (
            O => \N__44255\,
            I => \N__44252\
        );

    \I__9721\ : Span4Mux_v
    port map (
            O => \N__44252\,
            I => \N__44249\
        );

    \I__9720\ : Odrv4
    port map (
            O => \N__44249\,
            I => \sDAC_mem_3Z0Z_7\
        );

    \I__9719\ : CEMux
    port map (
            O => \N__44246\,
            I => \N__44240\
        );

    \I__9718\ : CEMux
    port map (
            O => \N__44245\,
            I => \N__44234\
        );

    \I__9717\ : CEMux
    port map (
            O => \N__44244\,
            I => \N__44231\
        );

    \I__9716\ : CEMux
    port map (
            O => \N__44243\,
            I => \N__44228\
        );

    \I__9715\ : LocalMux
    port map (
            O => \N__44240\,
            I => \N__44225\
        );

    \I__9714\ : CEMux
    port map (
            O => \N__44239\,
            I => \N__44221\
        );

    \I__9713\ : CEMux
    port map (
            O => \N__44238\,
            I => \N__44218\
        );

    \I__9712\ : CEMux
    port map (
            O => \N__44237\,
            I => \N__44215\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__44234\,
            I => \N__44212\
        );

    \I__9710\ : LocalMux
    port map (
            O => \N__44231\,
            I => \N__44209\
        );

    \I__9709\ : LocalMux
    port map (
            O => \N__44228\,
            I => \N__44206\
        );

    \I__9708\ : Span4Mux_h
    port map (
            O => \N__44225\,
            I => \N__44203\
        );

    \I__9707\ : CEMux
    port map (
            O => \N__44224\,
            I => \N__44200\
        );

    \I__9706\ : LocalMux
    port map (
            O => \N__44221\,
            I => \N__44197\
        );

    \I__9705\ : LocalMux
    port map (
            O => \N__44218\,
            I => \N__44194\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__44215\,
            I => \N__44191\
        );

    \I__9703\ : Span4Mux_v
    port map (
            O => \N__44212\,
            I => \N__44184\
        );

    \I__9702\ : Span4Mux_v
    port map (
            O => \N__44209\,
            I => \N__44184\
        );

    \I__9701\ : Span4Mux_v
    port map (
            O => \N__44206\,
            I => \N__44184\
        );

    \I__9700\ : Span4Mux_h
    port map (
            O => \N__44203\,
            I => \N__44181\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__44200\,
            I => \N__44178\
        );

    \I__9698\ : Span4Mux_v
    port map (
            O => \N__44197\,
            I => \N__44175\
        );

    \I__9697\ : Span4Mux_v
    port map (
            O => \N__44194\,
            I => \N__44170\
        );

    \I__9696\ : Span4Mux_h
    port map (
            O => \N__44191\,
            I => \N__44170\
        );

    \I__9695\ : Span4Mux_h
    port map (
            O => \N__44184\,
            I => \N__44167\
        );

    \I__9694\ : Span4Mux_h
    port map (
            O => \N__44181\,
            I => \N__44164\
        );

    \I__9693\ : Span4Mux_v
    port map (
            O => \N__44178\,
            I => \N__44161\
        );

    \I__9692\ : Sp12to4
    port map (
            O => \N__44175\,
            I => \N__44158\
        );

    \I__9691\ : Span4Mux_h
    port map (
            O => \N__44170\,
            I => \N__44155\
        );

    \I__9690\ : Span4Mux_h
    port map (
            O => \N__44167\,
            I => \N__44152\
        );

    \I__9689\ : Span4Mux_h
    port map (
            O => \N__44164\,
            I => \N__44149\
        );

    \I__9688\ : Sp12to4
    port map (
            O => \N__44161\,
            I => \N__44144\
        );

    \I__9687\ : Span12Mux_h
    port map (
            O => \N__44158\,
            I => \N__44144\
        );

    \I__9686\ : Odrv4
    port map (
            O => \N__44155\,
            I => \sDAC_mem_3_1_sqmuxa\
        );

    \I__9685\ : Odrv4
    port map (
            O => \N__44152\,
            I => \sDAC_mem_3_1_sqmuxa\
        );

    \I__9684\ : Odrv4
    port map (
            O => \N__44149\,
            I => \sDAC_mem_3_1_sqmuxa\
        );

    \I__9683\ : Odrv12
    port map (
            O => \N__44144\,
            I => \sDAC_mem_3_1_sqmuxa\
        );

    \I__9682\ : InMux
    port map (
            O => \N__44135\,
            I => \N__44132\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__44132\,
            I => \N__44129\
        );

    \I__9680\ : Span4Mux_h
    port map (
            O => \N__44129\,
            I => \N__44126\
        );

    \I__9679\ : Odrv4
    port map (
            O => \N__44126\,
            I => \sDAC_mem_1Z0Z_0\
        );

    \I__9678\ : InMux
    port map (
            O => \N__44123\,
            I => \N__44120\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__44120\,
            I => \N__44117\
        );

    \I__9676\ : Span4Mux_v
    port map (
            O => \N__44117\,
            I => \N__44114\
        );

    \I__9675\ : Odrv4
    port map (
            O => \N__44114\,
            I => \sDAC_mem_1Z0Z_1\
        );

    \I__9674\ : InMux
    port map (
            O => \N__44111\,
            I => \N__44108\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__44108\,
            I => \N__44105\
        );

    \I__9672\ : Odrv4
    port map (
            O => \N__44105\,
            I => \sDAC_mem_1Z0Z_2\
        );

    \I__9671\ : InMux
    port map (
            O => \N__44102\,
            I => \N__44099\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__44099\,
            I => \N__44096\
        );

    \I__9669\ : Odrv4
    port map (
            O => \N__44096\,
            I => \sDAC_mem_1Z0Z_3\
        );

    \I__9668\ : InMux
    port map (
            O => \N__44093\,
            I => \N__44090\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__44090\,
            I => \N__44087\
        );

    \I__9666\ : Odrv4
    port map (
            O => \N__44087\,
            I => \sDAC_mem_1Z0Z_4\
        );

    \I__9665\ : InMux
    port map (
            O => \N__44084\,
            I => \N__44081\
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__44081\,
            I => \N__44078\
        );

    \I__9663\ : Odrv4
    port map (
            O => \N__44078\,
            I => \sDAC_mem_1Z0Z_5\
        );

    \I__9662\ : IoInMux
    port map (
            O => \N__44075\,
            I => \N__44072\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__44072\,
            I => \N__44069\
        );

    \I__9660\ : IoSpan4Mux
    port map (
            O => \N__44069\,
            I => \N__44066\
        );

    \I__9659\ : Span4Mux_s3_h
    port map (
            O => \N__44066\,
            I => \N__44063\
        );

    \I__9658\ : Span4Mux_v
    port map (
            O => \N__44063\,
            I => \N__44060\
        );

    \I__9657\ : Span4Mux_v
    port map (
            O => \N__44060\,
            I => \N__44057\
        );

    \I__9656\ : Sp12to4
    port map (
            O => \N__44057\,
            I => \N__44053\
        );

    \I__9655\ : InMux
    port map (
            O => \N__44056\,
            I => \N__44050\
        );

    \I__9654\ : Odrv12
    port map (
            O => \N__44053\,
            I => \RAM_DATA_cl_10Z0Z_15\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__44050\,
            I => \RAM_DATA_cl_10Z0Z_15\
        );

    \I__9652\ : IoInMux
    port map (
            O => \N__44045\,
            I => \N__44042\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__44042\,
            I => \N__44039\
        );

    \I__9650\ : Span4Mux_s0_v
    port map (
            O => \N__44039\,
            I => \N__44036\
        );

    \I__9649\ : Span4Mux_v
    port map (
            O => \N__44036\,
            I => \N__44033\
        );

    \I__9648\ : Span4Mux_v
    port map (
            O => \N__44033\,
            I => \N__44029\
        );

    \I__9647\ : CascadeMux
    port map (
            O => \N__44032\,
            I => \N__44026\
        );

    \I__9646\ : Sp12to4
    port map (
            O => \N__44029\,
            I => \N__44023\
        );

    \I__9645\ : InMux
    port map (
            O => \N__44026\,
            I => \N__44020\
        );

    \I__9644\ : Odrv12
    port map (
            O => \N__44023\,
            I => \RAM_DATA_cl_3Z0Z_15\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__44020\,
            I => \RAM_DATA_cl_3Z0Z_15\
        );

    \I__9642\ : IoInMux
    port map (
            O => \N__44015\,
            I => \N__44012\
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__44012\,
            I => \N__44009\
        );

    \I__9640\ : IoSpan4Mux
    port map (
            O => \N__44009\,
            I => \N__44006\
        );

    \I__9639\ : Span4Mux_s0_v
    port map (
            O => \N__44006\,
            I => \N__44003\
        );

    \I__9638\ : Span4Mux_v
    port map (
            O => \N__44003\,
            I => \N__44000\
        );

    \I__9637\ : Span4Mux_v
    port map (
            O => \N__44000\,
            I => \N__43996\
        );

    \I__9636\ : InMux
    port map (
            O => \N__43999\,
            I => \N__43993\
        );

    \I__9635\ : Odrv4
    port map (
            O => \N__43996\,
            I => \RAM_DATA_cl_4Z0Z_15\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__43993\,
            I => \RAM_DATA_cl_4Z0Z_15\
        );

    \I__9633\ : IoInMux
    port map (
            O => \N__43988\,
            I => \N__43985\
        );

    \I__9632\ : LocalMux
    port map (
            O => \N__43985\,
            I => \N__43982\
        );

    \I__9631\ : Span4Mux_s3_h
    port map (
            O => \N__43982\,
            I => \N__43979\
        );

    \I__9630\ : Span4Mux_v
    port map (
            O => \N__43979\,
            I => \N__43976\
        );

    \I__9629\ : Span4Mux_v
    port map (
            O => \N__43976\,
            I => \N__43972\
        );

    \I__9628\ : CascadeMux
    port map (
            O => \N__43975\,
            I => \N__43969\
        );

    \I__9627\ : Span4Mux_h
    port map (
            O => \N__43972\,
            I => \N__43966\
        );

    \I__9626\ : InMux
    port map (
            O => \N__43969\,
            I => \N__43963\
        );

    \I__9625\ : Odrv4
    port map (
            O => \N__43966\,
            I => \RAM_DATA_cl_2Z0Z_15\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__43963\,
            I => \RAM_DATA_cl_2Z0Z_15\
        );

    \I__9623\ : CEMux
    port map (
            O => \N__43958\,
            I => \N__43922\
        );

    \I__9622\ : CEMux
    port map (
            O => \N__43957\,
            I => \N__43922\
        );

    \I__9621\ : CEMux
    port map (
            O => \N__43956\,
            I => \N__43922\
        );

    \I__9620\ : CEMux
    port map (
            O => \N__43955\,
            I => \N__43922\
        );

    \I__9619\ : CEMux
    port map (
            O => \N__43954\,
            I => \N__43922\
        );

    \I__9618\ : CEMux
    port map (
            O => \N__43953\,
            I => \N__43922\
        );

    \I__9617\ : CEMux
    port map (
            O => \N__43952\,
            I => \N__43922\
        );

    \I__9616\ : CEMux
    port map (
            O => \N__43951\,
            I => \N__43922\
        );

    \I__9615\ : CEMux
    port map (
            O => \N__43950\,
            I => \N__43922\
        );

    \I__9614\ : CEMux
    port map (
            O => \N__43949\,
            I => \N__43922\
        );

    \I__9613\ : CEMux
    port map (
            O => \N__43948\,
            I => \N__43922\
        );

    \I__9612\ : CEMux
    port map (
            O => \N__43947\,
            I => \N__43922\
        );

    \I__9611\ : GlobalMux
    port map (
            O => \N__43922\,
            I => \N__43919\
        );

    \I__9610\ : gio2CtrlBuf
    port map (
            O => \N__43919\,
            I => op_eq_scounterdac10_g
        );

    \I__9609\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43913\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__43913\,
            I => \N__43910\
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__43910\,
            I => \sDAC_dataZ0Z_2\
        );

    \I__9606\ : CEMux
    port map (
            O => \N__43907\,
            I => \N__43904\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__43904\,
            I => \N__43898\
        );

    \I__9604\ : CEMux
    port map (
            O => \N__43903\,
            I => \N__43895\
        );

    \I__9603\ : CEMux
    port map (
            O => \N__43902\,
            I => \N__43892\
        );

    \I__9602\ : CEMux
    port map (
            O => \N__43901\,
            I => \N__43889\
        );

    \I__9601\ : Span4Mux_h
    port map (
            O => \N__43898\,
            I => \N__43883\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__43895\,
            I => \N__43883\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__43892\,
            I => \N__43880\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__43889\,
            I => \N__43877\
        );

    \I__9597\ : CascadeMux
    port map (
            O => \N__43888\,
            I => \N__43874\
        );

    \I__9596\ : Span4Mux_h
    port map (
            O => \N__43883\,
            I => \N__43871\
        );

    \I__9595\ : Span4Mux_h
    port map (
            O => \N__43880\,
            I => \N__43868\
        );

    \I__9594\ : Span4Mux_h
    port map (
            O => \N__43877\,
            I => \N__43865\
        );

    \I__9593\ : InMux
    port map (
            O => \N__43874\,
            I => \N__43862\
        );

    \I__9592\ : Odrv4
    port map (
            O => \N__43871\,
            I => \spi_master_inst.spi_data_path_u1.tx_ready_iZ0\
        );

    \I__9591\ : Odrv4
    port map (
            O => \N__43868\,
            I => \spi_master_inst.spi_data_path_u1.tx_ready_iZ0\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__43865\,
            I => \spi_master_inst.spi_data_path_u1.tx_ready_iZ0\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__43862\,
            I => \spi_master_inst.spi_data_path_u1.tx_ready_iZ0\
        );

    \I__9588\ : InMux
    port map (
            O => \N__43853\,
            I => \N__43850\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__43850\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_2\
        );

    \I__9586\ : InMux
    port map (
            O => \N__43847\,
            I => \N__43844\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__43844\,
            I => \N__43841\
        );

    \I__9584\ : Span12Mux_h
    port map (
            O => \N__43841\,
            I => \N__43838\
        );

    \I__9583\ : Odrv12
    port map (
            O => \N__43838\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2\
        );

    \I__9582\ : InMux
    port map (
            O => \N__43835\,
            I => \N__43832\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__43832\,
            I => \N__43829\
        );

    \I__9580\ : Span4Mux_h
    port map (
            O => \N__43829\,
            I => \N__43826\
        );

    \I__9579\ : Span4Mux_h
    port map (
            O => \N__43826\,
            I => \N__43823\
        );

    \I__9578\ : Odrv4
    port map (
            O => \N__43823\,
            I => \sDAC_mem_7Z0Z_2\
        );

    \I__9577\ : InMux
    port map (
            O => \N__43820\,
            I => \N__43817\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__43817\,
            I => \N__43814\
        );

    \I__9575\ : Span12Mux_v
    port map (
            O => \N__43814\,
            I => \N__43811\
        );

    \I__9574\ : Odrv12
    port map (
            O => \N__43811\,
            I => \sDAC_mem_7Z0Z_3\
        );

    \I__9573\ : InMux
    port map (
            O => \N__43808\,
            I => \N__43805\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__43805\,
            I => \N__43802\
        );

    \I__9571\ : Span4Mux_h
    port map (
            O => \N__43802\,
            I => \N__43799\
        );

    \I__9570\ : Span4Mux_v
    port map (
            O => \N__43799\,
            I => \N__43796\
        );

    \I__9569\ : Span4Mux_v
    port map (
            O => \N__43796\,
            I => \N__43793\
        );

    \I__9568\ : IoSpan4Mux
    port map (
            O => \N__43793\,
            I => \N__43790\
        );

    \I__9567\ : Odrv4
    port map (
            O => \N__43790\,
            I => \RAM_DATA_in_1\
        );

    \I__9566\ : InMux
    port map (
            O => \N__43787\,
            I => \N__43784\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__43784\,
            I => \N__43781\
        );

    \I__9564\ : Span12Mux_h
    port map (
            O => \N__43781\,
            I => \N__43778\
        );

    \I__9563\ : Span12Mux_v
    port map (
            O => \N__43778\,
            I => \N__43775\
        );

    \I__9562\ : Odrv12
    port map (
            O => \N__43775\,
            I => \RAM_DATA_in_9\
        );

    \I__9561\ : CascadeMux
    port map (
            O => \N__43772\,
            I => \N__43762\
        );

    \I__9560\ : CascadeMux
    port map (
            O => \N__43771\,
            I => \N__43759\
        );

    \I__9559\ : CascadeMux
    port map (
            O => \N__43770\,
            I => \N__43756\
        );

    \I__9558\ : InMux
    port map (
            O => \N__43769\,
            I => \N__43751\
        );

    \I__9557\ : InMux
    port map (
            O => \N__43768\,
            I => \N__43751\
        );

    \I__9556\ : InMux
    port map (
            O => \N__43767\,
            I => \N__43748\
        );

    \I__9555\ : InMux
    port map (
            O => \N__43766\,
            I => \N__43737\
        );

    \I__9554\ : InMux
    port map (
            O => \N__43765\,
            I => \N__43737\
        );

    \I__9553\ : InMux
    port map (
            O => \N__43762\,
            I => \N__43737\
        );

    \I__9552\ : InMux
    port map (
            O => \N__43759\,
            I => \N__43737\
        );

    \I__9551\ : InMux
    port map (
            O => \N__43756\,
            I => \N__43737\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__43751\,
            I => \N__43732\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__43748\,
            I => \N__43729\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__43737\,
            I => \N__43726\
        );

    \I__9547\ : InMux
    port map (
            O => \N__43736\,
            I => \N__43723\
        );

    \I__9546\ : InMux
    port map (
            O => \N__43735\,
            I => \N__43720\
        );

    \I__9545\ : Span4Mux_h
    port map (
            O => \N__43732\,
            I => \N__43717\
        );

    \I__9544\ : Span4Mux_h
    port map (
            O => \N__43729\,
            I => \N__43714\
        );

    \I__9543\ : Span4Mux_v
    port map (
            O => \N__43726\,
            I => \N__43709\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__43723\,
            I => \N__43709\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__43720\,
            I => \N_75\
        );

    \I__9540\ : Odrv4
    port map (
            O => \N__43717\,
            I => \N_75\
        );

    \I__9539\ : Odrv4
    port map (
            O => \N__43714\,
            I => \N_75\
        );

    \I__9538\ : Odrv4
    port map (
            O => \N__43709\,
            I => \N_75\
        );

    \I__9537\ : InMux
    port map (
            O => \N__43700\,
            I => \N__43697\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__43697\,
            I => \N__43694\
        );

    \I__9535\ : Odrv4
    port map (
            O => \N__43694\,
            I => \spi_data_misoZ0Z_1\
        );

    \I__9534\ : CEMux
    port map (
            O => \N__43691\,
            I => \N__43688\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__43688\,
            I => \N__43683\
        );

    \I__9532\ : CEMux
    port map (
            O => \N__43687\,
            I => \N__43680\
        );

    \I__9531\ : CEMux
    port map (
            O => \N__43686\,
            I => \N__43677\
        );

    \I__9530\ : Span4Mux_v
    port map (
            O => \N__43683\,
            I => \N__43674\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__43680\,
            I => \N__43671\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__43677\,
            I => \N__43668\
        );

    \I__9527\ : Odrv4
    port map (
            O => \N__43674\,
            I => \sSPI_MSB0LSB1_RNIGRPGZ0Z4\
        );

    \I__9526\ : Odrv4
    port map (
            O => \N__43671\,
            I => \sSPI_MSB0LSB1_RNIGRPGZ0Z4\
        );

    \I__9525\ : Odrv12
    port map (
            O => \N__43668\,
            I => \sSPI_MSB0LSB1_RNIGRPGZ0Z4\
        );

    \I__9524\ : InMux
    port map (
            O => \N__43661\,
            I => \N__43658\
        );

    \I__9523\ : LocalMux
    port map (
            O => \N__43658\,
            I => \N__43655\
        );

    \I__9522\ : Span4Mux_v
    port map (
            O => \N__43655\,
            I => \N__43652\
        );

    \I__9521\ : Span4Mux_h
    port map (
            O => \N__43652\,
            I => \N__43649\
        );

    \I__9520\ : Sp12to4
    port map (
            O => \N__43649\,
            I => \N__43646\
        );

    \I__9519\ : Span12Mux_h
    port map (
            O => \N__43646\,
            I => \N__43642\
        );

    \I__9518\ : InMux
    port map (
            O => \N__43645\,
            I => \N__43639\
        );

    \I__9517\ : Odrv12
    port map (
            O => \N__43642\,
            I => \sRAM_pointer_writeZ0Z_8\
        );

    \I__9516\ : LocalMux
    port map (
            O => \N__43639\,
            I => \sRAM_pointer_writeZ0Z_8\
        );

    \I__9515\ : CascadeMux
    port map (
            O => \N__43634\,
            I => \N__43631\
        );

    \I__9514\ : InMux
    port map (
            O => \N__43631\,
            I => \N__43628\
        );

    \I__9513\ : LocalMux
    port map (
            O => \N__43628\,
            I => \N__43625\
        );

    \I__9512\ : Span4Mux_h
    port map (
            O => \N__43625\,
            I => \N__43622\
        );

    \I__9511\ : Span4Mux_h
    port map (
            O => \N__43622\,
            I => \N__43618\
        );

    \I__9510\ : InMux
    port map (
            O => \N__43621\,
            I => \N__43615\
        );

    \I__9509\ : Odrv4
    port map (
            O => \N__43618\,
            I => \sRAM_pointer_readZ0Z_8\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__43615\,
            I => \sRAM_pointer_readZ0Z_8\
        );

    \I__9507\ : IoInMux
    port map (
            O => \N__43610\,
            I => \N__43607\
        );

    \I__9506\ : LocalMux
    port map (
            O => \N__43607\,
            I => \N__43604\
        );

    \I__9505\ : IoSpan4Mux
    port map (
            O => \N__43604\,
            I => \N__43601\
        );

    \I__9504\ : Span4Mux_s3_h
    port map (
            O => \N__43601\,
            I => \N__43598\
        );

    \I__9503\ : Span4Mux_h
    port map (
            O => \N__43598\,
            I => \N__43595\
        );

    \I__9502\ : Span4Mux_v
    port map (
            O => \N__43595\,
            I => \N__43592\
        );

    \I__9501\ : Odrv4
    port map (
            O => \N__43592\,
            I => \RAM_ADD_c_8\
        );

    \I__9500\ : InMux
    port map (
            O => \N__43589\,
            I => \N__43586\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__43586\,
            I => \N__43583\
        );

    \I__9498\ : Span4Mux_h
    port map (
            O => \N__43583\,
            I => \N__43580\
        );

    \I__9497\ : Span4Mux_h
    port map (
            O => \N__43580\,
            I => \N__43577\
        );

    \I__9496\ : Sp12to4
    port map (
            O => \N__43577\,
            I => \N__43574\
        );

    \I__9495\ : Span12Mux_v
    port map (
            O => \N__43574\,
            I => \N__43570\
        );

    \I__9494\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43567\
        );

    \I__9493\ : Odrv12
    port map (
            O => \N__43570\,
            I => \sRAM_pointer_writeZ0Z_4\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__43567\,
            I => \sRAM_pointer_writeZ0Z_4\
        );

    \I__9491\ : CascadeMux
    port map (
            O => \N__43562\,
            I => \N__43559\
        );

    \I__9490\ : InMux
    port map (
            O => \N__43559\,
            I => \N__43556\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__43556\,
            I => \N__43553\
        );

    \I__9488\ : Span4Mux_h
    port map (
            O => \N__43553\,
            I => \N__43550\
        );

    \I__9487\ : Span4Mux_h
    port map (
            O => \N__43550\,
            I => \N__43546\
        );

    \I__9486\ : InMux
    port map (
            O => \N__43549\,
            I => \N__43543\
        );

    \I__9485\ : Odrv4
    port map (
            O => \N__43546\,
            I => \sRAM_pointer_readZ0Z_4\
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__43543\,
            I => \sRAM_pointer_readZ0Z_4\
        );

    \I__9483\ : IoInMux
    port map (
            O => \N__43538\,
            I => \N__43535\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__43535\,
            I => \N__43532\
        );

    \I__9481\ : Span4Mux_s2_v
    port map (
            O => \N__43532\,
            I => \N__43529\
        );

    \I__9480\ : Span4Mux_h
    port map (
            O => \N__43529\,
            I => \N__43526\
        );

    \I__9479\ : Span4Mux_v
    port map (
            O => \N__43526\,
            I => \N__43523\
        );

    \I__9478\ : Odrv4
    port map (
            O => \N__43523\,
            I => \RAM_ADD_c_4\
        );

    \I__9477\ : InMux
    port map (
            O => \N__43520\,
            I => \N__43517\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__43517\,
            I => \N__43514\
        );

    \I__9475\ : Span12Mux_v
    port map (
            O => \N__43514\,
            I => \N__43511\
        );

    \I__9474\ : Span12Mux_h
    port map (
            O => \N__43511\,
            I => \N__43507\
        );

    \I__9473\ : InMux
    port map (
            O => \N__43510\,
            I => \N__43504\
        );

    \I__9472\ : Odrv12
    port map (
            O => \N__43507\,
            I => \sRAM_pointer_writeZ0Z_3\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__43504\,
            I => \sRAM_pointer_writeZ0Z_3\
        );

    \I__9470\ : InMux
    port map (
            O => \N__43499\,
            I => \N__43478\
        );

    \I__9469\ : InMux
    port map (
            O => \N__43498\,
            I => \N__43478\
        );

    \I__9468\ : InMux
    port map (
            O => \N__43497\,
            I => \N__43478\
        );

    \I__9467\ : InMux
    port map (
            O => \N__43496\,
            I => \N__43478\
        );

    \I__9466\ : InMux
    port map (
            O => \N__43495\,
            I => \N__43469\
        );

    \I__9465\ : InMux
    port map (
            O => \N__43494\,
            I => \N__43469\
        );

    \I__9464\ : InMux
    port map (
            O => \N__43493\,
            I => \N__43469\
        );

    \I__9463\ : InMux
    port map (
            O => \N__43492\,
            I => \N__43469\
        );

    \I__9462\ : CascadeMux
    port map (
            O => \N__43491\,
            I => \N__43463\
        );

    \I__9461\ : CascadeMux
    port map (
            O => \N__43490\,
            I => \N__43459\
        );

    \I__9460\ : CascadeMux
    port map (
            O => \N__43489\,
            I => \N__43455\
        );

    \I__9459\ : CascadeMux
    port map (
            O => \N__43488\,
            I => \N__43451\
        );

    \I__9458\ : CascadeMux
    port map (
            O => \N__43487\,
            I => \N__43447\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__43478\,
            I => \N__43440\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__43469\,
            I => \N__43440\
        );

    \I__9455\ : InMux
    port map (
            O => \N__43468\,
            I => \N__43433\
        );

    \I__9454\ : InMux
    port map (
            O => \N__43467\,
            I => \N__43433\
        );

    \I__9453\ : InMux
    port map (
            O => \N__43466\,
            I => \N__43430\
        );

    \I__9452\ : InMux
    port map (
            O => \N__43463\,
            I => \N__43413\
        );

    \I__9451\ : InMux
    port map (
            O => \N__43462\,
            I => \N__43413\
        );

    \I__9450\ : InMux
    port map (
            O => \N__43459\,
            I => \N__43413\
        );

    \I__9449\ : InMux
    port map (
            O => \N__43458\,
            I => \N__43413\
        );

    \I__9448\ : InMux
    port map (
            O => \N__43455\,
            I => \N__43413\
        );

    \I__9447\ : InMux
    port map (
            O => \N__43454\,
            I => \N__43413\
        );

    \I__9446\ : InMux
    port map (
            O => \N__43451\,
            I => \N__43413\
        );

    \I__9445\ : InMux
    port map (
            O => \N__43450\,
            I => \N__43413\
        );

    \I__9444\ : InMux
    port map (
            O => \N__43447\,
            I => \N__43408\
        );

    \I__9443\ : InMux
    port map (
            O => \N__43446\,
            I => \N__43408\
        );

    \I__9442\ : InMux
    port map (
            O => \N__43445\,
            I => \N__43405\
        );

    \I__9441\ : Span4Mux_h
    port map (
            O => \N__43440\,
            I => \N__43402\
        );

    \I__9440\ : InMux
    port map (
            O => \N__43439\,
            I => \N__43399\
        );

    \I__9439\ : InMux
    port map (
            O => \N__43438\,
            I => \N__43396\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__43433\,
            I => \N__43385\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__43430\,
            I => \N__43385\
        );

    \I__9436\ : LocalMux
    port map (
            O => \N__43413\,
            I => \N__43385\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__43408\,
            I => \N__43385\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__43405\,
            I => \N__43385\
        );

    \I__9433\ : Odrv4
    port map (
            O => \N__43402\,
            I => \un1_sacqtime_cry_23_THRU_CO\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__43399\,
            I => \un1_sacqtime_cry_23_THRU_CO\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__43396\,
            I => \un1_sacqtime_cry_23_THRU_CO\
        );

    \I__9430\ : Odrv12
    port map (
            O => \N__43385\,
            I => \un1_sacqtime_cry_23_THRU_CO\
        );

    \I__9429\ : CascadeMux
    port map (
            O => \N__43376\,
            I => \N__43373\
        );

    \I__9428\ : InMux
    port map (
            O => \N__43373\,
            I => \N__43370\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__43370\,
            I => \N__43367\
        );

    \I__9426\ : Span12Mux_h
    port map (
            O => \N__43367\,
            I => \N__43363\
        );

    \I__9425\ : InMux
    port map (
            O => \N__43366\,
            I => \N__43360\
        );

    \I__9424\ : Odrv12
    port map (
            O => \N__43363\,
            I => \sRAM_pointer_readZ0Z_3\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__43360\,
            I => \sRAM_pointer_readZ0Z_3\
        );

    \I__9422\ : InMux
    port map (
            O => \N__43355\,
            I => \N__43317\
        );

    \I__9421\ : InMux
    port map (
            O => \N__43354\,
            I => \N__43317\
        );

    \I__9420\ : InMux
    port map (
            O => \N__43353\,
            I => \N__43317\
        );

    \I__9419\ : InMux
    port map (
            O => \N__43352\,
            I => \N__43317\
        );

    \I__9418\ : InMux
    port map (
            O => \N__43351\,
            I => \N__43317\
        );

    \I__9417\ : InMux
    port map (
            O => \N__43350\,
            I => \N__43317\
        );

    \I__9416\ : InMux
    port map (
            O => \N__43349\,
            I => \N__43317\
        );

    \I__9415\ : InMux
    port map (
            O => \N__43348\,
            I => \N__43317\
        );

    \I__9414\ : InMux
    port map (
            O => \N__43347\,
            I => \N__43308\
        );

    \I__9413\ : InMux
    port map (
            O => \N__43346\,
            I => \N__43308\
        );

    \I__9412\ : InMux
    port map (
            O => \N__43345\,
            I => \N__43308\
        );

    \I__9411\ : InMux
    port map (
            O => \N__43344\,
            I => \N__43291\
        );

    \I__9410\ : InMux
    port map (
            O => \N__43343\,
            I => \N__43291\
        );

    \I__9409\ : InMux
    port map (
            O => \N__43342\,
            I => \N__43291\
        );

    \I__9408\ : InMux
    port map (
            O => \N__43341\,
            I => \N__43291\
        );

    \I__9407\ : InMux
    port map (
            O => \N__43340\,
            I => \N__43291\
        );

    \I__9406\ : InMux
    port map (
            O => \N__43339\,
            I => \N__43291\
        );

    \I__9405\ : InMux
    port map (
            O => \N__43338\,
            I => \N__43291\
        );

    \I__9404\ : InMux
    port map (
            O => \N__43337\,
            I => \N__43291\
        );

    \I__9403\ : InMux
    port map (
            O => \N__43336\,
            I => \N__43286\
        );

    \I__9402\ : InMux
    port map (
            O => \N__43335\,
            I => \N__43286\
        );

    \I__9401\ : InMux
    port map (
            O => \N__43334\,
            I => \N__43283\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__43317\,
            I => \N__43280\
        );

    \I__9399\ : InMux
    port map (
            O => \N__43316\,
            I => \N__43277\
        );

    \I__9398\ : InMux
    port map (
            O => \N__43315\,
            I => \N__43274\
        );

    \I__9397\ : LocalMux
    port map (
            O => \N__43308\,
            I => \N__43265\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__43291\,
            I => \N__43265\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__43286\,
            I => \N__43265\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__43283\,
            I => \N__43265\
        );

    \I__9393\ : Span4Mux_h
    port map (
            O => \N__43280\,
            I => \N__43262\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__43277\,
            I => \N__43255\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__43274\,
            I => \N__43255\
        );

    \I__9390\ : Span4Mux_h
    port map (
            O => \N__43265\,
            I => \N__43255\
        );

    \I__9389\ : Span4Mux_h
    port map (
            O => \N__43262\,
            I => \N__43252\
        );

    \I__9388\ : Span4Mux_h
    port map (
            O => \N__43255\,
            I => \N__43249\
        );

    \I__9387\ : Odrv4
    port map (
            O => \N__43252\,
            I => \un4_sacqtime_cry_23_THRU_CO\
        );

    \I__9386\ : Odrv4
    port map (
            O => \N__43249\,
            I => \un4_sacqtime_cry_23_THRU_CO\
        );

    \I__9385\ : IoInMux
    port map (
            O => \N__43244\,
            I => \N__43241\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__43241\,
            I => \N__43238\
        );

    \I__9383\ : Span4Mux_s1_v
    port map (
            O => \N__43238\,
            I => \N__43235\
        );

    \I__9382\ : Span4Mux_v
    port map (
            O => \N__43235\,
            I => \N__43232\
        );

    \I__9381\ : Span4Mux_v
    port map (
            O => \N__43232\,
            I => \N__43229\
        );

    \I__9380\ : Odrv4
    port map (
            O => \N__43229\,
            I => \RAM_ADD_c_3\
        );

    \I__9379\ : CEMux
    port map (
            O => \N__43226\,
            I => \N__43222\
        );

    \I__9378\ : CEMux
    port map (
            O => \N__43225\,
            I => \N__43219\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__43222\,
            I => \N__43215\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__43219\,
            I => \N__43212\
        );

    \I__9375\ : CEMux
    port map (
            O => \N__43218\,
            I => \N__43209\
        );

    \I__9374\ : Span4Mux_v
    port map (
            O => \N__43215\,
            I => \N__43206\
        );

    \I__9373\ : Span4Mux_h
    port map (
            O => \N__43212\,
            I => \N__43203\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__43209\,
            I => \N__43200\
        );

    \I__9371\ : Span4Mux_h
    port map (
            O => \N__43206\,
            I => \N__43193\
        );

    \I__9370\ : Span4Mux_h
    port map (
            O => \N__43203\,
            I => \N__43193\
        );

    \I__9369\ : Span4Mux_v
    port map (
            O => \N__43200\,
            I => \N__43193\
        );

    \I__9368\ : Odrv4
    port map (
            O => \N__43193\,
            I => \N_67_i\
        );

    \I__9367\ : IoInMux
    port map (
            O => \N__43190\,
            I => \N__43187\
        );

    \I__9366\ : LocalMux
    port map (
            O => \N__43187\,
            I => \N__43184\
        );

    \I__9365\ : Span12Mux_s8_v
    port map (
            O => \N__43184\,
            I => \N__43180\
        );

    \I__9364\ : InMux
    port map (
            O => \N__43183\,
            I => \N__43177\
        );

    \I__9363\ : Odrv12
    port map (
            O => \N__43180\,
            I => \RAM_DATA_cl_13Z0Z_15\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__43177\,
            I => \RAM_DATA_cl_13Z0Z_15\
        );

    \I__9361\ : IoInMux
    port map (
            O => \N__43172\,
            I => \N__43169\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__43169\,
            I => \N__43166\
        );

    \I__9359\ : Span4Mux_s2_v
    port map (
            O => \N__43166\,
            I => \N__43163\
        );

    \I__9358\ : Span4Mux_h
    port map (
            O => \N__43163\,
            I => \N__43160\
        );

    \I__9357\ : Span4Mux_h
    port map (
            O => \N__43160\,
            I => \N__43156\
        );

    \I__9356\ : CascadeMux
    port map (
            O => \N__43159\,
            I => \N__43153\
        );

    \I__9355\ : Span4Mux_v
    port map (
            O => \N__43156\,
            I => \N__43150\
        );

    \I__9354\ : InMux
    port map (
            O => \N__43153\,
            I => \N__43147\
        );

    \I__9353\ : Odrv4
    port map (
            O => \N__43150\,
            I => \RAM_DATA_cl_14Z0Z_15\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__43147\,
            I => \RAM_DATA_cl_14Z0Z_15\
        );

    \I__9351\ : IoInMux
    port map (
            O => \N__43142\,
            I => \N__43139\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__43139\,
            I => \N__43136\
        );

    \I__9349\ : Span4Mux_s3_h
    port map (
            O => \N__43136\,
            I => \N__43133\
        );

    \I__9348\ : Span4Mux_v
    port map (
            O => \N__43133\,
            I => \N__43130\
        );

    \I__9347\ : Span4Mux_v
    port map (
            O => \N__43130\,
            I => \N__43127\
        );

    \I__9346\ : Span4Mux_h
    port map (
            O => \N__43127\,
            I => \N__43123\
        );

    \I__9345\ : InMux
    port map (
            O => \N__43126\,
            I => \N__43120\
        );

    \I__9344\ : Odrv4
    port map (
            O => \N__43123\,
            I => \RAM_DATA_cl_15Z0Z_15\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__43120\,
            I => \RAM_DATA_cl_15Z0Z_15\
        );

    \I__9342\ : IoInMux
    port map (
            O => \N__43115\,
            I => \N__43112\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__43112\,
            I => \N__43109\
        );

    \I__9340\ : IoSpan4Mux
    port map (
            O => \N__43109\,
            I => \N__43106\
        );

    \I__9339\ : Span4Mux_s2_h
    port map (
            O => \N__43106\,
            I => \N__43103\
        );

    \I__9338\ : Sp12to4
    port map (
            O => \N__43103\,
            I => \N__43100\
        );

    \I__9337\ : Span12Mux_s10_h
    port map (
            O => \N__43100\,
            I => \N__43096\
        );

    \I__9336\ : CascadeMux
    port map (
            O => \N__43099\,
            I => \N__43093\
        );

    \I__9335\ : Span12Mux_v
    port map (
            O => \N__43096\,
            I => \N__43090\
        );

    \I__9334\ : InMux
    port map (
            O => \N__43093\,
            I => \N__43087\
        );

    \I__9333\ : Odrv12
    port map (
            O => \N__43090\,
            I => \RAM_DATA_cl_1Z0Z_15\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__43087\,
            I => \RAM_DATA_cl_1Z0Z_15\
        );

    \I__9331\ : InMux
    port map (
            O => \N__43082\,
            I => \sCounterADC_cry_2\
        );

    \I__9330\ : InMux
    port map (
            O => \N__43079\,
            I => \N__43076\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__43076\,
            I => \N__43073\
        );

    \I__9328\ : Span4Mux_v
    port map (
            O => \N__43073\,
            I => \N__43070\
        );

    \I__9327\ : Span4Mux_h
    port map (
            O => \N__43070\,
            I => \N__43066\
        );

    \I__9326\ : InMux
    port map (
            O => \N__43069\,
            I => \N__43063\
        );

    \I__9325\ : Span4Mux_h
    port map (
            O => \N__43066\,
            I => \N__43060\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__43063\,
            I => \sCounterADCZ0Z_4\
        );

    \I__9323\ : Odrv4
    port map (
            O => \N__43060\,
            I => \sCounterADCZ0Z_4\
        );

    \I__9322\ : InMux
    port map (
            O => \N__43055\,
            I => \sCounterADC_cry_3\
        );

    \I__9321\ : InMux
    port map (
            O => \N__43052\,
            I => \N__43049\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__43049\,
            I => \N__43046\
        );

    \I__9319\ : Span4Mux_v
    port map (
            O => \N__43046\,
            I => \N__43043\
        );

    \I__9318\ : Span4Mux_h
    port map (
            O => \N__43043\,
            I => \N__43039\
        );

    \I__9317\ : InMux
    port map (
            O => \N__43042\,
            I => \N__43036\
        );

    \I__9316\ : Span4Mux_h
    port map (
            O => \N__43039\,
            I => \N__43033\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__43036\,
            I => \sCounterADCZ0Z_5\
        );

    \I__9314\ : Odrv4
    port map (
            O => \N__43033\,
            I => \sCounterADCZ0Z_5\
        );

    \I__9313\ : InMux
    port map (
            O => \N__43028\,
            I => \sCounterADC_cry_4\
        );

    \I__9312\ : InMux
    port map (
            O => \N__43025\,
            I => \sCounterADC_cry_5\
        );

    \I__9311\ : InMux
    port map (
            O => \N__43022\,
            I => \sCounterADC_cry_6\
        );

    \I__9310\ : InMux
    port map (
            O => \N__43019\,
            I => \N__43016\
        );

    \I__9309\ : LocalMux
    port map (
            O => \N__43016\,
            I => \N__43013\
        );

    \I__9308\ : Span4Mux_v
    port map (
            O => \N__43013\,
            I => \N__43010\
        );

    \I__9307\ : Sp12to4
    port map (
            O => \N__43010\,
            I => \N__43007\
        );

    \I__9306\ : Span12Mux_h
    port map (
            O => \N__43007\,
            I => \N__43004\
        );

    \I__9305\ : Odrv12
    port map (
            O => \N__43004\,
            I => \RAM_DATA_in_5\
        );

    \I__9304\ : InMux
    port map (
            O => \N__43001\,
            I => \N__42998\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__42998\,
            I => \N__42995\
        );

    \I__9302\ : Span12Mux_v
    port map (
            O => \N__42995\,
            I => \N__42992\
        );

    \I__9301\ : Odrv12
    port map (
            O => \N__42992\,
            I => \RAM_DATA_in_13\
        );

    \I__9300\ : InMux
    port map (
            O => \N__42989\,
            I => \N__42986\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__42986\,
            I => \N__42983\
        );

    \I__9298\ : Odrv4
    port map (
            O => \N__42983\,
            I => \spi_data_misoZ0Z_5\
        );

    \I__9297\ : InMux
    port map (
            O => \N__42980\,
            I => \N__42977\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__42977\,
            I => \N__42974\
        );

    \I__9295\ : Span12Mux_v
    port map (
            O => \N__42974\,
            I => \N__42971\
        );

    \I__9294\ : Odrv12
    port map (
            O => \N__42971\,
            I => \RAM_DATA_in_15\
        );

    \I__9293\ : CascadeMux
    port map (
            O => \N__42968\,
            I => \N__42965\
        );

    \I__9292\ : InMux
    port map (
            O => \N__42965\,
            I => \N__42962\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__42962\,
            I => \N__42959\
        );

    \I__9290\ : Span4Mux_v
    port map (
            O => \N__42959\,
            I => \N__42956\
        );

    \I__9289\ : Span4Mux_v
    port map (
            O => \N__42956\,
            I => \N__42953\
        );

    \I__9288\ : Span4Mux_h
    port map (
            O => \N__42953\,
            I => \N__42950\
        );

    \I__9287\ : Span4Mux_h
    port map (
            O => \N__42950\,
            I => \N__42947\
        );

    \I__9286\ : Odrv4
    port map (
            O => \N__42947\,
            I => \RAM_DATA_in_7\
        );

    \I__9285\ : InMux
    port map (
            O => \N__42944\,
            I => \N__42941\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__42941\,
            I => \N__42938\
        );

    \I__9283\ : Odrv4
    port map (
            O => \N__42938\,
            I => \spi_data_misoZ0Z_7\
        );

    \I__9282\ : InMux
    port map (
            O => \N__42935\,
            I => \N__42932\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__42932\,
            I => \N__42929\
        );

    \I__9280\ : Span4Mux_v
    port map (
            O => \N__42929\,
            I => \N__42926\
        );

    \I__9279\ : Sp12to4
    port map (
            O => \N__42926\,
            I => \N__42923\
        );

    \I__9278\ : Span12Mux_h
    port map (
            O => \N__42923\,
            I => \N__42920\
        );

    \I__9277\ : Odrv12
    port map (
            O => \N__42920\,
            I => \RAM_DATA_in_3\
        );

    \I__9276\ : CascadeMux
    port map (
            O => \N__42917\,
            I => \N__42914\
        );

    \I__9275\ : InMux
    port map (
            O => \N__42914\,
            I => \N__42911\
        );

    \I__9274\ : LocalMux
    port map (
            O => \N__42911\,
            I => \N__42908\
        );

    \I__9273\ : Span4Mux_h
    port map (
            O => \N__42908\,
            I => \N__42905\
        );

    \I__9272\ : Sp12to4
    port map (
            O => \N__42905\,
            I => \N__42902\
        );

    \I__9271\ : Span12Mux_v
    port map (
            O => \N__42902\,
            I => \N__42899\
        );

    \I__9270\ : Odrv12
    port map (
            O => \N__42899\,
            I => \RAM_DATA_in_11\
        );

    \I__9269\ : InMux
    port map (
            O => \N__42896\,
            I => \N__42893\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__42893\,
            I => \N__42890\
        );

    \I__9267\ : Odrv4
    port map (
            O => \N__42890\,
            I => \spi_data_misoZ0Z_3\
        );

    \I__9266\ : InMux
    port map (
            O => \N__42887\,
            I => \N__42884\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__42884\,
            I => \N__42881\
        );

    \I__9264\ : Span12Mux_v
    port map (
            O => \N__42881\,
            I => \N__42878\
        );

    \I__9263\ : Span12Mux_v
    port map (
            O => \N__42878\,
            I => \N__42875\
        );

    \I__9262\ : Odrv12
    port map (
            O => \N__42875\,
            I => \RAM_DATA_in_10\
        );

    \I__9261\ : InMux
    port map (
            O => \N__42872\,
            I => \N__42869\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__42869\,
            I => \N__42866\
        );

    \I__9259\ : Span4Mux_v
    port map (
            O => \N__42866\,
            I => \N__42863\
        );

    \I__9258\ : Sp12to4
    port map (
            O => \N__42863\,
            I => \N__42860\
        );

    \I__9257\ : Span12Mux_h
    port map (
            O => \N__42860\,
            I => \N__42857\
        );

    \I__9256\ : Odrv12
    port map (
            O => \N__42857\,
            I => \RAM_DATA_in_2\
        );

    \I__9255\ : InMux
    port map (
            O => \N__42854\,
            I => \N__42851\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__42851\,
            I => \N__42848\
        );

    \I__9253\ : Odrv4
    port map (
            O => \N__42848\,
            I => \spi_data_misoZ0Z_2\
        );

    \I__9252\ : InMux
    port map (
            O => \N__42845\,
            I => \N__42842\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__42842\,
            I => \N__42839\
        );

    \I__9250\ : Odrv4
    port map (
            O => \N__42839\,
            I => \spi_data_misoZ0Z_4\
        );

    \I__9249\ : InMux
    port map (
            O => \N__42836\,
            I => \N__42833\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__42833\,
            I => \spi_data_misoZ0Z_6\
        );

    \I__9247\ : CEMux
    port map (
            O => \N__42830\,
            I => \N__42827\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__42827\,
            I => \N__42824\
        );

    \I__9245\ : Span4Mux_v
    port map (
            O => \N__42824\,
            I => \N__42821\
        );

    \I__9244\ : Span4Mux_v
    port map (
            O => \N__42821\,
            I => \N__42818\
        );

    \I__9243\ : Sp12to4
    port map (
            O => \N__42818\,
            I => \N__42815\
        );

    \I__9242\ : Odrv12
    port map (
            O => \N__42815\,
            I => \spi_slave_inst.un4_i_wr\
        );

    \I__9241\ : InMux
    port map (
            O => \N__42812\,
            I => \bfn_18_15_0_\
        );

    \I__9240\ : InMux
    port map (
            O => \N__42809\,
            I => \sCounterADC_cry_0\
        );

    \I__9239\ : InMux
    port map (
            O => \N__42806\,
            I => \sCounterADC_cry_1\
        );

    \I__9238\ : InMux
    port map (
            O => \N__42803\,
            I => \N__42800\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__42800\,
            I => \N__42797\
        );

    \I__9236\ : Span4Mux_h
    port map (
            O => \N__42797\,
            I => \N__42794\
        );

    \I__9235\ : Odrv4
    port map (
            O => \N__42794\,
            I => \sDAC_mem_25Z0Z_7\
        );

    \I__9234\ : CascadeMux
    port map (
            O => \N__42791\,
            I => \N__42788\
        );

    \I__9233\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42784\
        );

    \I__9232\ : InMux
    port map (
            O => \N__42787\,
            I => \N__42781\
        );

    \I__9231\ : LocalMux
    port map (
            O => \N__42784\,
            I => \N__42776\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__42781\,
            I => \N__42776\
        );

    \I__9229\ : Odrv12
    port map (
            O => \N__42776\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa\
        );

    \I__9228\ : InMux
    port map (
            O => \N__42773\,
            I => \N__42769\
        );

    \I__9227\ : CascadeMux
    port map (
            O => \N__42772\,
            I => \N__42765\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__42769\,
            I => \N__42762\
        );

    \I__9225\ : InMux
    port map (
            O => \N__42768\,
            I => \N__42759\
        );

    \I__9224\ : InMux
    port map (
            O => \N__42765\,
            I => \N__42756\
        );

    \I__9223\ : Span12Mux_h
    port map (
            O => \N__42762\,
            I => \N__42753\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__42759\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__42756\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0\
        );

    \I__9220\ : Odrv12
    port map (
            O => \N__42753\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0\
        );

    \I__9219\ : InMux
    port map (
            O => \N__42746\,
            I => \N__42743\
        );

    \I__9218\ : LocalMux
    port map (
            O => \N__42743\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO\
        );

    \I__9217\ : CascadeMux
    port map (
            O => \N__42740\,
            I => \N__42737\
        );

    \I__9216\ : InMux
    port map (
            O => \N__42737\,
            I => \N__42733\
        );

    \I__9215\ : CascadeMux
    port map (
            O => \N__42736\,
            I => \N__42730\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__42733\,
            I => \N__42726\
        );

    \I__9213\ : InMux
    port map (
            O => \N__42730\,
            I => \N__42723\
        );

    \I__9212\ : InMux
    port map (
            O => \N__42729\,
            I => \N__42720\
        );

    \I__9211\ : Span12Mux_h
    port map (
            O => \N__42726\,
            I => \N__42717\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__42723\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1\
        );

    \I__9209\ : LocalMux
    port map (
            O => \N__42720\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1\
        );

    \I__9208\ : Odrv12
    port map (
            O => \N__42717\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1\
        );

    \I__9207\ : CascadeMux
    port map (
            O => \N__42710\,
            I => \N__42707\
        );

    \I__9206\ : InMux
    port map (
            O => \N__42707\,
            I => \N__42702\
        );

    \I__9205\ : InMux
    port map (
            O => \N__42706\,
            I => \N__42697\
        );

    \I__9204\ : InMux
    port map (
            O => \N__42705\,
            I => \N__42697\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__42702\,
            I => \N__42692\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__42697\,
            I => \N__42692\
        );

    \I__9201\ : Odrv12
    port map (
            O => \N__42692\,
            I => \spi_slave_inst.un23_i_ssn\
        );

    \I__9200\ : InMux
    port map (
            O => \N__42689\,
            I => \N__42686\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__42686\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO\
        );

    \I__9198\ : InMux
    port map (
            O => \N__42683\,
            I => \N__42680\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__42680\,
            I => \N__42675\
        );

    \I__9196\ : InMux
    port map (
            O => \N__42679\,
            I => \N__42672\
        );

    \I__9195\ : InMux
    port map (
            O => \N__42678\,
            I => \N__42669\
        );

    \I__9194\ : Span12Mux_h
    port map (
            O => \N__42675\,
            I => \N__42666\
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__42672\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__42669\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2\
        );

    \I__9191\ : Odrv12
    port map (
            O => \N__42666\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2\
        );

    \I__9190\ : InMux
    port map (
            O => \N__42659\,
            I => \N__42656\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__42656\,
            I => \N__42653\
        );

    \I__9188\ : Odrv4
    port map (
            O => \N__42653\,
            I => \spi_data_misoZ0Z_0\
        );

    \I__9187\ : CascadeMux
    port map (
            O => \N__42650\,
            I => \N__42647\
        );

    \I__9186\ : InMux
    port map (
            O => \N__42647\,
            I => \N__42644\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__42644\,
            I => \sDAC_mem_4Z0Z_1\
        );

    \I__9184\ : CEMux
    port map (
            O => \N__42641\,
            I => \N__42637\
        );

    \I__9183\ : CEMux
    port map (
            O => \N__42640\,
            I => \N__42633\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__42637\,
            I => \N__42630\
        );

    \I__9181\ : CEMux
    port map (
            O => \N__42636\,
            I => \N__42627\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__42633\,
            I => \N__42619\
        );

    \I__9179\ : Span4Mux_h
    port map (
            O => \N__42630\,
            I => \N__42619\
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__42627\,
            I => \N__42619\
        );

    \I__9177\ : CEMux
    port map (
            O => \N__42626\,
            I => \N__42616\
        );

    \I__9176\ : Span4Mux_v
    port map (
            O => \N__42619\,
            I => \N__42613\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__42616\,
            I => \N__42610\
        );

    \I__9174\ : Span4Mux_h
    port map (
            O => \N__42613\,
            I => \N__42607\
        );

    \I__9173\ : Span12Mux_h
    port map (
            O => \N__42610\,
            I => \N__42604\
        );

    \I__9172\ : Sp12to4
    port map (
            O => \N__42607\,
            I => \N__42601\
        );

    \I__9171\ : Odrv12
    port map (
            O => \N__42604\,
            I => \sDAC_mem_4_1_sqmuxa\
        );

    \I__9170\ : Odrv12
    port map (
            O => \N__42601\,
            I => \sDAC_mem_4_1_sqmuxa\
        );

    \I__9169\ : CascadeMux
    port map (
            O => \N__42596\,
            I => \N__42592\
        );

    \I__9168\ : CascadeMux
    port map (
            O => \N__42595\,
            I => \N__42589\
        );

    \I__9167\ : InMux
    port map (
            O => \N__42592\,
            I => \N__42581\
        );

    \I__9166\ : InMux
    port map (
            O => \N__42589\,
            I => \N__42581\
        );

    \I__9165\ : InMux
    port map (
            O => \N__42588\,
            I => \N__42581\
        );

    \I__9164\ : LocalMux
    port map (
            O => \N__42581\,
            I => \N__42577\
        );

    \I__9163\ : CascadeMux
    port map (
            O => \N__42580\,
            I => \N__42571\
        );

    \I__9162\ : Span4Mux_v
    port map (
            O => \N__42577\,
            I => \N__42563\
        );

    \I__9161\ : InMux
    port map (
            O => \N__42576\,
            I => \N__42560\
        );

    \I__9160\ : CascadeMux
    port map (
            O => \N__42575\,
            I => \N__42553\
        );

    \I__9159\ : CascadeMux
    port map (
            O => \N__42574\,
            I => \N__42546\
        );

    \I__9158\ : InMux
    port map (
            O => \N__42571\,
            I => \N__42538\
        );

    \I__9157\ : InMux
    port map (
            O => \N__42570\,
            I => \N__42538\
        );

    \I__9156\ : InMux
    port map (
            O => \N__42569\,
            I => \N__42538\
        );

    \I__9155\ : InMux
    port map (
            O => \N__42568\,
            I => \N__42533\
        );

    \I__9154\ : InMux
    port map (
            O => \N__42567\,
            I => \N__42533\
        );

    \I__9153\ : InMux
    port map (
            O => \N__42566\,
            I => \N__42530\
        );

    \I__9152\ : Span4Mux_h
    port map (
            O => \N__42563\,
            I => \N__42516\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__42560\,
            I => \N__42516\
        );

    \I__9150\ : InMux
    port map (
            O => \N__42559\,
            I => \N__42507\
        );

    \I__9149\ : InMux
    port map (
            O => \N__42558\,
            I => \N__42500\
        );

    \I__9148\ : InMux
    port map (
            O => \N__42557\,
            I => \N__42500\
        );

    \I__9147\ : InMux
    port map (
            O => \N__42556\,
            I => \N__42500\
        );

    \I__9146\ : InMux
    port map (
            O => \N__42553\,
            I => \N__42493\
        );

    \I__9145\ : InMux
    port map (
            O => \N__42552\,
            I => \N__42493\
        );

    \I__9144\ : InMux
    port map (
            O => \N__42551\,
            I => \N__42493\
        );

    \I__9143\ : InMux
    port map (
            O => \N__42550\,
            I => \N__42490\
        );

    \I__9142\ : InMux
    port map (
            O => \N__42549\,
            I => \N__42483\
        );

    \I__9141\ : InMux
    port map (
            O => \N__42546\,
            I => \N__42483\
        );

    \I__9140\ : InMux
    port map (
            O => \N__42545\,
            I => \N__42483\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__42538\,
            I => \N__42478\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__42533\,
            I => \N__42478\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__42530\,
            I => \N__42475\
        );

    \I__9136\ : InMux
    port map (
            O => \N__42529\,
            I => \N__42470\
        );

    \I__9135\ : InMux
    port map (
            O => \N__42528\,
            I => \N__42470\
        );

    \I__9134\ : InMux
    port map (
            O => \N__42527\,
            I => \N__42465\
        );

    \I__9133\ : InMux
    port map (
            O => \N__42526\,
            I => \N__42465\
        );

    \I__9132\ : InMux
    port map (
            O => \N__42525\,
            I => \N__42462\
        );

    \I__9131\ : InMux
    port map (
            O => \N__42524\,
            I => \N__42455\
        );

    \I__9130\ : InMux
    port map (
            O => \N__42523\,
            I => \N__42455\
        );

    \I__9129\ : InMux
    port map (
            O => \N__42522\,
            I => \N__42455\
        );

    \I__9128\ : InMux
    port map (
            O => \N__42521\,
            I => \N__42452\
        );

    \I__9127\ : Span4Mux_v
    port map (
            O => \N__42516\,
            I => \N__42449\
        );

    \I__9126\ : InMux
    port map (
            O => \N__42515\,
            I => \N__42446\
        );

    \I__9125\ : InMux
    port map (
            O => \N__42514\,
            I => \N__42441\
        );

    \I__9124\ : InMux
    port map (
            O => \N__42513\,
            I => \N__42441\
        );

    \I__9123\ : InMux
    port map (
            O => \N__42512\,
            I => \N__42434\
        );

    \I__9122\ : InMux
    port map (
            O => \N__42511\,
            I => \N__42434\
        );

    \I__9121\ : InMux
    port map (
            O => \N__42510\,
            I => \N__42434\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__42507\,
            I => \N__42418\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__42500\,
            I => \N__42415\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__42493\,
            I => \N__42412\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__42490\,
            I => \N__42408\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__42483\,
            I => \N__42403\
        );

    \I__9115\ : Span4Mux_v
    port map (
            O => \N__42478\,
            I => \N__42403\
        );

    \I__9114\ : Span4Mux_v
    port map (
            O => \N__42475\,
            I => \N__42400\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__42470\,
            I => \N__42395\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__42465\,
            I => \N__42395\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__42462\,
            I => \N__42388\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__42455\,
            I => \N__42388\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__42452\,
            I => \N__42388\
        );

    \I__9108\ : Span4Mux_h
    port map (
            O => \N__42449\,
            I => \N__42379\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__42446\,
            I => \N__42379\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__42441\,
            I => \N__42379\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__42434\,
            I => \N__42379\
        );

    \I__9104\ : InMux
    port map (
            O => \N__42433\,
            I => \N__42376\
        );

    \I__9103\ : InMux
    port map (
            O => \N__42432\,
            I => \N__42373\
        );

    \I__9102\ : InMux
    port map (
            O => \N__42431\,
            I => \N__42370\
        );

    \I__9101\ : InMux
    port map (
            O => \N__42430\,
            I => \N__42367\
        );

    \I__9100\ : InMux
    port map (
            O => \N__42429\,
            I => \N__42360\
        );

    \I__9099\ : InMux
    port map (
            O => \N__42428\,
            I => \N__42360\
        );

    \I__9098\ : InMux
    port map (
            O => \N__42427\,
            I => \N__42360\
        );

    \I__9097\ : InMux
    port map (
            O => \N__42426\,
            I => \N__42357\
        );

    \I__9096\ : InMux
    port map (
            O => \N__42425\,
            I => \N__42352\
        );

    \I__9095\ : InMux
    port map (
            O => \N__42424\,
            I => \N__42352\
        );

    \I__9094\ : InMux
    port map (
            O => \N__42423\,
            I => \N__42347\
        );

    \I__9093\ : InMux
    port map (
            O => \N__42422\,
            I => \N__42347\
        );

    \I__9092\ : InMux
    port map (
            O => \N__42421\,
            I => \N__42344\
        );

    \I__9091\ : Span4Mux_h
    port map (
            O => \N__42418\,
            I => \N__42337\
        );

    \I__9090\ : Span4Mux_v
    port map (
            O => \N__42415\,
            I => \N__42337\
        );

    \I__9089\ : Span4Mux_v
    port map (
            O => \N__42412\,
            I => \N__42337\
        );

    \I__9088\ : InMux
    port map (
            O => \N__42411\,
            I => \N__42334\
        );

    \I__9087\ : Span4Mux_v
    port map (
            O => \N__42408\,
            I => \N__42325\
        );

    \I__9086\ : Span4Mux_h
    port map (
            O => \N__42403\,
            I => \N__42325\
        );

    \I__9085\ : Span4Mux_h
    port map (
            O => \N__42400\,
            I => \N__42325\
        );

    \I__9084\ : Span4Mux_v
    port map (
            O => \N__42395\,
            I => \N__42325\
        );

    \I__9083\ : Span4Mux_v
    port map (
            O => \N__42388\,
            I => \N__42320\
        );

    \I__9082\ : Span4Mux_v
    port map (
            O => \N__42379\,
            I => \N__42320\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__42376\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__42373\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__42370\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__42367\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__42360\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9076\ : LocalMux
    port map (
            O => \N__42357\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__42352\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__42347\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__42344\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9072\ : Odrv4
    port map (
            O => \N__42337\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__42334\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9070\ : Odrv4
    port map (
            O => \N__42325\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9069\ : Odrv4
    port map (
            O => \N__42320\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9068\ : InMux
    port map (
            O => \N__42293\,
            I => \N__42290\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__42290\,
            I => \N__42287\
        );

    \I__9066\ : Span4Mux_v
    port map (
            O => \N__42287\,
            I => \N__42284\
        );

    \I__9065\ : Span4Mux_v
    port map (
            O => \N__42284\,
            I => \N__42281\
        );

    \I__9064\ : Odrv4
    port map (
            O => \N__42281\,
            I => \sDAC_mem_36Z0Z_2\
        );

    \I__9063\ : InMux
    port map (
            O => \N__42278\,
            I => \N__42275\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__42275\,
            I => \N__42272\
        );

    \I__9061\ : Span12Mux_s11_h
    port map (
            O => \N__42272\,
            I => \N__42269\
        );

    \I__9060\ : Odrv12
    port map (
            O => \N__42269\,
            I => \sDAC_mem_4Z0Z_2\
        );

    \I__9059\ : CascadeMux
    port map (
            O => \N__42266\,
            I => \N__42260\
        );

    \I__9058\ : CascadeMux
    port map (
            O => \N__42265\,
            I => \N__42256\
        );

    \I__9057\ : CascadeMux
    port map (
            O => \N__42264\,
            I => \N__42253\
        );

    \I__9056\ : CascadeMux
    port map (
            O => \N__42263\,
            I => \N__42250\
        );

    \I__9055\ : InMux
    port map (
            O => \N__42260\,
            I => \N__42235\
        );

    \I__9054\ : InMux
    port map (
            O => \N__42259\,
            I => \N__42222\
        );

    \I__9053\ : InMux
    port map (
            O => \N__42256\,
            I => \N__42222\
        );

    \I__9052\ : InMux
    port map (
            O => \N__42253\,
            I => \N__42222\
        );

    \I__9051\ : InMux
    port map (
            O => \N__42250\,
            I => \N__42219\
        );

    \I__9050\ : CascadeMux
    port map (
            O => \N__42249\,
            I => \N__42215\
        );

    \I__9049\ : CascadeMux
    port map (
            O => \N__42248\,
            I => \N__42206\
        );

    \I__9048\ : CascadeMux
    port map (
            O => \N__42247\,
            I => \N__42199\
        );

    \I__9047\ : CascadeMux
    port map (
            O => \N__42246\,
            I => \N__42194\
        );

    \I__9046\ : CascadeMux
    port map (
            O => \N__42245\,
            I => \N__42185\
        );

    \I__9045\ : CascadeMux
    port map (
            O => \N__42244\,
            I => \N__42182\
        );

    \I__9044\ : InMux
    port map (
            O => \N__42243\,
            I => \N__42176\
        );

    \I__9043\ : InMux
    port map (
            O => \N__42242\,
            I => \N__42176\
        );

    \I__9042\ : CascadeMux
    port map (
            O => \N__42241\,
            I => \N__42162\
        );

    \I__9041\ : CascadeMux
    port map (
            O => \N__42240\,
            I => \N__42158\
        );

    \I__9040\ : CascadeMux
    port map (
            O => \N__42239\,
            I => \N__42154\
        );

    \I__9039\ : CascadeMux
    port map (
            O => \N__42238\,
            I => \N__42150\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__42235\,
            I => \N__42139\
        );

    \I__9037\ : InMux
    port map (
            O => \N__42234\,
            I => \N__42132\
        );

    \I__9036\ : InMux
    port map (
            O => \N__42233\,
            I => \N__42132\
        );

    \I__9035\ : InMux
    port map (
            O => \N__42232\,
            I => \N__42132\
        );

    \I__9034\ : InMux
    port map (
            O => \N__42231\,
            I => \N__42125\
        );

    \I__9033\ : InMux
    port map (
            O => \N__42230\,
            I => \N__42125\
        );

    \I__9032\ : InMux
    port map (
            O => \N__42229\,
            I => \N__42125\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__42222\,
            I => \N__42120\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__42219\,
            I => \N__42120\
        );

    \I__9029\ : InMux
    port map (
            O => \N__42218\,
            I => \N__42115\
        );

    \I__9028\ : InMux
    port map (
            O => \N__42215\,
            I => \N__42115\
        );

    \I__9027\ : CascadeMux
    port map (
            O => \N__42214\,
            I => \N__42106\
        );

    \I__9026\ : CascadeMux
    port map (
            O => \N__42213\,
            I => \N__42101\
        );

    \I__9025\ : CascadeMux
    port map (
            O => \N__42212\,
            I => \N__42098\
        );

    \I__9024\ : InMux
    port map (
            O => \N__42211\,
            I => \N__42090\
        );

    \I__9023\ : InMux
    port map (
            O => \N__42210\,
            I => \N__42083\
        );

    \I__9022\ : InMux
    port map (
            O => \N__42209\,
            I => \N__42083\
        );

    \I__9021\ : InMux
    port map (
            O => \N__42206\,
            I => \N__42083\
        );

    \I__9020\ : CascadeMux
    port map (
            O => \N__42205\,
            I => \N__42077\
        );

    \I__9019\ : CascadeMux
    port map (
            O => \N__42204\,
            I => \N__42069\
        );

    \I__9018\ : CascadeMux
    port map (
            O => \N__42203\,
            I => \N__42064\
        );

    \I__9017\ : InMux
    port map (
            O => \N__42202\,
            I => \N__42053\
        );

    \I__9016\ : InMux
    port map (
            O => \N__42199\,
            I => \N__42053\
        );

    \I__9015\ : InMux
    port map (
            O => \N__42198\,
            I => \N__42053\
        );

    \I__9014\ : InMux
    port map (
            O => \N__42197\,
            I => \N__42053\
        );

    \I__9013\ : InMux
    port map (
            O => \N__42194\,
            I => \N__42053\
        );

    \I__9012\ : CascadeMux
    port map (
            O => \N__42193\,
            I => \N__42049\
        );

    \I__9011\ : CascadeMux
    port map (
            O => \N__42192\,
            I => \N__42046\
        );

    \I__9010\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42039\
        );

    \I__9009\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42039\
        );

    \I__9008\ : InMux
    port map (
            O => \N__42189\,
            I => \N__42039\
        );

    \I__9007\ : InMux
    port map (
            O => \N__42188\,
            I => \N__42029\
        );

    \I__9006\ : InMux
    port map (
            O => \N__42185\,
            I => \N__42022\
        );

    \I__9005\ : InMux
    port map (
            O => \N__42182\,
            I => \N__42022\
        );

    \I__9004\ : InMux
    port map (
            O => \N__42181\,
            I => \N__42022\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__42176\,
            I => \N__42019\
        );

    \I__9002\ : CascadeMux
    port map (
            O => \N__42175\,
            I => \N__42007\
        );

    \I__9001\ : CascadeMux
    port map (
            O => \N__42174\,
            I => \N__42003\
        );

    \I__9000\ : CascadeMux
    port map (
            O => \N__42173\,
            I => \N__41997\
        );

    \I__8999\ : CascadeMux
    port map (
            O => \N__42172\,
            I => \N__41994\
        );

    \I__8998\ : CascadeMux
    port map (
            O => \N__42171\,
            I => \N__41991\
        );

    \I__8997\ : CascadeMux
    port map (
            O => \N__42170\,
            I => \N__41979\
        );

    \I__8996\ : CascadeMux
    port map (
            O => \N__42169\,
            I => \N__41976\
        );

    \I__8995\ : InMux
    port map (
            O => \N__42168\,
            I => \N__41972\
        );

    \I__8994\ : InMux
    port map (
            O => \N__42167\,
            I => \N__41965\
        );

    \I__8993\ : InMux
    port map (
            O => \N__42166\,
            I => \N__41965\
        );

    \I__8992\ : InMux
    port map (
            O => \N__42165\,
            I => \N__41965\
        );

    \I__8991\ : InMux
    port map (
            O => \N__42162\,
            I => \N__41958\
        );

    \I__8990\ : InMux
    port map (
            O => \N__42161\,
            I => \N__41958\
        );

    \I__8989\ : InMux
    port map (
            O => \N__42158\,
            I => \N__41958\
        );

    \I__8988\ : InMux
    port map (
            O => \N__42157\,
            I => \N__41953\
        );

    \I__8987\ : InMux
    port map (
            O => \N__42154\,
            I => \N__41953\
        );

    \I__8986\ : InMux
    port map (
            O => \N__42153\,
            I => \N__41944\
        );

    \I__8985\ : InMux
    port map (
            O => \N__42150\,
            I => \N__41944\
        );

    \I__8984\ : InMux
    port map (
            O => \N__42149\,
            I => \N__41944\
        );

    \I__8983\ : InMux
    port map (
            O => \N__42148\,
            I => \N__41944\
        );

    \I__8982\ : InMux
    port map (
            O => \N__42147\,
            I => \N__41937\
        );

    \I__8981\ : InMux
    port map (
            O => \N__42146\,
            I => \N__41937\
        );

    \I__8980\ : InMux
    port map (
            O => \N__42145\,
            I => \N__41937\
        );

    \I__8979\ : InMux
    port map (
            O => \N__42144\,
            I => \N__41932\
        );

    \I__8978\ : InMux
    port map (
            O => \N__42143\,
            I => \N__41932\
        );

    \I__8977\ : InMux
    port map (
            O => \N__42142\,
            I => \N__41929\
        );

    \I__8976\ : Span4Mux_v
    port map (
            O => \N__42139\,
            I => \N__41918\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__42132\,
            I => \N__41918\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__42125\,
            I => \N__41918\
        );

    \I__8973\ : Span4Mux_h
    port map (
            O => \N__42120\,
            I => \N__41918\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__42115\,
            I => \N__41918\
        );

    \I__8971\ : InMux
    port map (
            O => \N__42114\,
            I => \N__41911\
        );

    \I__8970\ : InMux
    port map (
            O => \N__42113\,
            I => \N__41911\
        );

    \I__8969\ : InMux
    port map (
            O => \N__42112\,
            I => \N__41911\
        );

    \I__8968\ : InMux
    port map (
            O => \N__42111\,
            I => \N__41898\
        );

    \I__8967\ : InMux
    port map (
            O => \N__42110\,
            I => \N__41898\
        );

    \I__8966\ : InMux
    port map (
            O => \N__42109\,
            I => \N__41898\
        );

    \I__8965\ : InMux
    port map (
            O => \N__42106\,
            I => \N__41898\
        );

    \I__8964\ : InMux
    port map (
            O => \N__42105\,
            I => \N__41898\
        );

    \I__8963\ : InMux
    port map (
            O => \N__42104\,
            I => \N__41898\
        );

    \I__8962\ : InMux
    port map (
            O => \N__42101\,
            I => \N__41893\
        );

    \I__8961\ : InMux
    port map (
            O => \N__42098\,
            I => \N__41893\
        );

    \I__8960\ : CascadeMux
    port map (
            O => \N__42097\,
            I => \N__41888\
        );

    \I__8959\ : InMux
    port map (
            O => \N__42096\,
            I => \N__41879\
        );

    \I__8958\ : InMux
    port map (
            O => \N__42095\,
            I => \N__41879\
        );

    \I__8957\ : InMux
    port map (
            O => \N__42094\,
            I => \N__41876\
        );

    \I__8956\ : InMux
    port map (
            O => \N__42093\,
            I => \N__41869\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__42090\,
            I => \N__41856\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__42083\,
            I => \N__41856\
        );

    \I__8953\ : InMux
    port map (
            O => \N__42082\,
            I => \N__41851\
        );

    \I__8952\ : InMux
    port map (
            O => \N__42081\,
            I => \N__41851\
        );

    \I__8951\ : InMux
    port map (
            O => \N__42080\,
            I => \N__41842\
        );

    \I__8950\ : InMux
    port map (
            O => \N__42077\,
            I => \N__41842\
        );

    \I__8949\ : InMux
    port map (
            O => \N__42076\,
            I => \N__41842\
        );

    \I__8948\ : InMux
    port map (
            O => \N__42075\,
            I => \N__41842\
        );

    \I__8947\ : CascadeMux
    port map (
            O => \N__42074\,
            I => \N__41838\
        );

    \I__8946\ : InMux
    port map (
            O => \N__42073\,
            I => \N__41831\
        );

    \I__8945\ : InMux
    port map (
            O => \N__42072\,
            I => \N__41831\
        );

    \I__8944\ : InMux
    port map (
            O => \N__42069\,
            I => \N__41831\
        );

    \I__8943\ : InMux
    port map (
            O => \N__42068\,
            I => \N__41824\
        );

    \I__8942\ : InMux
    port map (
            O => \N__42067\,
            I => \N__41824\
        );

    \I__8941\ : InMux
    port map (
            O => \N__42064\,
            I => \N__41824\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__42053\,
            I => \N__41821\
        );

    \I__8939\ : InMux
    port map (
            O => \N__42052\,
            I => \N__41814\
        );

    \I__8938\ : InMux
    port map (
            O => \N__42049\,
            I => \N__41814\
        );

    \I__8937\ : InMux
    port map (
            O => \N__42046\,
            I => \N__41814\
        );

    \I__8936\ : LocalMux
    port map (
            O => \N__42039\,
            I => \N__41801\
        );

    \I__8935\ : InMux
    port map (
            O => \N__42038\,
            I => \N__41792\
        );

    \I__8934\ : InMux
    port map (
            O => \N__42037\,
            I => \N__41792\
        );

    \I__8933\ : InMux
    port map (
            O => \N__42036\,
            I => \N__41792\
        );

    \I__8932\ : InMux
    port map (
            O => \N__42035\,
            I => \N__41792\
        );

    \I__8931\ : InMux
    port map (
            O => \N__42034\,
            I => \N__41785\
        );

    \I__8930\ : InMux
    port map (
            O => \N__42033\,
            I => \N__41785\
        );

    \I__8929\ : InMux
    port map (
            O => \N__42032\,
            I => \N__41785\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__42029\,
            I => \N__41780\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__42022\,
            I => \N__41780\
        );

    \I__8926\ : Span4Mux_v
    port map (
            O => \N__42019\,
            I => \N__41777\
        );

    \I__8925\ : InMux
    port map (
            O => \N__42018\,
            I => \N__41768\
        );

    \I__8924\ : InMux
    port map (
            O => \N__42017\,
            I => \N__41768\
        );

    \I__8923\ : InMux
    port map (
            O => \N__42016\,
            I => \N__41768\
        );

    \I__8922\ : InMux
    port map (
            O => \N__42015\,
            I => \N__41768\
        );

    \I__8921\ : InMux
    port map (
            O => \N__42014\,
            I => \N__41763\
        );

    \I__8920\ : InMux
    port map (
            O => \N__42013\,
            I => \N__41763\
        );

    \I__8919\ : InMux
    port map (
            O => \N__42012\,
            I => \N__41756\
        );

    \I__8918\ : InMux
    port map (
            O => \N__42011\,
            I => \N__41756\
        );

    \I__8917\ : InMux
    port map (
            O => \N__42010\,
            I => \N__41756\
        );

    \I__8916\ : InMux
    port map (
            O => \N__42007\,
            I => \N__41749\
        );

    \I__8915\ : InMux
    port map (
            O => \N__42006\,
            I => \N__41749\
        );

    \I__8914\ : InMux
    port map (
            O => \N__42003\,
            I => \N__41749\
        );

    \I__8913\ : InMux
    port map (
            O => \N__42002\,
            I => \N__41744\
        );

    \I__8912\ : InMux
    port map (
            O => \N__42001\,
            I => \N__41744\
        );

    \I__8911\ : InMux
    port map (
            O => \N__42000\,
            I => \N__41735\
        );

    \I__8910\ : InMux
    port map (
            O => \N__41997\,
            I => \N__41735\
        );

    \I__8909\ : InMux
    port map (
            O => \N__41994\,
            I => \N__41735\
        );

    \I__8908\ : InMux
    port map (
            O => \N__41991\,
            I => \N__41735\
        );

    \I__8907\ : InMux
    port map (
            O => \N__41990\,
            I => \N__41730\
        );

    \I__8906\ : InMux
    port map (
            O => \N__41989\,
            I => \N__41730\
        );

    \I__8905\ : InMux
    port map (
            O => \N__41988\,
            I => \N__41723\
        );

    \I__8904\ : InMux
    port map (
            O => \N__41987\,
            I => \N__41723\
        );

    \I__8903\ : InMux
    port map (
            O => \N__41986\,
            I => \N__41723\
        );

    \I__8902\ : InMux
    port map (
            O => \N__41985\,
            I => \N__41717\
        );

    \I__8901\ : InMux
    port map (
            O => \N__41984\,
            I => \N__41712\
        );

    \I__8900\ : InMux
    port map (
            O => \N__41983\,
            I => \N__41712\
        );

    \I__8899\ : InMux
    port map (
            O => \N__41982\,
            I => \N__41709\
        );

    \I__8898\ : InMux
    port map (
            O => \N__41979\,
            I => \N__41702\
        );

    \I__8897\ : InMux
    port map (
            O => \N__41976\,
            I => \N__41702\
        );

    \I__8896\ : InMux
    port map (
            O => \N__41975\,
            I => \N__41702\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__41972\,
            I => \N__41689\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__41965\,
            I => \N__41689\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__41958\,
            I => \N__41689\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__41953\,
            I => \N__41689\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__41944\,
            I => \N__41689\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__41937\,
            I => \N__41689\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__41932\,
            I => \N__41684\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__41929\,
            I => \N__41684\
        );

    \I__8887\ : Span4Mux_h
    port map (
            O => \N__41918\,
            I => \N__41675\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__41911\,
            I => \N__41675\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__41898\,
            I => \N__41675\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__41893\,
            I => \N__41675\
        );

    \I__8883\ : InMux
    port map (
            O => \N__41892\,
            I => \N__41666\
        );

    \I__8882\ : InMux
    port map (
            O => \N__41891\,
            I => \N__41666\
        );

    \I__8881\ : InMux
    port map (
            O => \N__41888\,
            I => \N__41666\
        );

    \I__8880\ : InMux
    port map (
            O => \N__41887\,
            I => \N__41666\
        );

    \I__8879\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41659\
        );

    \I__8878\ : InMux
    port map (
            O => \N__41885\,
            I => \N__41659\
        );

    \I__8877\ : InMux
    port map (
            O => \N__41884\,
            I => \N__41659\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__41879\,
            I => \N__41652\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__41876\,
            I => \N__41652\
        );

    \I__8874\ : InMux
    port map (
            O => \N__41875\,
            I => \N__41643\
        );

    \I__8873\ : InMux
    port map (
            O => \N__41874\,
            I => \N__41643\
        );

    \I__8872\ : InMux
    port map (
            O => \N__41873\,
            I => \N__41643\
        );

    \I__8871\ : InMux
    port map (
            O => \N__41872\,
            I => \N__41643\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__41869\,
            I => \N__41640\
        );

    \I__8869\ : InMux
    port map (
            O => \N__41868\,
            I => \N__41631\
        );

    \I__8868\ : InMux
    port map (
            O => \N__41867\,
            I => \N__41631\
        );

    \I__8867\ : InMux
    port map (
            O => \N__41866\,
            I => \N__41631\
        );

    \I__8866\ : InMux
    port map (
            O => \N__41865\,
            I => \N__41631\
        );

    \I__8865\ : InMux
    port map (
            O => \N__41864\,
            I => \N__41622\
        );

    \I__8864\ : InMux
    port map (
            O => \N__41863\,
            I => \N__41622\
        );

    \I__8863\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41622\
        );

    \I__8862\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41622\
        );

    \I__8861\ : Span4Mux_v
    port map (
            O => \N__41856\,
            I => \N__41615\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__41851\,
            I => \N__41615\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__41842\,
            I => \N__41615\
        );

    \I__8858\ : InMux
    port map (
            O => \N__41841\,
            I => \N__41610\
        );

    \I__8857\ : InMux
    port map (
            O => \N__41838\,
            I => \N__41610\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__41831\,
            I => \N__41596\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__41824\,
            I => \N__41596\
        );

    \I__8854\ : Span4Mux_v
    port map (
            O => \N__41821\,
            I => \N__41596\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__41814\,
            I => \N__41596\
        );

    \I__8852\ : InMux
    port map (
            O => \N__41813\,
            I => \N__41587\
        );

    \I__8851\ : InMux
    port map (
            O => \N__41812\,
            I => \N__41587\
        );

    \I__8850\ : InMux
    port map (
            O => \N__41811\,
            I => \N__41587\
        );

    \I__8849\ : InMux
    port map (
            O => \N__41810\,
            I => \N__41587\
        );

    \I__8848\ : InMux
    port map (
            O => \N__41809\,
            I => \N__41582\
        );

    \I__8847\ : InMux
    port map (
            O => \N__41808\,
            I => \N__41582\
        );

    \I__8846\ : InMux
    port map (
            O => \N__41807\,
            I => \N__41579\
        );

    \I__8845\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41572\
        );

    \I__8844\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41572\
        );

    \I__8843\ : InMux
    port map (
            O => \N__41804\,
            I => \N__41572\
        );

    \I__8842\ : Span4Mux_v
    port map (
            O => \N__41801\,
            I => \N__41567\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__41792\,
            I => \N__41567\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__41785\,
            I => \N__41560\
        );

    \I__8839\ : Span4Mux_v
    port map (
            O => \N__41780\,
            I => \N__41557\
        );

    \I__8838\ : Span4Mux_h
    port map (
            O => \N__41777\,
            I => \N__41548\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__41768\,
            I => \N__41548\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__41763\,
            I => \N__41548\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__41756\,
            I => \N__41548\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__41749\,
            I => \N__41541\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__41744\,
            I => \N__41541\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__41735\,
            I => \N__41541\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__41730\,
            I => \N__41538\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__41723\,
            I => \N__41533\
        );

    \I__8829\ : InMux
    port map (
            O => \N__41722\,
            I => \N__41526\
        );

    \I__8828\ : InMux
    port map (
            O => \N__41721\,
            I => \N__41526\
        );

    \I__8827\ : InMux
    port map (
            O => \N__41720\,
            I => \N__41526\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__41717\,
            I => \N__41523\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__41712\,
            I => \N__41506\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__41709\,
            I => \N__41506\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__41702\,
            I => \N__41506\
        );

    \I__8822\ : Span4Mux_v
    port map (
            O => \N__41689\,
            I => \N__41506\
        );

    \I__8821\ : Span4Mux_h
    port map (
            O => \N__41684\,
            I => \N__41506\
        );

    \I__8820\ : Span4Mux_v
    port map (
            O => \N__41675\,
            I => \N__41506\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__41666\,
            I => \N__41506\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__41659\,
            I => \N__41506\
        );

    \I__8817\ : InMux
    port map (
            O => \N__41658\,
            I => \N__41501\
        );

    \I__8816\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41501\
        );

    \I__8815\ : Span4Mux_h
    port map (
            O => \N__41652\,
            I => \N__41494\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__41643\,
            I => \N__41494\
        );

    \I__8813\ : Span4Mux_v
    port map (
            O => \N__41640\,
            I => \N__41494\
        );

    \I__8812\ : LocalMux
    port map (
            O => \N__41631\,
            I => \N__41489\
        );

    \I__8811\ : LocalMux
    port map (
            O => \N__41622\,
            I => \N__41489\
        );

    \I__8810\ : Span4Mux_h
    port map (
            O => \N__41615\,
            I => \N__41484\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__41610\,
            I => \N__41484\
        );

    \I__8808\ : InMux
    port map (
            O => \N__41609\,
            I => \N__41479\
        );

    \I__8807\ : InMux
    port map (
            O => \N__41608\,
            I => \N__41479\
        );

    \I__8806\ : InMux
    port map (
            O => \N__41607\,
            I => \N__41476\
        );

    \I__8805\ : InMux
    port map (
            O => \N__41606\,
            I => \N__41471\
        );

    \I__8804\ : InMux
    port map (
            O => \N__41605\,
            I => \N__41471\
        );

    \I__8803\ : Sp12to4
    port map (
            O => \N__41596\,
            I => \N__41464\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__41587\,
            I => \N__41464\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__41582\,
            I => \N__41464\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__41579\,
            I => \N__41457\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__41572\,
            I => \N__41457\
        );

    \I__8798\ : Span4Mux_v
    port map (
            O => \N__41567\,
            I => \N__41457\
        );

    \I__8797\ : InMux
    port map (
            O => \N__41566\,
            I => \N__41448\
        );

    \I__8796\ : InMux
    port map (
            O => \N__41565\,
            I => \N__41448\
        );

    \I__8795\ : InMux
    port map (
            O => \N__41564\,
            I => \N__41448\
        );

    \I__8794\ : InMux
    port map (
            O => \N__41563\,
            I => \N__41448\
        );

    \I__8793\ : Span4Mux_v
    port map (
            O => \N__41560\,
            I => \N__41441\
        );

    \I__8792\ : Span4Mux_h
    port map (
            O => \N__41557\,
            I => \N__41441\
        );

    \I__8791\ : Span4Mux_v
    port map (
            O => \N__41548\,
            I => \N__41441\
        );

    \I__8790\ : Span12Mux_h
    port map (
            O => \N__41541\,
            I => \N__41436\
        );

    \I__8789\ : Span12Mux_h
    port map (
            O => \N__41538\,
            I => \N__41436\
        );

    \I__8788\ : InMux
    port map (
            O => \N__41537\,
            I => \N__41431\
        );

    \I__8787\ : InMux
    port map (
            O => \N__41536\,
            I => \N__41431\
        );

    \I__8786\ : Span4Mux_h
    port map (
            O => \N__41533\,
            I => \N__41424\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__41526\,
            I => \N__41424\
        );

    \I__8784\ : Span4Mux_v
    port map (
            O => \N__41523\,
            I => \N__41424\
        );

    \I__8783\ : Span4Mux_v
    port map (
            O => \N__41506\,
            I => \N__41419\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__41501\,
            I => \N__41419\
        );

    \I__8781\ : Span4Mux_v
    port map (
            O => \N__41494\,
            I => \N__41412\
        );

    \I__8780\ : Span4Mux_v
    port map (
            O => \N__41489\,
            I => \N__41412\
        );

    \I__8779\ : Span4Mux_h
    port map (
            O => \N__41484\,
            I => \N__41412\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__41479\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__41476\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__41471\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8775\ : Odrv12
    port map (
            O => \N__41464\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8774\ : Odrv4
    port map (
            O => \N__41457\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__41448\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8772\ : Odrv4
    port map (
            O => \N__41441\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8771\ : Odrv12
    port map (
            O => \N__41436\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__41431\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8769\ : Odrv4
    port map (
            O => \N__41424\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8768\ : Odrv4
    port map (
            O => \N__41419\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8767\ : Odrv4
    port map (
            O => \N__41412\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__8766\ : InMux
    port map (
            O => \N__41387\,
            I => \N__41384\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__41384\,
            I => \N__41381\
        );

    \I__8764\ : Odrv4
    port map (
            O => \N__41381\,
            I => \sDAC_mem_37Z0Z_2\
        );

    \I__8763\ : CascadeMux
    port map (
            O => \N__41378\,
            I => \sDAC_data_2_13_am_1_5_cascade_\
        );

    \I__8762\ : InMux
    port map (
            O => \N__41375\,
            I => \N__41372\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__41372\,
            I => \sDAC_data_RNO_4Z0Z_5\
        );

    \I__8760\ : InMux
    port map (
            O => \N__41369\,
            I => \N__41366\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__41366\,
            I => \N__41363\
        );

    \I__8758\ : Span4Mux_h
    port map (
            O => \N__41363\,
            I => \N__41360\
        );

    \I__8757\ : Odrv4
    port map (
            O => \N__41360\,
            I => \sDAC_mem_25Z0Z_5\
        );

    \I__8756\ : InMux
    port map (
            O => \N__41357\,
            I => \N__41354\
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__41354\,
            I => \N__41351\
        );

    \I__8754\ : Span4Mux_h
    port map (
            O => \N__41351\,
            I => \N__41348\
        );

    \I__8753\ : Odrv4
    port map (
            O => \N__41348\,
            I => \sDAC_mem_25Z0Z_2\
        );

    \I__8752\ : InMux
    port map (
            O => \N__41345\,
            I => \N__41342\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__41342\,
            I => \sDAC_mem_25Z0Z_3\
        );

    \I__8750\ : InMux
    port map (
            O => \N__41339\,
            I => \N__41336\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__41336\,
            I => \N__41333\
        );

    \I__8748\ : Span4Mux_h
    port map (
            O => \N__41333\,
            I => \N__41330\
        );

    \I__8747\ : Span4Mux_h
    port map (
            O => \N__41330\,
            I => \N__41327\
        );

    \I__8746\ : Odrv4
    port map (
            O => \N__41327\,
            I => \sDAC_mem_25Z0Z_4\
        );

    \I__8745\ : InMux
    port map (
            O => \N__41324\,
            I => \N__41321\
        );

    \I__8744\ : LocalMux
    port map (
            O => \N__41321\,
            I => \N__41318\
        );

    \I__8743\ : Span4Mux_h
    port map (
            O => \N__41318\,
            I => \N__41315\
        );

    \I__8742\ : Odrv4
    port map (
            O => \N__41315\,
            I => \sDAC_mem_25Z0Z_0\
        );

    \I__8741\ : InMux
    port map (
            O => \N__41312\,
            I => \N__41309\
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__41309\,
            I => \N__41306\
        );

    \I__8739\ : Span4Mux_h
    port map (
            O => \N__41306\,
            I => \N__41303\
        );

    \I__8738\ : Span4Mux_h
    port map (
            O => \N__41303\,
            I => \N__41300\
        );

    \I__8737\ : Odrv4
    port map (
            O => \N__41300\,
            I => \sDAC_mem_25Z0Z_6\
        );

    \I__8736\ : InMux
    port map (
            O => \N__41297\,
            I => \N__41294\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__41294\,
            I => \sDAC_mem_32Z0Z_1\
        );

    \I__8734\ : CascadeMux
    port map (
            O => \N__41291\,
            I => \sDAC_data_RNO_26Z0Z_5_cascade_\
        );

    \I__8733\ : InMux
    port map (
            O => \N__41288\,
            I => \N__41285\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__41285\,
            I => \sDAC_data_RNO_14Z0Z_5\
        );

    \I__8731\ : InMux
    port map (
            O => \N__41282\,
            I => \N__41279\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__41279\,
            I => \sDAC_mem_32Z0Z_2\
        );

    \I__8729\ : CEMux
    port map (
            O => \N__41276\,
            I => \N__41272\
        );

    \I__8728\ : CEMux
    port map (
            O => \N__41275\,
            I => \N__41269\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__41272\,
            I => \N__41266\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__41269\,
            I => \N__41262\
        );

    \I__8725\ : Span4Mux_h
    port map (
            O => \N__41266\,
            I => \N__41259\
        );

    \I__8724\ : CEMux
    port map (
            O => \N__41265\,
            I => \N__41255\
        );

    \I__8723\ : Span4Mux_h
    port map (
            O => \N__41262\,
            I => \N__41252\
        );

    \I__8722\ : Span4Mux_v
    port map (
            O => \N__41259\,
            I => \N__41249\
        );

    \I__8721\ : CEMux
    port map (
            O => \N__41258\,
            I => \N__41246\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__41255\,
            I => \N__41243\
        );

    \I__8719\ : Span4Mux_h
    port map (
            O => \N__41252\,
            I => \N__41240\
        );

    \I__8718\ : Span4Mux_h
    port map (
            O => \N__41249\,
            I => \N__41237\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__41246\,
            I => \N__41234\
        );

    \I__8716\ : Span4Mux_v
    port map (
            O => \N__41243\,
            I => \N__41231\
        );

    \I__8715\ : Span4Mux_h
    port map (
            O => \N__41240\,
            I => \N__41226\
        );

    \I__8714\ : Span4Mux_h
    port map (
            O => \N__41237\,
            I => \N__41226\
        );

    \I__8713\ : Span12Mux_h
    port map (
            O => \N__41234\,
            I => \N__41223\
        );

    \I__8712\ : Span4Mux_h
    port map (
            O => \N__41231\,
            I => \N__41220\
        );

    \I__8711\ : Odrv4
    port map (
            O => \N__41226\,
            I => \sDAC_mem_32_1_sqmuxa\
        );

    \I__8710\ : Odrv12
    port map (
            O => \N__41223\,
            I => \sDAC_mem_32_1_sqmuxa\
        );

    \I__8709\ : Odrv4
    port map (
            O => \N__41220\,
            I => \sDAC_mem_32_1_sqmuxa\
        );

    \I__8708\ : InMux
    port map (
            O => \N__41213\,
            I => \N__41210\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__41210\,
            I => \N__41207\
        );

    \I__8706\ : Span12Mux_h
    port map (
            O => \N__41207\,
            I => \N__41204\
        );

    \I__8705\ : Odrv12
    port map (
            O => \N__41204\,
            I => \sDAC_mem_36Z0Z_0\
        );

    \I__8704\ : InMux
    port map (
            O => \N__41201\,
            I => \N__41198\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__41198\,
            I => \N__41195\
        );

    \I__8702\ : Odrv4
    port map (
            O => \N__41195\,
            I => \sDAC_mem_37Z0Z_0\
        );

    \I__8701\ : CascadeMux
    port map (
            O => \N__41192\,
            I => \sDAC_data_2_13_am_1_3_cascade_\
        );

    \I__8700\ : CascadeMux
    port map (
            O => \N__41189\,
            I => \N__41186\
        );

    \I__8699\ : InMux
    port map (
            O => \N__41186\,
            I => \N__41183\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__41183\,
            I => \N__41180\
        );

    \I__8697\ : Odrv4
    port map (
            O => \N__41180\,
            I => \sDAC_data_RNO_4Z0Z_3\
        );

    \I__8696\ : InMux
    port map (
            O => \N__41177\,
            I => \N__41174\
        );

    \I__8695\ : LocalMux
    port map (
            O => \N__41174\,
            I => \sDAC_mem_4Z0Z_0\
        );

    \I__8694\ : InMux
    port map (
            O => \N__41171\,
            I => \N__41168\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__41168\,
            I => \N__41165\
        );

    \I__8692\ : Span4Mux_v
    port map (
            O => \N__41165\,
            I => \N__41162\
        );

    \I__8691\ : Span4Mux_v
    port map (
            O => \N__41162\,
            I => \N__41159\
        );

    \I__8690\ : Odrv4
    port map (
            O => \N__41159\,
            I => \sDAC_mem_36Z0Z_1\
        );

    \I__8689\ : CascadeMux
    port map (
            O => \N__41156\,
            I => \sDAC_data_2_13_am_1_4_cascade_\
        );

    \I__8688\ : InMux
    port map (
            O => \N__41153\,
            I => \N__41150\
        );

    \I__8687\ : LocalMux
    port map (
            O => \N__41150\,
            I => \N__41147\
        );

    \I__8686\ : Odrv4
    port map (
            O => \N__41147\,
            I => \sDAC_mem_37Z0Z_1\
        );

    \I__8685\ : InMux
    port map (
            O => \N__41144\,
            I => \N__41141\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__41141\,
            I => \N__41138\
        );

    \I__8683\ : Span4Mux_v
    port map (
            O => \N__41138\,
            I => \N__41135\
        );

    \I__8682\ : Odrv4
    port map (
            O => \N__41135\,
            I => \sDAC_data_RNO_4Z0Z_4\
        );

    \I__8681\ : InMux
    port map (
            O => \N__41132\,
            I => \N__41129\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__41129\,
            I => \N__41126\
        );

    \I__8679\ : Odrv12
    port map (
            O => \N__41126\,
            I => \sDAC_mem_37Z0Z_3\
        );

    \I__8678\ : InMux
    port map (
            O => \N__41123\,
            I => \N__41120\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__41120\,
            I => \N__41117\
        );

    \I__8676\ : Span4Mux_h
    port map (
            O => \N__41117\,
            I => \N__41114\
        );

    \I__8675\ : Odrv4
    port map (
            O => \N__41114\,
            I => \sDAC_mem_37Z0Z_4\
        );

    \I__8674\ : InMux
    port map (
            O => \N__41111\,
            I => \N__41108\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__41108\,
            I => \N__41105\
        );

    \I__8672\ : Span4Mux_h
    port map (
            O => \N__41105\,
            I => \N__41102\
        );

    \I__8671\ : Odrv4
    port map (
            O => \N__41102\,
            I => \sDAC_mem_37Z0Z_5\
        );

    \I__8670\ : InMux
    port map (
            O => \N__41099\,
            I => \N__41096\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__41096\,
            I => \N__41093\
        );

    \I__8668\ : Span4Mux_v
    port map (
            O => \N__41093\,
            I => \N__41090\
        );

    \I__8667\ : Odrv4
    port map (
            O => \N__41090\,
            I => \sDAC_mem_37Z0Z_6\
        );

    \I__8666\ : InMux
    port map (
            O => \N__41087\,
            I => \N__41084\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__41084\,
            I => \N__41081\
        );

    \I__8664\ : Span4Mux_h
    port map (
            O => \N__41081\,
            I => \N__41078\
        );

    \I__8663\ : Odrv4
    port map (
            O => \N__41078\,
            I => \sDAC_mem_37Z0Z_7\
        );

    \I__8662\ : CEMux
    port map (
            O => \N__41075\,
            I => \N__41072\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__41072\,
            I => \N__41069\
        );

    \I__8660\ : Span4Mux_h
    port map (
            O => \N__41069\,
            I => \N__41066\
        );

    \I__8659\ : Span4Mux_h
    port map (
            O => \N__41066\,
            I => \N__41063\
        );

    \I__8658\ : Odrv4
    port map (
            O => \N__41063\,
            I => \sDAC_mem_37_1_sqmuxa\
        );

    \I__8657\ : InMux
    port map (
            O => \N__41060\,
            I => \N__41057\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__41057\,
            I => \sDAC_data_RNO_26Z0Z_3\
        );

    \I__8655\ : InMux
    port map (
            O => \N__41054\,
            I => \N__41051\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__41051\,
            I => \sDAC_data_RNO_14Z0Z_3\
        );

    \I__8653\ : CascadeMux
    port map (
            O => \N__41048\,
            I => \sDAC_data_RNO_26Z0Z_4_cascade_\
        );

    \I__8652\ : InMux
    port map (
            O => \N__41045\,
            I => \N__41042\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__41042\,
            I => \N__41039\
        );

    \I__8650\ : Span4Mux_v
    port map (
            O => \N__41039\,
            I => \N__41036\
        );

    \I__8649\ : Odrv4
    port map (
            O => \N__41036\,
            I => \sDAC_data_RNO_14Z0Z_4\
        );

    \I__8648\ : InMux
    port map (
            O => \N__41033\,
            I => \N__41030\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__41030\,
            I => \sDAC_mem_32Z0Z_0\
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__41027\,
            I => \N__41023\
        );

    \I__8645\ : InMux
    port map (
            O => \N__41026\,
            I => \N__41018\
        );

    \I__8644\ : InMux
    port map (
            O => \N__41023\,
            I => \N__41018\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__41018\,
            I => \sAddress_RNI6VH7_6Z0Z_1\
        );

    \I__8642\ : CascadeMux
    port map (
            O => \N__41015\,
            I => \sAddress_RNI6VH7_6Z0Z_1_cascade_\
        );

    \I__8641\ : CascadeMux
    port map (
            O => \N__41012\,
            I => \N__41007\
        );

    \I__8640\ : CascadeMux
    port map (
            O => \N__41011\,
            I => \N__41004\
        );

    \I__8639\ : CascadeMux
    port map (
            O => \N__41010\,
            I => \N__41001\
        );

    \I__8638\ : InMux
    port map (
            O => \N__41007\,
            I => \N__40991\
        );

    \I__8637\ : InMux
    port map (
            O => \N__41004\,
            I => \N__40986\
        );

    \I__8636\ : InMux
    port map (
            O => \N__41001\,
            I => \N__40986\
        );

    \I__8635\ : CascadeMux
    port map (
            O => \N__41000\,
            I => \N__40982\
        );

    \I__8634\ : CascadeMux
    port map (
            O => \N__40999\,
            I => \N__40979\
        );

    \I__8633\ : CascadeMux
    port map (
            O => \N__40998\,
            I => \N__40973\
        );

    \I__8632\ : CascadeMux
    port map (
            O => \N__40997\,
            I => \N__40970\
        );

    \I__8631\ : CascadeMux
    port map (
            O => \N__40996\,
            I => \N__40965\
        );

    \I__8630\ : CascadeMux
    port map (
            O => \N__40995\,
            I => \N__40962\
        );

    \I__8629\ : CascadeMux
    port map (
            O => \N__40994\,
            I => \N__40957\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__40991\,
            I => \N__40951\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__40986\,
            I => \N__40951\
        );

    \I__8626\ : InMux
    port map (
            O => \N__40985\,
            I => \N__40940\
        );

    \I__8625\ : InMux
    port map (
            O => \N__40982\,
            I => \N__40940\
        );

    \I__8624\ : InMux
    port map (
            O => \N__40979\,
            I => \N__40940\
        );

    \I__8623\ : InMux
    port map (
            O => \N__40978\,
            I => \N__40940\
        );

    \I__8622\ : CascadeMux
    port map (
            O => \N__40977\,
            I => \N__40937\
        );

    \I__8621\ : CascadeMux
    port map (
            O => \N__40976\,
            I => \N__40934\
        );

    \I__8620\ : InMux
    port map (
            O => \N__40973\,
            I => \N__40931\
        );

    \I__8619\ : InMux
    port map (
            O => \N__40970\,
            I => \N__40922\
        );

    \I__8618\ : InMux
    port map (
            O => \N__40969\,
            I => \N__40922\
        );

    \I__8617\ : InMux
    port map (
            O => \N__40968\,
            I => \N__40922\
        );

    \I__8616\ : InMux
    port map (
            O => \N__40965\,
            I => \N__40922\
        );

    \I__8615\ : InMux
    port map (
            O => \N__40962\,
            I => \N__40915\
        );

    \I__8614\ : InMux
    port map (
            O => \N__40961\,
            I => \N__40915\
        );

    \I__8613\ : InMux
    port map (
            O => \N__40960\,
            I => \N__40915\
        );

    \I__8612\ : InMux
    port map (
            O => \N__40957\,
            I => \N__40910\
        );

    \I__8611\ : InMux
    port map (
            O => \N__40956\,
            I => \N__40910\
        );

    \I__8610\ : Span4Mux_v
    port map (
            O => \N__40951\,
            I => \N__40907\
        );

    \I__8609\ : InMux
    port map (
            O => \N__40950\,
            I => \N__40904\
        );

    \I__8608\ : InMux
    port map (
            O => \N__40949\,
            I => \N__40901\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__40940\,
            I => \N__40897\
        );

    \I__8606\ : InMux
    port map (
            O => \N__40937\,
            I => \N__40889\
        );

    \I__8605\ : InMux
    port map (
            O => \N__40934\,
            I => \N__40889\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__40931\,
            I => \N__40882\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__40922\,
            I => \N__40882\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__40915\,
            I => \N__40882\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__40910\,
            I => \N__40877\
        );

    \I__8600\ : Span4Mux_v
    port map (
            O => \N__40907\,
            I => \N__40877\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__40904\,
            I => \N__40872\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__40901\,
            I => \N__40872\
        );

    \I__8597\ : CascadeMux
    port map (
            O => \N__40900\,
            I => \N__40868\
        );

    \I__8596\ : Span4Mux_v
    port map (
            O => \N__40897\,
            I => \N__40865\
        );

    \I__8595\ : InMux
    port map (
            O => \N__40896\,
            I => \N__40854\
        );

    \I__8594\ : InMux
    port map (
            O => \N__40895\,
            I => \N__40854\
        );

    \I__8593\ : InMux
    port map (
            O => \N__40894\,
            I => \N__40854\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__40889\,
            I => \N__40851\
        );

    \I__8591\ : Span4Mux_v
    port map (
            O => \N__40882\,
            I => \N__40844\
        );

    \I__8590\ : Span4Mux_h
    port map (
            O => \N__40877\,
            I => \N__40844\
        );

    \I__8589\ : Span4Mux_v
    port map (
            O => \N__40872\,
            I => \N__40844\
        );

    \I__8588\ : InMux
    port map (
            O => \N__40871\,
            I => \N__40839\
        );

    \I__8587\ : InMux
    port map (
            O => \N__40868\,
            I => \N__40839\
        );

    \I__8586\ : Sp12to4
    port map (
            O => \N__40865\,
            I => \N__40836\
        );

    \I__8585\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40829\
        );

    \I__8584\ : InMux
    port map (
            O => \N__40863\,
            I => \N__40829\
        );

    \I__8583\ : InMux
    port map (
            O => \N__40862\,
            I => \N__40829\
        );

    \I__8582\ : InMux
    port map (
            O => \N__40861\,
            I => \N__40826\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__40854\,
            I => \sAddressZ0Z_5\
        );

    \I__8580\ : Odrv4
    port map (
            O => \N__40851\,
            I => \sAddressZ0Z_5\
        );

    \I__8579\ : Odrv4
    port map (
            O => \N__40844\,
            I => \sAddressZ0Z_5\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__40839\,
            I => \sAddressZ0Z_5\
        );

    \I__8577\ : Odrv12
    port map (
            O => \N__40836\,
            I => \sAddressZ0Z_5\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__40829\,
            I => \sAddressZ0Z_5\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__40826\,
            I => \sAddressZ0Z_5\
        );

    \I__8574\ : InMux
    port map (
            O => \N__40811\,
            I => \N__40806\
        );

    \I__8573\ : InMux
    port map (
            O => \N__40810\,
            I => \N__40801\
        );

    \I__8572\ : InMux
    port map (
            O => \N__40809\,
            I => \N__40801\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__40806\,
            I => \N__40790\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__40801\,
            I => \N__40787\
        );

    \I__8569\ : InMux
    port map (
            O => \N__40800\,
            I => \N__40775\
        );

    \I__8568\ : InMux
    port map (
            O => \N__40799\,
            I => \N__40775\
        );

    \I__8567\ : InMux
    port map (
            O => \N__40798\,
            I => \N__40775\
        );

    \I__8566\ : InMux
    port map (
            O => \N__40797\,
            I => \N__40775\
        );

    \I__8565\ : InMux
    port map (
            O => \N__40796\,
            I => \N__40766\
        );

    \I__8564\ : InMux
    port map (
            O => \N__40795\,
            I => \N__40766\
        );

    \I__8563\ : InMux
    port map (
            O => \N__40794\,
            I => \N__40766\
        );

    \I__8562\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40766\
        );

    \I__8561\ : Span4Mux_v
    port map (
            O => \N__40790\,
            I => \N__40761\
        );

    \I__8560\ : Span4Mux_v
    port map (
            O => \N__40787\,
            I => \N__40761\
        );

    \I__8559\ : InMux
    port map (
            O => \N__40786\,
            I => \N__40754\
        );

    \I__8558\ : InMux
    port map (
            O => \N__40785\,
            I => \N__40754\
        );

    \I__8557\ : InMux
    port map (
            O => \N__40784\,
            I => \N__40754\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__40775\,
            I => \N__40748\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__40766\,
            I => \N__40733\
        );

    \I__8554\ : Span4Mux_h
    port map (
            O => \N__40761\,
            I => \N__40733\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__40754\,
            I => \N__40733\
        );

    \I__8552\ : InMux
    port map (
            O => \N__40753\,
            I => \N__40726\
        );

    \I__8551\ : InMux
    port map (
            O => \N__40752\,
            I => \N__40726\
        );

    \I__8550\ : InMux
    port map (
            O => \N__40751\,
            I => \N__40726\
        );

    \I__8549\ : Span4Mux_v
    port map (
            O => \N__40748\,
            I => \N__40723\
        );

    \I__8548\ : InMux
    port map (
            O => \N__40747\,
            I => \N__40720\
        );

    \I__8547\ : InMux
    port map (
            O => \N__40746\,
            I => \N__40715\
        );

    \I__8546\ : InMux
    port map (
            O => \N__40745\,
            I => \N__40715\
        );

    \I__8545\ : InMux
    port map (
            O => \N__40744\,
            I => \N__40708\
        );

    \I__8544\ : InMux
    port map (
            O => \N__40743\,
            I => \N__40708\
        );

    \I__8543\ : InMux
    port map (
            O => \N__40742\,
            I => \N__40708\
        );

    \I__8542\ : InMux
    port map (
            O => \N__40741\,
            I => \N__40705\
        );

    \I__8541\ : InMux
    port map (
            O => \N__40740\,
            I => \N__40702\
        );

    \I__8540\ : Span4Mux_v
    port map (
            O => \N__40733\,
            I => \N__40699\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__40726\,
            I => \N__40696\
        );

    \I__8538\ : Sp12to4
    port map (
            O => \N__40723\,
            I => \N__40693\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__40720\,
            I => \sAddress_RNIP2UK1Z0Z_4\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__40715\,
            I => \sAddress_RNIP2UK1Z0Z_4\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__40708\,
            I => \sAddress_RNIP2UK1Z0Z_4\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__40705\,
            I => \sAddress_RNIP2UK1Z0Z_4\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__40702\,
            I => \sAddress_RNIP2UK1Z0Z_4\
        );

    \I__8532\ : Odrv4
    port map (
            O => \N__40699\,
            I => \sAddress_RNIP2UK1Z0Z_4\
        );

    \I__8531\ : Odrv4
    port map (
            O => \N__40696\,
            I => \sAddress_RNIP2UK1Z0Z_4\
        );

    \I__8530\ : Odrv12
    port map (
            O => \N__40693\,
            I => \sAddress_RNIP2UK1Z0Z_4\
        );

    \I__8529\ : CascadeMux
    port map (
            O => \N__40676\,
            I => \N__40670\
        );

    \I__8528\ : InMux
    port map (
            O => \N__40675\,
            I => \N__40660\
        );

    \I__8527\ : InMux
    port map (
            O => \N__40674\,
            I => \N__40660\
        );

    \I__8526\ : InMux
    port map (
            O => \N__40673\,
            I => \N__40660\
        );

    \I__8525\ : InMux
    port map (
            O => \N__40670\,
            I => \N__40660\
        );

    \I__8524\ : CascadeMux
    port map (
            O => \N__40669\,
            I => \N__40655\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__40660\,
            I => \N__40648\
        );

    \I__8522\ : InMux
    port map (
            O => \N__40659\,
            I => \N__40642\
        );

    \I__8521\ : InMux
    port map (
            O => \N__40658\,
            I => \N__40633\
        );

    \I__8520\ : InMux
    port map (
            O => \N__40655\,
            I => \N__40633\
        );

    \I__8519\ : InMux
    port map (
            O => \N__40654\,
            I => \N__40633\
        );

    \I__8518\ : InMux
    port map (
            O => \N__40653\,
            I => \N__40633\
        );

    \I__8517\ : InMux
    port map (
            O => \N__40652\,
            I => \N__40627\
        );

    \I__8516\ : InMux
    port map (
            O => \N__40651\,
            I => \N__40627\
        );

    \I__8515\ : Span4Mux_v
    port map (
            O => \N__40648\,
            I => \N__40624\
        );

    \I__8514\ : InMux
    port map (
            O => \N__40647\,
            I => \N__40621\
        );

    \I__8513\ : InMux
    port map (
            O => \N__40646\,
            I => \N__40610\
        );

    \I__8512\ : InMux
    port map (
            O => \N__40645\,
            I => \N__40610\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__40642\,
            I => \N__40605\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__40633\,
            I => \N__40605\
        );

    \I__8509\ : InMux
    port map (
            O => \N__40632\,
            I => \N__40600\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__40627\,
            I => \N__40597\
        );

    \I__8507\ : Span4Mux_h
    port map (
            O => \N__40624\,
            I => \N__40592\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__40621\,
            I => \N__40592\
        );

    \I__8505\ : InMux
    port map (
            O => \N__40620\,
            I => \N__40589\
        );

    \I__8504\ : InMux
    port map (
            O => \N__40619\,
            I => \N__40580\
        );

    \I__8503\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40580\
        );

    \I__8502\ : InMux
    port map (
            O => \N__40617\,
            I => \N__40580\
        );

    \I__8501\ : InMux
    port map (
            O => \N__40616\,
            I => \N__40580\
        );

    \I__8500\ : InMux
    port map (
            O => \N__40615\,
            I => \N__40577\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__40610\,
            I => \N__40572\
        );

    \I__8498\ : Span12Mux_h
    port map (
            O => \N__40605\,
            I => \N__40572\
        );

    \I__8497\ : InMux
    port map (
            O => \N__40604\,
            I => \N__40567\
        );

    \I__8496\ : InMux
    port map (
            O => \N__40603\,
            I => \N__40567\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__40600\,
            I => \N__40562\
        );

    \I__8494\ : Sp12to4
    port map (
            O => \N__40597\,
            I => \N__40562\
        );

    \I__8493\ : Odrv4
    port map (
            O => \N__40592\,
            I => \sAddressZ0Z_2\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__40589\,
            I => \sAddressZ0Z_2\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__40580\,
            I => \sAddressZ0Z_2\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__40577\,
            I => \sAddressZ0Z_2\
        );

    \I__8489\ : Odrv12
    port map (
            O => \N__40572\,
            I => \sAddressZ0Z_2\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__40567\,
            I => \sAddressZ0Z_2\
        );

    \I__8487\ : Odrv12
    port map (
            O => \N__40562\,
            I => \sAddressZ0Z_2\
        );

    \I__8486\ : InMux
    port map (
            O => \N__40547\,
            I => \N__40540\
        );

    \I__8485\ : InMux
    port map (
            O => \N__40546\,
            I => \N__40540\
        );

    \I__8484\ : InMux
    port map (
            O => \N__40545\,
            I => \N__40537\
        );

    \I__8483\ : LocalMux
    port map (
            O => \N__40540\,
            I => \N__40534\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__40537\,
            I => \N__40528\
        );

    \I__8481\ : Span4Mux_h
    port map (
            O => \N__40534\,
            I => \N__40525\
        );

    \I__8480\ : InMux
    port map (
            O => \N__40533\,
            I => \N__40522\
        );

    \I__8479\ : CascadeMux
    port map (
            O => \N__40532\,
            I => \N__40517\
        );

    \I__8478\ : CascadeMux
    port map (
            O => \N__40531\,
            I => \N__40513\
        );

    \I__8477\ : Span4Mux_h
    port map (
            O => \N__40528\,
            I => \N__40510\
        );

    \I__8476\ : Span4Mux_h
    port map (
            O => \N__40525\,
            I => \N__40504\
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__40522\,
            I => \N__40501\
        );

    \I__8474\ : CascadeMux
    port map (
            O => \N__40521\,
            I => \N__40497\
        );

    \I__8473\ : InMux
    port map (
            O => \N__40520\,
            I => \N__40493\
        );

    \I__8472\ : InMux
    port map (
            O => \N__40517\,
            I => \N__40488\
        );

    \I__8471\ : InMux
    port map (
            O => \N__40516\,
            I => \N__40488\
        );

    \I__8470\ : InMux
    port map (
            O => \N__40513\,
            I => \N__40485\
        );

    \I__8469\ : Span4Mux_v
    port map (
            O => \N__40510\,
            I => \N__40482\
        );

    \I__8468\ : InMux
    port map (
            O => \N__40509\,
            I => \N__40479\
        );

    \I__8467\ : InMux
    port map (
            O => \N__40508\,
            I => \N__40474\
        );

    \I__8466\ : InMux
    port map (
            O => \N__40507\,
            I => \N__40474\
        );

    \I__8465\ : Span4Mux_h
    port map (
            O => \N__40504\,
            I => \N__40469\
        );

    \I__8464\ : Span4Mux_h
    port map (
            O => \N__40501\,
            I => \N__40469\
        );

    \I__8463\ : InMux
    port map (
            O => \N__40500\,
            I => \N__40466\
        );

    \I__8462\ : InMux
    port map (
            O => \N__40497\,
            I => \N__40461\
        );

    \I__8461\ : InMux
    port map (
            O => \N__40496\,
            I => \N__40461\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__40493\,
            I => \N__40456\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__40488\,
            I => \N__40456\
        );

    \I__8458\ : LocalMux
    port map (
            O => \N__40485\,
            I => \sAddressZ0Z_1\
        );

    \I__8457\ : Odrv4
    port map (
            O => \N__40482\,
            I => \sAddressZ0Z_1\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__40479\,
            I => \sAddressZ0Z_1\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__40474\,
            I => \sAddressZ0Z_1\
        );

    \I__8454\ : Odrv4
    port map (
            O => \N__40469\,
            I => \sAddressZ0Z_1\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__40466\,
            I => \sAddressZ0Z_1\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__40461\,
            I => \sAddressZ0Z_1\
        );

    \I__8451\ : Odrv12
    port map (
            O => \N__40456\,
            I => \sAddressZ0Z_1\
        );

    \I__8450\ : CascadeMux
    port map (
            O => \N__40439\,
            I => \N__40434\
        );

    \I__8449\ : CascadeMux
    port map (
            O => \N__40438\,
            I => \N__40430\
        );

    \I__8448\ : InMux
    port map (
            O => \N__40437\,
            I => \N__40419\
        );

    \I__8447\ : InMux
    port map (
            O => \N__40434\,
            I => \N__40419\
        );

    \I__8446\ : InMux
    port map (
            O => \N__40433\,
            I => \N__40419\
        );

    \I__8445\ : InMux
    port map (
            O => \N__40430\,
            I => \N__40419\
        );

    \I__8444\ : CascadeMux
    port map (
            O => \N__40429\,
            I => \N__40413\
        );

    \I__8443\ : InMux
    port map (
            O => \N__40428\,
            I => \N__40399\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__40419\,
            I => \N__40396\
        );

    \I__8441\ : InMux
    port map (
            O => \N__40418\,
            I => \N__40391\
        );

    \I__8440\ : InMux
    port map (
            O => \N__40417\,
            I => \N__40391\
        );

    \I__8439\ : InMux
    port map (
            O => \N__40416\,
            I => \N__40386\
        );

    \I__8438\ : InMux
    port map (
            O => \N__40413\,
            I => \N__40386\
        );

    \I__8437\ : CascadeMux
    port map (
            O => \N__40412\,
            I => \N__40381\
        );

    \I__8436\ : CascadeMux
    port map (
            O => \N__40411\,
            I => \N__40378\
        );

    \I__8435\ : InMux
    port map (
            O => \N__40410\,
            I => \N__40374\
        );

    \I__8434\ : InMux
    port map (
            O => \N__40409\,
            I => \N__40367\
        );

    \I__8433\ : InMux
    port map (
            O => \N__40408\,
            I => \N__40367\
        );

    \I__8432\ : InMux
    port map (
            O => \N__40407\,
            I => \N__40367\
        );

    \I__8431\ : InMux
    port map (
            O => \N__40406\,
            I => \N__40364\
        );

    \I__8430\ : InMux
    port map (
            O => \N__40405\,
            I => \N__40357\
        );

    \I__8429\ : InMux
    port map (
            O => \N__40404\,
            I => \N__40357\
        );

    \I__8428\ : InMux
    port map (
            O => \N__40403\,
            I => \N__40357\
        );

    \I__8427\ : InMux
    port map (
            O => \N__40402\,
            I => \N__40354\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__40399\,
            I => \N__40351\
        );

    \I__8425\ : Span4Mux_v
    port map (
            O => \N__40396\,
            I => \N__40348\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__40391\,
            I => \N__40343\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__40386\,
            I => \N__40343\
        );

    \I__8422\ : InMux
    port map (
            O => \N__40385\,
            I => \N__40340\
        );

    \I__8421\ : InMux
    port map (
            O => \N__40384\,
            I => \N__40337\
        );

    \I__8420\ : InMux
    port map (
            O => \N__40381\,
            I => \N__40329\
        );

    \I__8419\ : InMux
    port map (
            O => \N__40378\,
            I => \N__40329\
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__40377\,
            I => \N__40326\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__40374\,
            I => \N__40315\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__40367\,
            I => \N__40315\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__40364\,
            I => \N__40315\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__40357\,
            I => \N__40315\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__40354\,
            I => \N__40315\
        );

    \I__8412\ : Span4Mux_v
    port map (
            O => \N__40351\,
            I => \N__40308\
        );

    \I__8411\ : Span4Mux_v
    port map (
            O => \N__40348\,
            I => \N__40308\
        );

    \I__8410\ : Span4Mux_h
    port map (
            O => \N__40343\,
            I => \N__40308\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__40340\,
            I => \N__40289\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__40337\,
            I => \N__40289\
        );

    \I__8407\ : InMux
    port map (
            O => \N__40336\,
            I => \N__40286\
        );

    \I__8406\ : InMux
    port map (
            O => \N__40335\,
            I => \N__40281\
        );

    \I__8405\ : InMux
    port map (
            O => \N__40334\,
            I => \N__40281\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__40329\,
            I => \N__40278\
        );

    \I__8403\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40275\
        );

    \I__8402\ : Span4Mux_v
    port map (
            O => \N__40315\,
            I => \N__40270\
        );

    \I__8401\ : Span4Mux_h
    port map (
            O => \N__40308\,
            I => \N__40270\
        );

    \I__8400\ : InMux
    port map (
            O => \N__40307\,
            I => \N__40264\
        );

    \I__8399\ : InMux
    port map (
            O => \N__40306\,
            I => \N__40264\
        );

    \I__8398\ : InMux
    port map (
            O => \N__40305\,
            I => \N__40255\
        );

    \I__8397\ : InMux
    port map (
            O => \N__40304\,
            I => \N__40255\
        );

    \I__8396\ : InMux
    port map (
            O => \N__40303\,
            I => \N__40255\
        );

    \I__8395\ : InMux
    port map (
            O => \N__40302\,
            I => \N__40255\
        );

    \I__8394\ : InMux
    port map (
            O => \N__40301\,
            I => \N__40252\
        );

    \I__8393\ : InMux
    port map (
            O => \N__40300\,
            I => \N__40241\
        );

    \I__8392\ : InMux
    port map (
            O => \N__40299\,
            I => \N__40241\
        );

    \I__8391\ : InMux
    port map (
            O => \N__40298\,
            I => \N__40241\
        );

    \I__8390\ : InMux
    port map (
            O => \N__40297\,
            I => \N__40241\
        );

    \I__8389\ : InMux
    port map (
            O => \N__40296\,
            I => \N__40241\
        );

    \I__8388\ : InMux
    port map (
            O => \N__40295\,
            I => \N__40236\
        );

    \I__8387\ : InMux
    port map (
            O => \N__40294\,
            I => \N__40236\
        );

    \I__8386\ : Span4Mux_v
    port map (
            O => \N__40289\,
            I => \N__40233\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__40286\,
            I => \N__40224\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__40281\,
            I => \N__40224\
        );

    \I__8383\ : Span4Mux_v
    port map (
            O => \N__40278\,
            I => \N__40224\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__40275\,
            I => \N__40224\
        );

    \I__8381\ : Span4Mux_h
    port map (
            O => \N__40270\,
            I => \N__40221\
        );

    \I__8380\ : InMux
    port map (
            O => \N__40269\,
            I => \N__40218\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__40264\,
            I => \sAddressZ0Z_3\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__40255\,
            I => \sAddressZ0Z_3\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__40252\,
            I => \sAddressZ0Z_3\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__40241\,
            I => \sAddressZ0Z_3\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__40236\,
            I => \sAddressZ0Z_3\
        );

    \I__8374\ : Odrv4
    port map (
            O => \N__40233\,
            I => \sAddressZ0Z_3\
        );

    \I__8373\ : Odrv4
    port map (
            O => \N__40224\,
            I => \sAddressZ0Z_3\
        );

    \I__8372\ : Odrv4
    port map (
            O => \N__40221\,
            I => \sAddressZ0Z_3\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__40218\,
            I => \sAddressZ0Z_3\
        );

    \I__8370\ : CascadeMux
    port map (
            O => \N__40199\,
            I => \N__40192\
        );

    \I__8369\ : CascadeMux
    port map (
            O => \N__40198\,
            I => \N__40186\
        );

    \I__8368\ : InMux
    port map (
            O => \N__40197\,
            I => \N__40181\
        );

    \I__8367\ : InMux
    port map (
            O => \N__40196\,
            I => \N__40181\
        );

    \I__8366\ : CascadeMux
    port map (
            O => \N__40195\,
            I => \N__40177\
        );

    \I__8365\ : InMux
    port map (
            O => \N__40192\,
            I => \N__40164\
        );

    \I__8364\ : InMux
    port map (
            O => \N__40191\,
            I => \N__40164\
        );

    \I__8363\ : InMux
    port map (
            O => \N__40190\,
            I => \N__40164\
        );

    \I__8362\ : InMux
    port map (
            O => \N__40189\,
            I => \N__40164\
        );

    \I__8361\ : InMux
    port map (
            O => \N__40186\,
            I => \N__40164\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__40181\,
            I => \N__40154\
        );

    \I__8359\ : InMux
    port map (
            O => \N__40180\,
            I => \N__40151\
        );

    \I__8358\ : InMux
    port map (
            O => \N__40177\,
            I => \N__40148\
        );

    \I__8357\ : InMux
    port map (
            O => \N__40176\,
            I => \N__40143\
        );

    \I__8356\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40143\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__40164\,
            I => \N__40140\
        );

    \I__8354\ : InMux
    port map (
            O => \N__40163\,
            I => \N__40134\
        );

    \I__8353\ : InMux
    port map (
            O => \N__40162\,
            I => \N__40134\
        );

    \I__8352\ : InMux
    port map (
            O => \N__40161\,
            I => \N__40129\
        );

    \I__8351\ : InMux
    port map (
            O => \N__40160\,
            I => \N__40129\
        );

    \I__8350\ : InMux
    port map (
            O => \N__40159\,
            I => \N__40124\
        );

    \I__8349\ : InMux
    port map (
            O => \N__40158\,
            I => \N__40124\
        );

    \I__8348\ : CascadeMux
    port map (
            O => \N__40157\,
            I => \N__40121\
        );

    \I__8347\ : Span4Mux_v
    port map (
            O => \N__40154\,
            I => \N__40117\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__40151\,
            I => \N__40110\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__40148\,
            I => \N__40110\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__40143\,
            I => \N__40110\
        );

    \I__8343\ : Span4Mux_v
    port map (
            O => \N__40140\,
            I => \N__40107\
        );

    \I__8342\ : InMux
    port map (
            O => \N__40139\,
            I => \N__40104\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__40134\,
            I => \N__40097\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__40129\,
            I => \N__40097\
        );

    \I__8339\ : LocalMux
    port map (
            O => \N__40124\,
            I => \N__40097\
        );

    \I__8338\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40092\
        );

    \I__8337\ : InMux
    port map (
            O => \N__40120\,
            I => \N__40092\
        );

    \I__8336\ : Sp12to4
    port map (
            O => \N__40117\,
            I => \N__40089\
        );

    \I__8335\ : Span4Mux_v
    port map (
            O => \N__40110\,
            I => \N__40084\
        );

    \I__8334\ : Span4Mux_v
    port map (
            O => \N__40107\,
            I => \N__40084\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__40104\,
            I => \sAddressZ0Z_0\
        );

    \I__8332\ : Odrv12
    port map (
            O => \N__40097\,
            I => \sAddressZ0Z_0\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__40092\,
            I => \sAddressZ0Z_0\
        );

    \I__8330\ : Odrv12
    port map (
            O => \N__40089\,
            I => \sAddressZ0Z_0\
        );

    \I__8329\ : Odrv4
    port map (
            O => \N__40084\,
            I => \sAddressZ0Z_0\
        );

    \I__8328\ : InMux
    port map (
            O => \N__40073\,
            I => \N__40069\
        );

    \I__8327\ : InMux
    port map (
            O => \N__40072\,
            I => \N__40066\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__40069\,
            I => \N__40063\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__40066\,
            I => \N__40060\
        );

    \I__8324\ : Span4Mux_v
    port map (
            O => \N__40063\,
            I => \N__40057\
        );

    \I__8323\ : Span4Mux_h
    port map (
            O => \N__40060\,
            I => \N__40054\
        );

    \I__8322\ : Span4Mux_h
    port map (
            O => \N__40057\,
            I => \N__40049\
        );

    \I__8321\ : Span4Mux_v
    port map (
            O => \N__40054\,
            I => \N__40046\
        );

    \I__8320\ : InMux
    port map (
            O => \N__40053\,
            I => \N__40041\
        );

    \I__8319\ : InMux
    port map (
            O => \N__40052\,
            I => \N__40041\
        );

    \I__8318\ : Span4Mux_h
    port map (
            O => \N__40049\,
            I => \N__40034\
        );

    \I__8317\ : Span4Mux_v
    port map (
            O => \N__40046\,
            I => \N__40034\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__40041\,
            I => \N__40034\
        );

    \I__8315\ : Odrv4
    port map (
            O => \N__40034\,
            I => \sAddress_RNIAM2A_1Z0Z_1\
        );

    \I__8314\ : CascadeMux
    port map (
            O => \N__40031\,
            I => \sAddress_RNIAM2A_1Z0Z_1_cascade_\
        );

    \I__8313\ : InMux
    port map (
            O => \N__40028\,
            I => \N__40021\
        );

    \I__8312\ : InMux
    port map (
            O => \N__40027\,
            I => \N__40016\
        );

    \I__8311\ : InMux
    port map (
            O => \N__40026\,
            I => \N__40016\
        );

    \I__8310\ : InMux
    port map (
            O => \N__40025\,
            I => \N__40011\
        );

    \I__8309\ : InMux
    port map (
            O => \N__40024\,
            I => \N__40011\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__40021\,
            I => \N__40006\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__40016\,
            I => \N__40003\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__40011\,
            I => \N__39999\
        );

    \I__8305\ : InMux
    port map (
            O => \N__40010\,
            I => \N__39992\
        );

    \I__8304\ : InMux
    port map (
            O => \N__40009\,
            I => \N__39992\
        );

    \I__8303\ : Span4Mux_v
    port map (
            O => \N__40006\,
            I => \N__39988\
        );

    \I__8302\ : Span4Mux_v
    port map (
            O => \N__40003\,
            I => \N__39985\
        );

    \I__8301\ : InMux
    port map (
            O => \N__40002\,
            I => \N__39982\
        );

    \I__8300\ : Span4Mux_v
    port map (
            O => \N__39999\,
            I => \N__39979\
        );

    \I__8299\ : InMux
    port map (
            O => \N__39998\,
            I => \N__39974\
        );

    \I__8298\ : InMux
    port map (
            O => \N__39997\,
            I => \N__39974\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__39992\,
            I => \N__39966\
        );

    \I__8296\ : InMux
    port map (
            O => \N__39991\,
            I => \N__39963\
        );

    \I__8295\ : Sp12to4
    port map (
            O => \N__39988\,
            I => \N__39958\
        );

    \I__8294\ : Sp12to4
    port map (
            O => \N__39985\,
            I => \N__39958\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__39982\,
            I => \N__39951\
        );

    \I__8292\ : Span4Mux_h
    port map (
            O => \N__39979\,
            I => \N__39951\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__39974\,
            I => \N__39951\
        );

    \I__8290\ : InMux
    port map (
            O => \N__39973\,
            I => \N__39948\
        );

    \I__8289\ : InMux
    port map (
            O => \N__39972\,
            I => \N__39945\
        );

    \I__8288\ : InMux
    port map (
            O => \N__39971\,
            I => \N__39940\
        );

    \I__8287\ : InMux
    port map (
            O => \N__39970\,
            I => \N__39940\
        );

    \I__8286\ : InMux
    port map (
            O => \N__39969\,
            I => \N__39937\
        );

    \I__8285\ : Odrv4
    port map (
            O => \N__39966\,
            I => \sAddress_RNIVREN1Z0Z_4\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__39963\,
            I => \sAddress_RNIVREN1Z0Z_4\
        );

    \I__8283\ : Odrv12
    port map (
            O => \N__39958\,
            I => \sAddress_RNIVREN1Z0Z_4\
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__39951\,
            I => \sAddress_RNIVREN1Z0Z_4\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__39948\,
            I => \sAddress_RNIVREN1Z0Z_4\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__39945\,
            I => \sAddress_RNIVREN1Z0Z_4\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__39940\,
            I => \sAddress_RNIVREN1Z0Z_4\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__39937\,
            I => \sAddress_RNIVREN1Z0Z_4\
        );

    \I__8277\ : CEMux
    port map (
            O => \N__39920\,
            I => \N__39917\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__39917\,
            I => \N__39914\
        );

    \I__8275\ : Sp12to4
    port map (
            O => \N__39914\,
            I => \N__39911\
        );

    \I__8274\ : Odrv12
    port map (
            O => \N__39911\,
            I => \sDAC_mem_17_1_sqmuxa\
        );

    \I__8273\ : InMux
    port map (
            O => \N__39908\,
            I => \N__39905\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__39905\,
            I => \N__39902\
        );

    \I__8271\ : Span4Mux_v
    port map (
            O => \N__39902\,
            I => \N__39899\
        );

    \I__8270\ : Odrv4
    port map (
            O => \N__39899\,
            I => \sDAC_mem_41Z0Z_0\
        );

    \I__8269\ : InMux
    port map (
            O => \N__39896\,
            I => \N__39893\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__39893\,
            I => \N__39890\
        );

    \I__8267\ : Span12Mux_v
    port map (
            O => \N__39890\,
            I => \N__39887\
        );

    \I__8266\ : Odrv12
    port map (
            O => \N__39887\,
            I => \sDAC_mem_41Z0Z_1\
        );

    \I__8265\ : InMux
    port map (
            O => \N__39884\,
            I => \N__39881\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__39881\,
            I => \N__39878\
        );

    \I__8263\ : Span4Mux_v
    port map (
            O => \N__39878\,
            I => \N__39875\
        );

    \I__8262\ : Odrv4
    port map (
            O => \N__39875\,
            I => \sDAC_mem_41Z0Z_2\
        );

    \I__8261\ : InMux
    port map (
            O => \N__39872\,
            I => \N__39869\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__39869\,
            I => \N__39866\
        );

    \I__8259\ : Span4Mux_v
    port map (
            O => \N__39866\,
            I => \N__39863\
        );

    \I__8258\ : Span4Mux_h
    port map (
            O => \N__39863\,
            I => \N__39860\
        );

    \I__8257\ : Odrv4
    port map (
            O => \N__39860\,
            I => \sDAC_mem_41Z0Z_3\
        );

    \I__8256\ : InMux
    port map (
            O => \N__39857\,
            I => \N__39854\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__39854\,
            I => \N__39851\
        );

    \I__8254\ : Span4Mux_h
    port map (
            O => \N__39851\,
            I => \N__39848\
        );

    \I__8253\ : Span4Mux_h
    port map (
            O => \N__39848\,
            I => \N__39845\
        );

    \I__8252\ : Odrv4
    port map (
            O => \N__39845\,
            I => \sDAC_mem_41Z0Z_5\
        );

    \I__8251\ : InMux
    port map (
            O => \N__39842\,
            I => \N__39839\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__39839\,
            I => \N__39836\
        );

    \I__8249\ : Span4Mux_h
    port map (
            O => \N__39836\,
            I => \N__39833\
        );

    \I__8248\ : Odrv4
    port map (
            O => \N__39833\,
            I => \sDAC_mem_41Z0Z_6\
        );

    \I__8247\ : InMux
    port map (
            O => \N__39830\,
            I => \N__39827\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__39827\,
            I => \N__39824\
        );

    \I__8245\ : Span4Mux_v
    port map (
            O => \N__39824\,
            I => \N__39821\
        );

    \I__8244\ : Odrv4
    port map (
            O => \N__39821\,
            I => \sDAC_mem_41Z0Z_7\
        );

    \I__8243\ : CEMux
    port map (
            O => \N__39818\,
            I => \N__39815\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__39815\,
            I => \N__39812\
        );

    \I__8241\ : Span4Mux_v
    port map (
            O => \N__39812\,
            I => \N__39809\
        );

    \I__8240\ : Odrv4
    port map (
            O => \N__39809\,
            I => \sDAC_mem_9_1_sqmuxa\
        );

    \I__8239\ : CEMux
    port map (
            O => \N__39806\,
            I => \N__39803\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__39803\,
            I => \N__39799\
        );

    \I__8237\ : CEMux
    port map (
            O => \N__39802\,
            I => \N__39796\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__39799\,
            I => \N__39791\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__39796\,
            I => \N__39791\
        );

    \I__8234\ : Span4Mux_v
    port map (
            O => \N__39791\,
            I => \N__39788\
        );

    \I__8233\ : Odrv4
    port map (
            O => \N__39788\,
            I => \sDAC_mem_41_1_sqmuxa\
        );

    \I__8232\ : IoInMux
    port map (
            O => \N__39785\,
            I => \N__39782\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__39782\,
            I => \N__39779\
        );

    \I__8230\ : IoSpan4Mux
    port map (
            O => \N__39779\,
            I => \N__39776\
        );

    \I__8229\ : Span4Mux_s3_v
    port map (
            O => \N__39776\,
            I => \N__39773\
        );

    \I__8228\ : Span4Mux_h
    port map (
            O => \N__39773\,
            I => \N__39769\
        );

    \I__8227\ : CascadeMux
    port map (
            O => \N__39772\,
            I => \N__39766\
        );

    \I__8226\ : Span4Mux_v
    port map (
            O => \N__39769\,
            I => \N__39763\
        );

    \I__8225\ : InMux
    port map (
            O => \N__39766\,
            I => \N__39760\
        );

    \I__8224\ : Odrv4
    port map (
            O => \N__39763\,
            I => \RAM_DATA_cl_8Z0Z_15\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__39760\,
            I => \RAM_DATA_cl_8Z0Z_15\
        );

    \I__8222\ : IoInMux
    port map (
            O => \N__39755\,
            I => \N__39752\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__39752\,
            I => \N__39749\
        );

    \I__8220\ : Span4Mux_s3_v
    port map (
            O => \N__39749\,
            I => \N__39746\
        );

    \I__8219\ : Span4Mux_h
    port map (
            O => \N__39746\,
            I => \N__39743\
        );

    \I__8218\ : Span4Mux_h
    port map (
            O => \N__39743\,
            I => \N__39739\
        );

    \I__8217\ : CascadeMux
    port map (
            O => \N__39742\,
            I => \N__39736\
        );

    \I__8216\ : Span4Mux_v
    port map (
            O => \N__39739\,
            I => \N__39733\
        );

    \I__8215\ : InMux
    port map (
            O => \N__39736\,
            I => \N__39730\
        );

    \I__8214\ : Odrv4
    port map (
            O => \N__39733\,
            I => \RAM_DATA_cl_9Z0Z_15\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__39730\,
            I => \RAM_DATA_cl_9Z0Z_15\
        );

    \I__8212\ : IoInMux
    port map (
            O => \N__39725\,
            I => \N__39722\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__39722\,
            I => \N__39719\
        );

    \I__8210\ : Span4Mux_s3_v
    port map (
            O => \N__39719\,
            I => \N__39716\
        );

    \I__8209\ : Span4Mux_h
    port map (
            O => \N__39716\,
            I => \N__39713\
        );

    \I__8208\ : Span4Mux_v
    port map (
            O => \N__39713\,
            I => \N__39709\
        );

    \I__8207\ : InMux
    port map (
            O => \N__39712\,
            I => \N__39706\
        );

    \I__8206\ : Odrv4
    port map (
            O => \N__39709\,
            I => \RAM_DATA_clZ0Z_15\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__39706\,
            I => \RAM_DATA_clZ0Z_15\
        );

    \I__8204\ : IoInMux
    port map (
            O => \N__39701\,
            I => \N__39698\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__39698\,
            I => \N__39695\
        );

    \I__8202\ : IoSpan4Mux
    port map (
            O => \N__39695\,
            I => \N__39692\
        );

    \I__8201\ : IoSpan4Mux
    port map (
            O => \N__39692\,
            I => \N__39689\
        );

    \I__8200\ : IoSpan4Mux
    port map (
            O => \N__39689\,
            I => \N__39686\
        );

    \I__8199\ : Span4Mux_s3_v
    port map (
            O => \N__39686\,
            I => \N__39683\
        );

    \I__8198\ : Odrv4
    port map (
            O => \N__39683\,
            I => \RAM_DATA_1Z0Z_7\
        );

    \I__8197\ : InMux
    port map (
            O => \N__39680\,
            I => \N__39677\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__39677\,
            I => \N__39674\
        );

    \I__8195\ : Span4Mux_h
    port map (
            O => \N__39674\,
            I => \N__39671\
        );

    \I__8194\ : Odrv4
    port map (
            O => \N__39671\,
            I => \sDAC_mem_41Z0Z_4\
        );

    \I__8193\ : InMux
    port map (
            O => \N__39668\,
            I => \N__39665\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__39665\,
            I => \N__39662\
        );

    \I__8191\ : Span4Mux_v
    port map (
            O => \N__39662\,
            I => \N__39659\
        );

    \I__8190\ : Odrv4
    port map (
            O => \N__39659\,
            I => \sDAC_mem_36Z0Z_3\
        );

    \I__8189\ : InMux
    port map (
            O => \N__39656\,
            I => \N__39653\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__39653\,
            I => \N__39650\
        );

    \I__8187\ : Span4Mux_h
    port map (
            O => \N__39650\,
            I => \N__39647\
        );

    \I__8186\ : Odrv4
    port map (
            O => \N__39647\,
            I => \sDAC_mem_4Z0Z_3\
        );

    \I__8185\ : CascadeMux
    port map (
            O => \N__39644\,
            I => \sDAC_data_2_13_am_1_6_cascade_\
        );

    \I__8184\ : InMux
    port map (
            O => \N__39641\,
            I => \N__39638\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__39638\,
            I => \N__39635\
        );

    \I__8182\ : Odrv12
    port map (
            O => \N__39635\,
            I => \sDAC_data_RNO_4Z0Z_6\
        );

    \I__8181\ : InMux
    port map (
            O => \N__39632\,
            I => \N__39629\
        );

    \I__8180\ : LocalMux
    port map (
            O => \N__39629\,
            I => \N__39626\
        );

    \I__8179\ : Odrv4
    port map (
            O => \N__39626\,
            I => \sDAC_mem_32Z0Z_5\
        );

    \I__8178\ : InMux
    port map (
            O => \N__39623\,
            I => \N__39620\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__39620\,
            I => \N__39617\
        );

    \I__8176\ : Span4Mux_h
    port map (
            O => \N__39617\,
            I => \N__39614\
        );

    \I__8175\ : Span4Mux_v
    port map (
            O => \N__39614\,
            I => \N__39611\
        );

    \I__8174\ : Odrv4
    port map (
            O => \N__39611\,
            I => \sDAC_mem_32Z0Z_7\
        );

    \I__8173\ : CascadeMux
    port map (
            O => \N__39608\,
            I => \N__39605\
        );

    \I__8172\ : InMux
    port map (
            O => \N__39605\,
            I => \N__39602\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__39602\,
            I => \N__39598\
        );

    \I__8170\ : InMux
    port map (
            O => \N__39601\,
            I => \N__39595\
        );

    \I__8169\ : Span4Mux_h
    port map (
            O => \N__39598\,
            I => \N__39592\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__39595\,
            I => \sCounterRAMZ0Z_2\
        );

    \I__8167\ : Odrv4
    port map (
            O => \N__39592\,
            I => \sCounterRAMZ0Z_2\
        );

    \I__8166\ : InMux
    port map (
            O => \N__39587\,
            I => \sCounterRAM_cry_1\
        );

    \I__8165\ : InMux
    port map (
            O => \N__39584\,
            I => \N__39580\
        );

    \I__8164\ : InMux
    port map (
            O => \N__39583\,
            I => \N__39577\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__39580\,
            I => \N__39574\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__39577\,
            I => \sCounterRAMZ0Z_3\
        );

    \I__8161\ : Odrv4
    port map (
            O => \N__39574\,
            I => \sCounterRAMZ0Z_3\
        );

    \I__8160\ : InMux
    port map (
            O => \N__39569\,
            I => \sCounterRAM_cry_2\
        );

    \I__8159\ : InMux
    port map (
            O => \N__39566\,
            I => \N__39562\
        );

    \I__8158\ : InMux
    port map (
            O => \N__39565\,
            I => \N__39559\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__39562\,
            I => \N__39556\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__39559\,
            I => \sCounterRAMZ0Z_4\
        );

    \I__8155\ : Odrv4
    port map (
            O => \N__39556\,
            I => \sCounterRAMZ0Z_4\
        );

    \I__8154\ : InMux
    port map (
            O => \N__39551\,
            I => \sCounterRAM_cry_3\
        );

    \I__8153\ : InMux
    port map (
            O => \N__39548\,
            I => \N__39544\
        );

    \I__8152\ : InMux
    port map (
            O => \N__39547\,
            I => \N__39541\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__39544\,
            I => \N__39538\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__39541\,
            I => \sCounterRAMZ0Z_5\
        );

    \I__8149\ : Odrv4
    port map (
            O => \N__39538\,
            I => \sCounterRAMZ0Z_5\
        );

    \I__8148\ : InMux
    port map (
            O => \N__39533\,
            I => \sCounterRAM_cry_4\
        );

    \I__8147\ : InMux
    port map (
            O => \N__39530\,
            I => \N__39526\
        );

    \I__8146\ : InMux
    port map (
            O => \N__39529\,
            I => \N__39523\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__39526\,
            I => \N__39520\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__39523\,
            I => \sCounterRAMZ0Z_6\
        );

    \I__8143\ : Odrv4
    port map (
            O => \N__39520\,
            I => \sCounterRAMZ0Z_6\
        );

    \I__8142\ : InMux
    port map (
            O => \N__39515\,
            I => \sCounterRAM_cry_5\
        );

    \I__8141\ : InMux
    port map (
            O => \N__39512\,
            I => \N__39496\
        );

    \I__8140\ : InMux
    port map (
            O => \N__39511\,
            I => \N__39496\
        );

    \I__8139\ : InMux
    port map (
            O => \N__39510\,
            I => \N__39496\
        );

    \I__8138\ : InMux
    port map (
            O => \N__39509\,
            I => \N__39496\
        );

    \I__8137\ : InMux
    port map (
            O => \N__39508\,
            I => \N__39487\
        );

    \I__8136\ : InMux
    port map (
            O => \N__39507\,
            I => \N__39487\
        );

    \I__8135\ : InMux
    port map (
            O => \N__39506\,
            I => \N__39487\
        );

    \I__8134\ : InMux
    port map (
            O => \N__39505\,
            I => \N__39487\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__39496\,
            I => \N_70_i\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__39487\,
            I => \N_70_i\
        );

    \I__8131\ : InMux
    port map (
            O => \N__39482\,
            I => \sCounterRAM_cry_6\
        );

    \I__8130\ : CascadeMux
    port map (
            O => \N__39479\,
            I => \N__39476\
        );

    \I__8129\ : InMux
    port map (
            O => \N__39476\,
            I => \N__39472\
        );

    \I__8128\ : InMux
    port map (
            O => \N__39475\,
            I => \N__39469\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__39472\,
            I => \N__39466\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__39469\,
            I => \sCounterRAMZ0Z_7\
        );

    \I__8125\ : Odrv4
    port map (
            O => \N__39466\,
            I => \sCounterRAMZ0Z_7\
        );

    \I__8124\ : IoInMux
    port map (
            O => \N__39461\,
            I => \N__39458\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__39458\,
            I => \N__39455\
        );

    \I__8122\ : IoSpan4Mux
    port map (
            O => \N__39455\,
            I => \N__39452\
        );

    \I__8121\ : Span4Mux_s3_h
    port map (
            O => \N__39452\,
            I => \N__39449\
        );

    \I__8120\ : Sp12to4
    port map (
            O => \N__39449\,
            I => \N__39446\
        );

    \I__8119\ : Span12Mux_v
    port map (
            O => \N__39446\,
            I => \N__39442\
        );

    \I__8118\ : CascadeMux
    port map (
            O => \N__39445\,
            I => \N__39439\
        );

    \I__8117\ : Span12Mux_v
    port map (
            O => \N__39442\,
            I => \N__39436\
        );

    \I__8116\ : InMux
    port map (
            O => \N__39439\,
            I => \N__39433\
        );

    \I__8115\ : Odrv12
    port map (
            O => \N__39436\,
            I => \RAM_DATA_cl_6Z0Z_15\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__39433\,
            I => \RAM_DATA_cl_6Z0Z_15\
        );

    \I__8113\ : IoInMux
    port map (
            O => \N__39428\,
            I => \N__39425\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__39425\,
            I => \N__39422\
        );

    \I__8111\ : Span12Mux_s11_h
    port map (
            O => \N__39422\,
            I => \N__39418\
        );

    \I__8110\ : InMux
    port map (
            O => \N__39421\,
            I => \N__39415\
        );

    \I__8109\ : Odrv12
    port map (
            O => \N__39418\,
            I => \RAM_DATA_cl_7Z0Z_15\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__39415\,
            I => \RAM_DATA_cl_7Z0Z_15\
        );

    \I__8107\ : InMux
    port map (
            O => \N__39410\,
            I => \N__39378\
        );

    \I__8106\ : InMux
    port map (
            O => \N__39409\,
            I => \N__39378\
        );

    \I__8105\ : InMux
    port map (
            O => \N__39408\,
            I => \N__39378\
        );

    \I__8104\ : InMux
    port map (
            O => \N__39407\,
            I => \N__39378\
        );

    \I__8103\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39369\
        );

    \I__8102\ : InMux
    port map (
            O => \N__39405\,
            I => \N__39369\
        );

    \I__8101\ : InMux
    port map (
            O => \N__39404\,
            I => \N__39369\
        );

    \I__8100\ : InMux
    port map (
            O => \N__39403\,
            I => \N__39369\
        );

    \I__8099\ : InMux
    port map (
            O => \N__39402\,
            I => \N__39360\
        );

    \I__8098\ : InMux
    port map (
            O => \N__39401\,
            I => \N__39360\
        );

    \I__8097\ : InMux
    port map (
            O => \N__39400\,
            I => \N__39360\
        );

    \I__8096\ : InMux
    port map (
            O => \N__39399\,
            I => \N__39360\
        );

    \I__8095\ : InMux
    port map (
            O => \N__39398\,
            I => \N__39351\
        );

    \I__8094\ : InMux
    port map (
            O => \N__39397\,
            I => \N__39351\
        );

    \I__8093\ : InMux
    port map (
            O => \N__39396\,
            I => \N__39348\
        );

    \I__8092\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39331\
        );

    \I__8091\ : InMux
    port map (
            O => \N__39394\,
            I => \N__39331\
        );

    \I__8090\ : InMux
    port map (
            O => \N__39393\,
            I => \N__39331\
        );

    \I__8089\ : InMux
    port map (
            O => \N__39392\,
            I => \N__39331\
        );

    \I__8088\ : InMux
    port map (
            O => \N__39391\,
            I => \N__39322\
        );

    \I__8087\ : InMux
    port map (
            O => \N__39390\,
            I => \N__39322\
        );

    \I__8086\ : InMux
    port map (
            O => \N__39389\,
            I => \N__39322\
        );

    \I__8085\ : InMux
    port map (
            O => \N__39388\,
            I => \N__39322\
        );

    \I__8084\ : CascadeMux
    port map (
            O => \N__39387\,
            I => \N__39319\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__39378\,
            I => \N__39312\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__39369\,
            I => \N__39312\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__39360\,
            I => \N__39312\
        );

    \I__8080\ : InMux
    port map (
            O => \N__39359\,
            I => \N__39303\
        );

    \I__8079\ : InMux
    port map (
            O => \N__39358\,
            I => \N__39303\
        );

    \I__8078\ : InMux
    port map (
            O => \N__39357\,
            I => \N__39303\
        );

    \I__8077\ : InMux
    port map (
            O => \N__39356\,
            I => \N__39303\
        );

    \I__8076\ : LocalMux
    port map (
            O => \N__39351\,
            I => \N__39298\
        );

    \I__8075\ : LocalMux
    port map (
            O => \N__39348\,
            I => \N__39298\
        );

    \I__8074\ : InMux
    port map (
            O => \N__39347\,
            I => \N__39286\
        );

    \I__8073\ : InMux
    port map (
            O => \N__39346\,
            I => \N__39286\
        );

    \I__8072\ : InMux
    port map (
            O => \N__39345\,
            I => \N__39286\
        );

    \I__8071\ : InMux
    port map (
            O => \N__39344\,
            I => \N__39286\
        );

    \I__8070\ : InMux
    port map (
            O => \N__39343\,
            I => \N__39277\
        );

    \I__8069\ : InMux
    port map (
            O => \N__39342\,
            I => \N__39277\
        );

    \I__8068\ : InMux
    port map (
            O => \N__39341\,
            I => \N__39277\
        );

    \I__8067\ : InMux
    port map (
            O => \N__39340\,
            I => \N__39277\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__39331\,
            I => \N__39272\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__39322\,
            I => \N__39272\
        );

    \I__8064\ : InMux
    port map (
            O => \N__39319\,
            I => \N__39269\
        );

    \I__8063\ : Span4Mux_v
    port map (
            O => \N__39312\,
            I => \N__39262\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__39303\,
            I => \N__39262\
        );

    \I__8061\ : Span4Mux_v
    port map (
            O => \N__39298\,
            I => \N__39262\
        );

    \I__8060\ : InMux
    port map (
            O => \N__39297\,
            I => \N__39257\
        );

    \I__8059\ : InMux
    port map (
            O => \N__39296\,
            I => \N__39257\
        );

    \I__8058\ : InMux
    port map (
            O => \N__39295\,
            I => \N__39254\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__39286\,
            I => \N__39249\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__39277\,
            I => \N__39249\
        );

    \I__8055\ : Span4Mux_h
    port map (
            O => \N__39272\,
            I => \N__39243\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__39269\,
            I => \N__39243\
        );

    \I__8053\ : Span4Mux_h
    port map (
            O => \N__39262\,
            I => \N__39240\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__39257\,
            I => \N__39235\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__39254\,
            I => \N__39235\
        );

    \I__8050\ : Span4Mux_h
    port map (
            O => \N__39249\,
            I => \N__39232\
        );

    \I__8049\ : InMux
    port map (
            O => \N__39248\,
            I => \N__39229\
        );

    \I__8048\ : Span4Mux_v
    port map (
            O => \N__39243\,
            I => \N__39226\
        );

    \I__8047\ : Sp12to4
    port map (
            O => \N__39240\,
            I => \N__39220\
        );

    \I__8046\ : Span12Mux_h
    port map (
            O => \N__39235\,
            I => \N__39220\
        );

    \I__8045\ : Sp12to4
    port map (
            O => \N__39232\,
            I => \N__39215\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__39229\,
            I => \N__39215\
        );

    \I__8043\ : Span4Mux_h
    port map (
            O => \N__39226\,
            I => \N__39212\
        );

    \I__8042\ : InMux
    port map (
            O => \N__39225\,
            I => \N__39209\
        );

    \I__8041\ : Span12Mux_v
    port map (
            O => \N__39220\,
            I => \N__39204\
        );

    \I__8040\ : Span12Mux_v
    port map (
            O => \N__39215\,
            I => \N__39204\
        );

    \I__8039\ : Span4Mux_v
    port map (
            O => \N__39212\,
            I => \N__39201\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__39209\,
            I => \sEEPointerResetZ0\
        );

    \I__8037\ : Odrv12
    port map (
            O => \N__39204\,
            I => \sEEPointerResetZ0\
        );

    \I__8036\ : Odrv4
    port map (
            O => \N__39201\,
            I => \sEEPointerResetZ0\
        );

    \I__8035\ : CascadeMux
    port map (
            O => \N__39194\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3_cascade_\
        );

    \I__8034\ : IoInMux
    port map (
            O => \N__39191\,
            I => \N__39188\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__39188\,
            I => \N__39185\
        );

    \I__8032\ : IoSpan4Mux
    port map (
            O => \N__39185\,
            I => \N__39182\
        );

    \I__8031\ : Span4Mux_s2_v
    port map (
            O => \N__39182\,
            I => \N__39179\
        );

    \I__8030\ : Span4Mux_v
    port map (
            O => \N__39179\,
            I => \N__39176\
        );

    \I__8029\ : Odrv4
    port map (
            O => \N__39176\,
            I => \N_28\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__39173\,
            I => \N__39169\
        );

    \I__8027\ : CascadeMux
    port map (
            O => \N__39172\,
            I => \N__39166\
        );

    \I__8026\ : InMux
    port map (
            O => \N__39169\,
            I => \N__39160\
        );

    \I__8025\ : InMux
    port map (
            O => \N__39166\,
            I => \N__39155\
        );

    \I__8024\ : InMux
    port map (
            O => \N__39165\,
            I => \N__39155\
        );

    \I__8023\ : InMux
    port map (
            O => \N__39164\,
            I => \N__39150\
        );

    \I__8022\ : InMux
    port map (
            O => \N__39163\,
            I => \N__39150\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__39160\,
            I => \N__39145\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__39155\,
            I => \N__39145\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__39150\,
            I => \sSPI_MSB0LSBZ0Z1\
        );

    \I__8018\ : Odrv12
    port map (
            O => \N__39145\,
            I => \sSPI_MSB0LSBZ0Z1\
        );

    \I__8017\ : InMux
    port map (
            O => \N__39140\,
            I => \N__39134\
        );

    \I__8016\ : InMux
    port map (
            O => \N__39139\,
            I => \N__39134\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__39134\,
            I => \N__39131\
        );

    \I__8014\ : Span4Mux_v
    port map (
            O => \N__39131\,
            I => \N__39124\
        );

    \I__8013\ : InMux
    port map (
            O => \N__39130\,
            I => \N__39115\
        );

    \I__8012\ : InMux
    port map (
            O => \N__39129\,
            I => \N__39115\
        );

    \I__8011\ : InMux
    port map (
            O => \N__39128\,
            I => \N__39115\
        );

    \I__8010\ : InMux
    port map (
            O => \N__39127\,
            I => \N__39115\
        );

    \I__8009\ : Span4Mux_v
    port map (
            O => \N__39124\,
            I => \N__39112\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__39115\,
            I => \N__39109\
        );

    \I__8007\ : Sp12to4
    port map (
            O => \N__39112\,
            I => \N__39104\
        );

    \I__8006\ : Span12Mux_v
    port map (
            O => \N__39109\,
            I => \N__39104\
        );

    \I__8005\ : Odrv12
    port map (
            O => \N__39104\,
            I => \spi_mosi_ready_prev3_RNILKERZ0\
        );

    \I__8004\ : IoInMux
    port map (
            O => \N__39101\,
            I => \N__39098\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__39098\,
            I => \N__39095\
        );

    \I__8002\ : IoSpan4Mux
    port map (
            O => \N__39095\,
            I => \N__39092\
        );

    \I__8001\ : IoSpan4Mux
    port map (
            O => \N__39092\,
            I => \N__39089\
        );

    \I__8000\ : Span4Mux_s1_h
    port map (
            O => \N__39089\,
            I => \N__39086\
        );

    \I__7999\ : Sp12to4
    port map (
            O => \N__39086\,
            I => \N__39083\
        );

    \I__7998\ : Span12Mux_v
    port map (
            O => \N__39083\,
            I => \N__39079\
        );

    \I__7997\ : InMux
    port map (
            O => \N__39082\,
            I => \N__39076\
        );

    \I__7996\ : Odrv12
    port map (
            O => \N__39079\,
            I => \RAM_DATA_cl_11Z0Z_15\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__39076\,
            I => \RAM_DATA_cl_11Z0Z_15\
        );

    \I__7994\ : IoInMux
    port map (
            O => \N__39071\,
            I => \N__39068\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__39068\,
            I => \N__39065\
        );

    \I__7992\ : Span4Mux_s2_v
    port map (
            O => \N__39065\,
            I => \N__39062\
        );

    \I__7991\ : Sp12to4
    port map (
            O => \N__39062\,
            I => \N__39059\
        );

    \I__7990\ : Span12Mux_s11_h
    port map (
            O => \N__39059\,
            I => \N__39055\
        );

    \I__7989\ : InMux
    port map (
            O => \N__39058\,
            I => \N__39052\
        );

    \I__7988\ : Odrv12
    port map (
            O => \N__39055\,
            I => \RAM_DATA_cl_12Z0Z_15\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__39052\,
            I => \RAM_DATA_cl_12Z0Z_15\
        );

    \I__7986\ : InMux
    port map (
            O => \N__39047\,
            I => \N__39043\
        );

    \I__7985\ : InMux
    port map (
            O => \N__39046\,
            I => \N__39040\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__39043\,
            I => \N__39037\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__39040\,
            I => \sCounterRAMZ0Z_0\
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__39037\,
            I => \sCounterRAMZ0Z_0\
        );

    \I__7981\ : InMux
    port map (
            O => \N__39032\,
            I => \bfn_17_18_0_\
        );

    \I__7980\ : InMux
    port map (
            O => \N__39029\,
            I => \N__39026\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__39026\,
            I => \N__39022\
        );

    \I__7978\ : InMux
    port map (
            O => \N__39025\,
            I => \N__39019\
        );

    \I__7977\ : Span4Mux_v
    port map (
            O => \N__39022\,
            I => \N__39016\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__39019\,
            I => \sCounterRAMZ0Z_1\
        );

    \I__7975\ : Odrv4
    port map (
            O => \N__39016\,
            I => \sCounterRAMZ0Z_1\
        );

    \I__7974\ : InMux
    port map (
            O => \N__39011\,
            I => \sCounterRAM_cry_0\
        );

    \I__7973\ : InMux
    port map (
            O => \N__39008\,
            I => \N__39005\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__39005\,
            I => \N__39002\
        );

    \I__7971\ : Span4Mux_v
    port map (
            O => \N__39002\,
            I => \N__38999\
        );

    \I__7970\ : Span4Mux_v
    port map (
            O => \N__38999\,
            I => \N__38996\
        );

    \I__7969\ : Odrv4
    port map (
            O => \N__38996\,
            I => \sDAC_mem_17Z0Z_4\
        );

    \I__7968\ : InMux
    port map (
            O => \N__38993\,
            I => \N__38990\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__38990\,
            I => \N__38987\
        );

    \I__7966\ : Span4Mux_v
    port map (
            O => \N__38987\,
            I => \N__38984\
        );

    \I__7965\ : Span4Mux_h
    port map (
            O => \N__38984\,
            I => \N__38981\
        );

    \I__7964\ : Odrv4
    port map (
            O => \N__38981\,
            I => \sDAC_mem_17Z0Z_5\
        );

    \I__7963\ : InMux
    port map (
            O => \N__38978\,
            I => \N__38975\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__38975\,
            I => \N__38972\
        );

    \I__7961\ : Span4Mux_h
    port map (
            O => \N__38972\,
            I => \N__38969\
        );

    \I__7960\ : Span4Mux_v
    port map (
            O => \N__38969\,
            I => \N__38966\
        );

    \I__7959\ : Odrv4
    port map (
            O => \N__38966\,
            I => \sDAC_mem_17Z0Z_6\
        );

    \I__7958\ : InMux
    port map (
            O => \N__38963\,
            I => \N__38960\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__38960\,
            I => \N__38957\
        );

    \I__7956\ : Span4Mux_h
    port map (
            O => \N__38957\,
            I => \N__38954\
        );

    \I__7955\ : Odrv4
    port map (
            O => \N__38954\,
            I => \sDAC_mem_17Z0Z_7\
        );

    \I__7954\ : InMux
    port map (
            O => \N__38951\,
            I => \N__38948\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__38948\,
            I => \N__38945\
        );

    \I__7952\ : Span4Mux_v
    port map (
            O => \N__38945\,
            I => \N__38942\
        );

    \I__7951\ : Span4Mux_h
    port map (
            O => \N__38942\,
            I => \N__38939\
        );

    \I__7950\ : Span4Mux_h
    port map (
            O => \N__38939\,
            I => \N__38936\
        );

    \I__7949\ : Span4Mux_v
    port map (
            O => \N__38936\,
            I => \N__38933\
        );

    \I__7948\ : Odrv4
    port map (
            O => \N__38933\,
            I => \RAM_DATA_in_14\
        );

    \I__7947\ : CascadeMux
    port map (
            O => \N__38930\,
            I => \N__38927\
        );

    \I__7946\ : InMux
    port map (
            O => \N__38927\,
            I => \N__38924\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__38924\,
            I => \N__38921\
        );

    \I__7944\ : Span4Mux_v
    port map (
            O => \N__38921\,
            I => \N__38918\
        );

    \I__7943\ : Sp12to4
    port map (
            O => \N__38918\,
            I => \N__38915\
        );

    \I__7942\ : Span12Mux_h
    port map (
            O => \N__38915\,
            I => \N__38912\
        );

    \I__7941\ : Span12Mux_v
    port map (
            O => \N__38912\,
            I => \N__38909\
        );

    \I__7940\ : Odrv12
    port map (
            O => \N__38909\,
            I => \RAM_DATA_in_6\
        );

    \I__7939\ : InMux
    port map (
            O => \N__38906\,
            I => \N__38902\
        );

    \I__7938\ : InMux
    port map (
            O => \N__38905\,
            I => \N__38899\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__38902\,
            I => \N__38896\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__38899\,
            I => \button_debounce_counterZ0Z_13\
        );

    \I__7935\ : Odrv4
    port map (
            O => \N__38896\,
            I => \button_debounce_counterZ0Z_13\
        );

    \I__7934\ : InMux
    port map (
            O => \N__38891\,
            I => \N__38887\
        );

    \I__7933\ : InMux
    port map (
            O => \N__38890\,
            I => \N__38884\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__38887\,
            I => \N__38881\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__38884\,
            I => \button_debounce_counterZ0Z_12\
        );

    \I__7930\ : Odrv4
    port map (
            O => \N__38881\,
            I => \button_debounce_counterZ0Z_12\
        );

    \I__7929\ : CascadeMux
    port map (
            O => \N__38876\,
            I => \N__38873\
        );

    \I__7928\ : InMux
    port map (
            O => \N__38873\,
            I => \N__38869\
        );

    \I__7927\ : InMux
    port map (
            O => \N__38872\,
            I => \N__38866\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__38869\,
            I => \N__38863\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__38866\,
            I => \button_debounce_counterZ0Z_14\
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__38863\,
            I => \button_debounce_counterZ0Z_14\
        );

    \I__7923\ : InMux
    port map (
            O => \N__38858\,
            I => \N__38854\
        );

    \I__7922\ : InMux
    port map (
            O => \N__38857\,
            I => \N__38851\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__38854\,
            I => \N__38848\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__38851\,
            I => \button_debounce_counterZ0Z_11\
        );

    \I__7919\ : Odrv4
    port map (
            O => \N__38848\,
            I => \button_debounce_counterZ0Z_11\
        );

    \I__7918\ : InMux
    port map (
            O => \N__38843\,
            I => \N__38840\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__38840\,
            I => \N__38837\
        );

    \I__7916\ : Odrv4
    port map (
            O => \N__38837\,
            I => \sbuttonModeStatus_0_sqmuxa_15\
        );

    \I__7915\ : InMux
    port map (
            O => \N__38834\,
            I => \N__38831\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__38831\,
            I => \N__38827\
        );

    \I__7913\ : InMux
    port map (
            O => \N__38830\,
            I => \N__38824\
        );

    \I__7912\ : Span4Mux_h
    port map (
            O => \N__38827\,
            I => \N__38821\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__38824\,
            I => \button_debounce_counterZ0Z_9\
        );

    \I__7910\ : Odrv4
    port map (
            O => \N__38821\,
            I => \button_debounce_counterZ0Z_9\
        );

    \I__7909\ : InMux
    port map (
            O => \N__38816\,
            I => \N__38812\
        );

    \I__7908\ : InMux
    port map (
            O => \N__38815\,
            I => \N__38809\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__38812\,
            I => \N__38806\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__38809\,
            I => \button_debounce_counterZ0Z_7\
        );

    \I__7905\ : Odrv4
    port map (
            O => \N__38806\,
            I => \button_debounce_counterZ0Z_7\
        );

    \I__7904\ : CascadeMux
    port map (
            O => \N__38801\,
            I => \N__38798\
        );

    \I__7903\ : InMux
    port map (
            O => \N__38798\,
            I => \N__38795\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__38795\,
            I => \N__38791\
        );

    \I__7901\ : InMux
    port map (
            O => \N__38794\,
            I => \N__38788\
        );

    \I__7900\ : Span4Mux_v
    port map (
            O => \N__38791\,
            I => \N__38785\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__38788\,
            I => \button_debounce_counterZ0Z_10\
        );

    \I__7898\ : Odrv4
    port map (
            O => \N__38785\,
            I => \button_debounce_counterZ0Z_10\
        );

    \I__7897\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38776\
        );

    \I__7896\ : InMux
    port map (
            O => \N__38779\,
            I => \N__38773\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__38776\,
            I => \N__38770\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__38773\,
            I => \button_debounce_counterZ0Z_8\
        );

    \I__7893\ : Odrv4
    port map (
            O => \N__38770\,
            I => \button_debounce_counterZ0Z_8\
        );

    \I__7892\ : InMux
    port map (
            O => \N__38765\,
            I => \N__38762\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__38762\,
            I => \N__38759\
        );

    \I__7890\ : Odrv12
    port map (
            O => \N__38759\,
            I => \sbuttonModeStatus_0_sqmuxa_16\
        );

    \I__7889\ : InMux
    port map (
            O => \N__38756\,
            I => \N__38753\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__38753\,
            I => \N__38750\
        );

    \I__7887\ : Span4Mux_v
    port map (
            O => \N__38750\,
            I => \N__38747\
        );

    \I__7886\ : Sp12to4
    port map (
            O => \N__38747\,
            I => \N__38744\
        );

    \I__7885\ : Span12Mux_h
    port map (
            O => \N__38744\,
            I => \N__38741\
        );

    \I__7884\ : Odrv12
    port map (
            O => \N__38741\,
            I => \RAM_DATA_in_0\
        );

    \I__7883\ : CascadeMux
    port map (
            O => \N__38738\,
            I => \N__38735\
        );

    \I__7882\ : InMux
    port map (
            O => \N__38735\,
            I => \N__38732\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__38732\,
            I => \N__38729\
        );

    \I__7880\ : Span4Mux_v
    port map (
            O => \N__38729\,
            I => \N__38726\
        );

    \I__7879\ : Span4Mux_h
    port map (
            O => \N__38726\,
            I => \N__38723\
        );

    \I__7878\ : Sp12to4
    port map (
            O => \N__38723\,
            I => \N__38720\
        );

    \I__7877\ : Span12Mux_v
    port map (
            O => \N__38720\,
            I => \N__38717\
        );

    \I__7876\ : Odrv12
    port map (
            O => \N__38717\,
            I => \RAM_DATA_in_8\
        );

    \I__7875\ : InMux
    port map (
            O => \N__38714\,
            I => \N__38711\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__38711\,
            I => \N__38708\
        );

    \I__7873\ : Span4Mux_v
    port map (
            O => \N__38708\,
            I => \N__38705\
        );

    \I__7872\ : Span4Mux_h
    port map (
            O => \N__38705\,
            I => \N__38702\
        );

    \I__7871\ : Span4Mux_h
    port map (
            O => \N__38702\,
            I => \N__38699\
        );

    \I__7870\ : IoSpan4Mux
    port map (
            O => \N__38699\,
            I => \N__38696\
        );

    \I__7869\ : Odrv4
    port map (
            O => \N__38696\,
            I => \RAM_DATA_in_12\
        );

    \I__7868\ : CascadeMux
    port map (
            O => \N__38693\,
            I => \N__38690\
        );

    \I__7867\ : InMux
    port map (
            O => \N__38690\,
            I => \N__38687\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__38687\,
            I => \N__38684\
        );

    \I__7865\ : Span4Mux_v
    port map (
            O => \N__38684\,
            I => \N__38681\
        );

    \I__7864\ : Sp12to4
    port map (
            O => \N__38681\,
            I => \N__38678\
        );

    \I__7863\ : Span12Mux_h
    port map (
            O => \N__38678\,
            I => \N__38675\
        );

    \I__7862\ : Odrv12
    port map (
            O => \N__38675\,
            I => \RAM_DATA_in_4\
        );

    \I__7861\ : InMux
    port map (
            O => \N__38672\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0\
        );

    \I__7860\ : InMux
    port map (
            O => \N__38669\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1\
        );

    \I__7859\ : InMux
    port map (
            O => \N__38666\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2\
        );

    \I__7858\ : InMux
    port map (
            O => \N__38663\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3\
        );

    \I__7857\ : InMux
    port map (
            O => \N__38660\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4\
        );

    \I__7856\ : InMux
    port map (
            O => \N__38657\,
            I => \N__38654\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__38654\,
            I => \N__38650\
        );

    \I__7854\ : InMux
    port map (
            O => \N__38653\,
            I => \N__38647\
        );

    \I__7853\ : Span4Mux_h
    port map (
            O => \N__38650\,
            I => \N__38644\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__38647\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5\
        );

    \I__7851\ : Odrv4
    port map (
            O => \N__38644\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5\
        );

    \I__7850\ : InMux
    port map (
            O => \N__38639\,
            I => \N__38636\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__38636\,
            I => \N__38633\
        );

    \I__7848\ : Odrv12
    port map (
            O => \N__38633\,
            I => \sDAC_mem_17Z0Z_0\
        );

    \I__7847\ : InMux
    port map (
            O => \N__38630\,
            I => \N__38627\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__38627\,
            I => \N__38624\
        );

    \I__7845\ : Odrv12
    port map (
            O => \N__38624\,
            I => \sDAC_mem_17Z0Z_1\
        );

    \I__7844\ : InMux
    port map (
            O => \N__38621\,
            I => \N__38618\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__38618\,
            I => \N__38615\
        );

    \I__7842\ : Odrv4
    port map (
            O => \N__38615\,
            I => \sDAC_mem_17Z0Z_2\
        );

    \I__7841\ : InMux
    port map (
            O => \N__38612\,
            I => \N__38609\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__38609\,
            I => \N__38606\
        );

    \I__7839\ : Span4Mux_h
    port map (
            O => \N__38606\,
            I => \N__38603\
        );

    \I__7838\ : Span4Mux_v
    port map (
            O => \N__38603\,
            I => \N__38600\
        );

    \I__7837\ : Odrv4
    port map (
            O => \N__38600\,
            I => \sDAC_mem_17Z0Z_3\
        );

    \I__7836\ : InMux
    port map (
            O => \N__38597\,
            I => \N__38594\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__38594\,
            I => \N__38591\
        );

    \I__7834\ : Span4Mux_h
    port map (
            O => \N__38591\,
            I => \N__38588\
        );

    \I__7833\ : Span4Mux_h
    port map (
            O => \N__38588\,
            I => \N__38585\
        );

    \I__7832\ : Span4Mux_h
    port map (
            O => \N__38585\,
            I => \N__38582\
        );

    \I__7831\ : Odrv4
    port map (
            O => \N__38582\,
            I => \sDAC_mem_29Z0Z_2\
        );

    \I__7830\ : InMux
    port map (
            O => \N__38579\,
            I => \N__38576\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__38576\,
            I => \sDAC_data_RNO_23Z0Z_5\
        );

    \I__7828\ : InMux
    port map (
            O => \N__38573\,
            I => \N__38570\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__38570\,
            I => \N__38567\
        );

    \I__7826\ : Span4Mux_v
    port map (
            O => \N__38567\,
            I => \N__38564\
        );

    \I__7825\ : Span4Mux_h
    port map (
            O => \N__38564\,
            I => \N__38561\
        );

    \I__7824\ : Odrv4
    port map (
            O => \N__38561\,
            I => \sDAC_mem_24Z0Z_3\
        );

    \I__7823\ : InMux
    port map (
            O => \N__38558\,
            I => \N__38547\
        );

    \I__7822\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38542\
        );

    \I__7821\ : InMux
    port map (
            O => \N__38556\,
            I => \N__38542\
        );

    \I__7820\ : InMux
    port map (
            O => \N__38555\,
            I => \N__38539\
        );

    \I__7819\ : InMux
    port map (
            O => \N__38554\,
            I => \N__38534\
        );

    \I__7818\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38534\
        );

    \I__7817\ : CascadeMux
    port map (
            O => \N__38552\,
            I => \N__38527\
        );

    \I__7816\ : InMux
    port map (
            O => \N__38551\,
            I => \N__38521\
        );

    \I__7815\ : InMux
    port map (
            O => \N__38550\,
            I => \N__38521\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__38547\,
            I => \N__38512\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__38542\,
            I => \N__38512\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__38539\,
            I => \N__38512\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__38534\,
            I => \N__38512\
        );

    \I__7810\ : InMux
    port map (
            O => \N__38533\,
            I => \N__38501\
        );

    \I__7809\ : InMux
    port map (
            O => \N__38532\,
            I => \N__38501\
        );

    \I__7808\ : CascadeMux
    port map (
            O => \N__38531\,
            I => \N__38497\
        );

    \I__7807\ : InMux
    port map (
            O => \N__38530\,
            I => \N__38494\
        );

    \I__7806\ : InMux
    port map (
            O => \N__38527\,
            I => \N__38491\
        );

    \I__7805\ : InMux
    port map (
            O => \N__38526\,
            I => \N__38486\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__38521\,
            I => \N__38481\
        );

    \I__7803\ : Span4Mux_v
    port map (
            O => \N__38512\,
            I => \N__38481\
        );

    \I__7802\ : InMux
    port map (
            O => \N__38511\,
            I => \N__38478\
        );

    \I__7801\ : CascadeMux
    port map (
            O => \N__38510\,
            I => \N__38473\
        );

    \I__7800\ : InMux
    port map (
            O => \N__38509\,
            I => \N__38470\
        );

    \I__7799\ : InMux
    port map (
            O => \N__38508\,
            I => \N__38467\
        );

    \I__7798\ : InMux
    port map (
            O => \N__38507\,
            I => \N__38464\
        );

    \I__7797\ : InMux
    port map (
            O => \N__38506\,
            I => \N__38461\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__38501\,
            I => \N__38456\
        );

    \I__7795\ : InMux
    port map (
            O => \N__38500\,
            I => \N__38453\
        );

    \I__7794\ : InMux
    port map (
            O => \N__38497\,
            I => \N__38449\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__38494\,
            I => \N__38445\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__38491\,
            I => \N__38442\
        );

    \I__7791\ : InMux
    port map (
            O => \N__38490\,
            I => \N__38437\
        );

    \I__7790\ : InMux
    port map (
            O => \N__38489\,
            I => \N__38437\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__38486\,
            I => \N__38430\
        );

    \I__7788\ : Span4Mux_v
    port map (
            O => \N__38481\,
            I => \N__38430\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__38478\,
            I => \N__38430\
        );

    \I__7786\ : InMux
    port map (
            O => \N__38477\,
            I => \N__38427\
        );

    \I__7785\ : InMux
    port map (
            O => \N__38476\,
            I => \N__38420\
        );

    \I__7784\ : InMux
    port map (
            O => \N__38473\,
            I => \N__38420\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__38470\,
            I => \N__38415\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__38467\,
            I => \N__38415\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__38464\,
            I => \N__38409\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__38461\,
            I => \N__38409\
        );

    \I__7779\ : InMux
    port map (
            O => \N__38460\,
            I => \N__38404\
        );

    \I__7778\ : InMux
    port map (
            O => \N__38459\,
            I => \N__38404\
        );

    \I__7777\ : Span4Mux_v
    port map (
            O => \N__38456\,
            I => \N__38397\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__38453\,
            I => \N__38397\
        );

    \I__7775\ : InMux
    port map (
            O => \N__38452\,
            I => \N__38394\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__38449\,
            I => \N__38391\
        );

    \I__7773\ : InMux
    port map (
            O => \N__38448\,
            I => \N__38388\
        );

    \I__7772\ : Span4Mux_v
    port map (
            O => \N__38445\,
            I => \N__38384\
        );

    \I__7771\ : Span4Mux_h
    port map (
            O => \N__38442\,
            I => \N__38375\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__38437\,
            I => \N__38375\
        );

    \I__7769\ : Span4Mux_h
    port map (
            O => \N__38430\,
            I => \N__38375\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__38427\,
            I => \N__38375\
        );

    \I__7767\ : InMux
    port map (
            O => \N__38426\,
            I => \N__38372\
        );

    \I__7766\ : InMux
    port map (
            O => \N__38425\,
            I => \N__38369\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__38420\,
            I => \N__38364\
        );

    \I__7764\ : Span4Mux_h
    port map (
            O => \N__38415\,
            I => \N__38364\
        );

    \I__7763\ : InMux
    port map (
            O => \N__38414\,
            I => \N__38361\
        );

    \I__7762\ : Span4Mux_v
    port map (
            O => \N__38409\,
            I => \N__38356\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__38404\,
            I => \N__38356\
        );

    \I__7760\ : InMux
    port map (
            O => \N__38403\,
            I => \N__38353\
        );

    \I__7759\ : InMux
    port map (
            O => \N__38402\,
            I => \N__38350\
        );

    \I__7758\ : Span4Mux_v
    port map (
            O => \N__38397\,
            I => \N__38347\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__38394\,
            I => \N__38340\
        );

    \I__7756\ : Span4Mux_v
    port map (
            O => \N__38391\,
            I => \N__38340\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__38388\,
            I => \N__38340\
        );

    \I__7754\ : InMux
    port map (
            O => \N__38387\,
            I => \N__38337\
        );

    \I__7753\ : Span4Mux_h
    port map (
            O => \N__38384\,
            I => \N__38332\
        );

    \I__7752\ : Span4Mux_v
    port map (
            O => \N__38375\,
            I => \N__38332\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__38372\,
            I => \N__38321\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__38369\,
            I => \N__38321\
        );

    \I__7749\ : Span4Mux_v
    port map (
            O => \N__38364\,
            I => \N__38321\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__38361\,
            I => \N__38321\
        );

    \I__7747\ : Span4Mux_h
    port map (
            O => \N__38356\,
            I => \N__38321\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__38353\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__38350\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__7744\ : Odrv4
    port map (
            O => \N__38347\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__7743\ : Odrv4
    port map (
            O => \N__38340\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__38337\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__7741\ : Odrv4
    port map (
            O => \N__38332\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__7740\ : Odrv4
    port map (
            O => \N__38321\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__7739\ : CascadeMux
    port map (
            O => \N__38306\,
            I => \sDAC_data_RNO_30Z0Z_6_cascade_\
        );

    \I__7738\ : InMux
    port map (
            O => \N__38303\,
            I => \N__38297\
        );

    \I__7737\ : InMux
    port map (
            O => \N__38302\,
            I => \N__38292\
        );

    \I__7736\ : InMux
    port map (
            O => \N__38301\,
            I => \N__38292\
        );

    \I__7735\ : InMux
    port map (
            O => \N__38300\,
            I => \N__38282\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__38297\,
            I => \N__38277\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__38292\,
            I => \N__38277\
        );

    \I__7732\ : InMux
    port map (
            O => \N__38291\,
            I => \N__38272\
        );

    \I__7731\ : InMux
    port map (
            O => \N__38290\,
            I => \N__38272\
        );

    \I__7730\ : InMux
    port map (
            O => \N__38289\,
            I => \N__38263\
        );

    \I__7729\ : InMux
    port map (
            O => \N__38288\,
            I => \N__38263\
        );

    \I__7728\ : InMux
    port map (
            O => \N__38287\,
            I => \N__38263\
        );

    \I__7727\ : InMux
    port map (
            O => \N__38286\,
            I => \N__38263\
        );

    \I__7726\ : CascadeMux
    port map (
            O => \N__38285\,
            I => \N__38259\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__38282\,
            I => \N__38246\
        );

    \I__7724\ : Span4Mux_v
    port map (
            O => \N__38277\,
            I => \N__38239\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__38272\,
            I => \N__38239\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__38263\,
            I => \N__38239\
        );

    \I__7721\ : InMux
    port map (
            O => \N__38262\,
            I => \N__38234\
        );

    \I__7720\ : InMux
    port map (
            O => \N__38259\,
            I => \N__38234\
        );

    \I__7719\ : CascadeMux
    port map (
            O => \N__38258\,
            I => \N__38227\
        );

    \I__7718\ : CascadeMux
    port map (
            O => \N__38257\,
            I => \N__38224\
        );

    \I__7717\ : CascadeMux
    port map (
            O => \N__38256\,
            I => \N__38221\
        );

    \I__7716\ : CascadeMux
    port map (
            O => \N__38255\,
            I => \N__38218\
        );

    \I__7715\ : CascadeMux
    port map (
            O => \N__38254\,
            I => \N__38213\
        );

    \I__7714\ : CascadeMux
    port map (
            O => \N__38253\,
            I => \N__38204\
        );

    \I__7713\ : InMux
    port map (
            O => \N__38252\,
            I => \N__38197\
        );

    \I__7712\ : CascadeMux
    port map (
            O => \N__38251\,
            I => \N__38191\
        );

    \I__7711\ : InMux
    port map (
            O => \N__38250\,
            I => \N__38185\
        );

    \I__7710\ : InMux
    port map (
            O => \N__38249\,
            I => \N__38185\
        );

    \I__7709\ : Span4Mux_h
    port map (
            O => \N__38246\,
            I => \N__38178\
        );

    \I__7708\ : Span4Mux_v
    port map (
            O => \N__38239\,
            I => \N__38178\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__38234\,
            I => \N__38178\
        );

    \I__7706\ : CascadeMux
    port map (
            O => \N__38233\,
            I => \N__38174\
        );

    \I__7705\ : CascadeMux
    port map (
            O => \N__38232\,
            I => \N__38171\
        );

    \I__7704\ : InMux
    port map (
            O => \N__38231\,
            I => \N__38163\
        );

    \I__7703\ : InMux
    port map (
            O => \N__38230\,
            I => \N__38156\
        );

    \I__7702\ : InMux
    port map (
            O => \N__38227\,
            I => \N__38156\
        );

    \I__7701\ : InMux
    port map (
            O => \N__38224\,
            I => \N__38156\
        );

    \I__7700\ : InMux
    port map (
            O => \N__38221\,
            I => \N__38151\
        );

    \I__7699\ : InMux
    port map (
            O => \N__38218\,
            I => \N__38151\
        );

    \I__7698\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38144\
        );

    \I__7697\ : InMux
    port map (
            O => \N__38216\,
            I => \N__38144\
        );

    \I__7696\ : InMux
    port map (
            O => \N__38213\,
            I => \N__38144\
        );

    \I__7695\ : CascadeMux
    port map (
            O => \N__38212\,
            I => \N__38141\
        );

    \I__7694\ : CascadeMux
    port map (
            O => \N__38211\,
            I => \N__38138\
        );

    \I__7693\ : CascadeMux
    port map (
            O => \N__38210\,
            I => \N__38135\
        );

    \I__7692\ : CascadeMux
    port map (
            O => \N__38209\,
            I => \N__38132\
        );

    \I__7691\ : CascadeMux
    port map (
            O => \N__38208\,
            I => \N__38126\
        );

    \I__7690\ : CascadeMux
    port map (
            O => \N__38207\,
            I => \N__38123\
        );

    \I__7689\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38118\
        );

    \I__7688\ : CascadeMux
    port map (
            O => \N__38203\,
            I => \N__38112\
        );

    \I__7687\ : InMux
    port map (
            O => \N__38202\,
            I => \N__38108\
        );

    \I__7686\ : CascadeMux
    port map (
            O => \N__38201\,
            I => \N__38105\
        );

    \I__7685\ : CascadeMux
    port map (
            O => \N__38200\,
            I => \N__38101\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__38197\,
            I => \N__38098\
        );

    \I__7683\ : CascadeMux
    port map (
            O => \N__38196\,
            I => \N__38092\
        );

    \I__7682\ : CascadeMux
    port map (
            O => \N__38195\,
            I => \N__38088\
        );

    \I__7681\ : InMux
    port map (
            O => \N__38194\,
            I => \N__38083\
        );

    \I__7680\ : InMux
    port map (
            O => \N__38191\,
            I => \N__38083\
        );

    \I__7679\ : InMux
    port map (
            O => \N__38190\,
            I => \N__38080\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__38185\,
            I => \N__38075\
        );

    \I__7677\ : Span4Mux_v
    port map (
            O => \N__38178\,
            I => \N__38075\
        );

    \I__7676\ : InMux
    port map (
            O => \N__38177\,
            I => \N__38066\
        );

    \I__7675\ : InMux
    port map (
            O => \N__38174\,
            I => \N__38066\
        );

    \I__7674\ : InMux
    port map (
            O => \N__38171\,
            I => \N__38066\
        );

    \I__7673\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38066\
        );

    \I__7672\ : InMux
    port map (
            O => \N__38169\,
            I => \N__38061\
        );

    \I__7671\ : InMux
    port map (
            O => \N__38168\,
            I => \N__38061\
        );

    \I__7670\ : InMux
    port map (
            O => \N__38167\,
            I => \N__38056\
        );

    \I__7669\ : InMux
    port map (
            O => \N__38166\,
            I => \N__38056\
        );

    \I__7668\ : LocalMux
    port map (
            O => \N__38163\,
            I => \N__38053\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__38156\,
            I => \N__38048\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__38151\,
            I => \N__38048\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__38144\,
            I => \N__38045\
        );

    \I__7664\ : InMux
    port map (
            O => \N__38141\,
            I => \N__38042\
        );

    \I__7663\ : InMux
    port map (
            O => \N__38138\,
            I => \N__38035\
        );

    \I__7662\ : InMux
    port map (
            O => \N__38135\,
            I => \N__38035\
        );

    \I__7661\ : InMux
    port map (
            O => \N__38132\,
            I => \N__38035\
        );

    \I__7660\ : InMux
    port map (
            O => \N__38131\,
            I => \N__38032\
        );

    \I__7659\ : InMux
    port map (
            O => \N__38130\,
            I => \N__38025\
        );

    \I__7658\ : InMux
    port map (
            O => \N__38129\,
            I => \N__38025\
        );

    \I__7657\ : InMux
    port map (
            O => \N__38126\,
            I => \N__38020\
        );

    \I__7656\ : InMux
    port map (
            O => \N__38123\,
            I => \N__38020\
        );

    \I__7655\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38015\
        );

    \I__7654\ : InMux
    port map (
            O => \N__38121\,
            I => \N__38015\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__38118\,
            I => \N__38012\
        );

    \I__7652\ : InMux
    port map (
            O => \N__38117\,
            I => \N__38009\
        );

    \I__7651\ : InMux
    port map (
            O => \N__38116\,
            I => \N__38002\
        );

    \I__7650\ : InMux
    port map (
            O => \N__38115\,
            I => \N__38002\
        );

    \I__7649\ : InMux
    port map (
            O => \N__38112\,
            I => \N__38002\
        );

    \I__7648\ : InMux
    port map (
            O => \N__38111\,
            I => \N__37998\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__38108\,
            I => \N__37994\
        );

    \I__7646\ : InMux
    port map (
            O => \N__38105\,
            I => \N__37989\
        );

    \I__7645\ : InMux
    port map (
            O => \N__38104\,
            I => \N__37989\
        );

    \I__7644\ : InMux
    port map (
            O => \N__38101\,
            I => \N__37986\
        );

    \I__7643\ : Span4Mux_v
    port map (
            O => \N__38098\,
            I => \N__37983\
        );

    \I__7642\ : InMux
    port map (
            O => \N__38097\,
            I => \N__37980\
        );

    \I__7641\ : InMux
    port map (
            O => \N__38096\,
            I => \N__37975\
        );

    \I__7640\ : InMux
    port map (
            O => \N__38095\,
            I => \N__37975\
        );

    \I__7639\ : InMux
    port map (
            O => \N__38092\,
            I => \N__37968\
        );

    \I__7638\ : InMux
    port map (
            O => \N__38091\,
            I => \N__37968\
        );

    \I__7637\ : InMux
    port map (
            O => \N__38088\,
            I => \N__37968\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__38083\,
            I => \N__37959\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__38080\,
            I => \N__37959\
        );

    \I__7634\ : Span4Mux_h
    port map (
            O => \N__38075\,
            I => \N__37959\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__38066\,
            I => \N__37959\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__38061\,
            I => \N__37948\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__38056\,
            I => \N__37948\
        );

    \I__7630\ : Span4Mux_h
    port map (
            O => \N__38053\,
            I => \N__37948\
        );

    \I__7629\ : Span4Mux_v
    port map (
            O => \N__38048\,
            I => \N__37948\
        );

    \I__7628\ : Span4Mux_h
    port map (
            O => \N__38045\,
            I => \N__37948\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__38042\,
            I => \N__37943\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__38035\,
            I => \N__37943\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__38032\,
            I => \N__37940\
        );

    \I__7624\ : InMux
    port map (
            O => \N__38031\,
            I => \N__37937\
        );

    \I__7623\ : InMux
    port map (
            O => \N__38030\,
            I => \N__37934\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__38025\,
            I => \N__37929\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__38020\,
            I => \N__37929\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__38015\,
            I => \N__37926\
        );

    \I__7619\ : Span4Mux_h
    port map (
            O => \N__38012\,
            I => \N__37919\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__38009\,
            I => \N__37919\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__38002\,
            I => \N__37919\
        );

    \I__7616\ : InMux
    port map (
            O => \N__38001\,
            I => \N__37916\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__37998\,
            I => \N__37913\
        );

    \I__7614\ : InMux
    port map (
            O => \N__37997\,
            I => \N__37910\
        );

    \I__7613\ : Span4Mux_v
    port map (
            O => \N__37994\,
            I => \N__37907\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__37989\,
            I => \N__37902\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__37986\,
            I => \N__37902\
        );

    \I__7610\ : Span4Mux_h
    port map (
            O => \N__37983\,
            I => \N__37891\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__37980\,
            I => \N__37891\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__37975\,
            I => \N__37891\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__37968\,
            I => \N__37891\
        );

    \I__7606\ : Span4Mux_v
    port map (
            O => \N__37959\,
            I => \N__37891\
        );

    \I__7605\ : Span4Mux_v
    port map (
            O => \N__37948\,
            I => \N__37886\
        );

    \I__7604\ : Span4Mux_h
    port map (
            O => \N__37943\,
            I => \N__37886\
        );

    \I__7603\ : Span12Mux_h
    port map (
            O => \N__37940\,
            I => \N__37873\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__37937\,
            I => \N__37873\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__37934\,
            I => \N__37873\
        );

    \I__7600\ : Span12Mux_h
    port map (
            O => \N__37929\,
            I => \N__37873\
        );

    \I__7599\ : Sp12to4
    port map (
            O => \N__37926\,
            I => \N__37873\
        );

    \I__7598\ : Sp12to4
    port map (
            O => \N__37919\,
            I => \N__37873\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__37916\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__7596\ : Odrv12
    port map (
            O => \N__37913\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__37910\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__7594\ : Odrv4
    port map (
            O => \N__37907\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__7593\ : Odrv4
    port map (
            O => \N__37902\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__7592\ : Odrv4
    port map (
            O => \N__37891\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__7591\ : Odrv4
    port map (
            O => \N__37886\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__7590\ : Odrv12
    port map (
            O => \N__37873\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__7589\ : InMux
    port map (
            O => \N__37856\,
            I => \N__37853\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__37853\,
            I => \N__37850\
        );

    \I__7587\ : Span4Mux_v
    port map (
            O => \N__37850\,
            I => \N__37847\
        );

    \I__7586\ : Odrv4
    port map (
            O => \N__37847\,
            I => \sDAC_data_RNO_24Z0Z_6\
        );

    \I__7585\ : CascadeMux
    port map (
            O => \N__37844\,
            I => \sDAC_data_2_39_ns_1_6_cascade_\
        );

    \I__7584\ : InMux
    port map (
            O => \N__37841\,
            I => \N__37838\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__37838\,
            I => \N__37835\
        );

    \I__7582\ : Span4Mux_h
    port map (
            O => \N__37835\,
            I => \N__37832\
        );

    \I__7581\ : Odrv4
    port map (
            O => \N__37832\,
            I => \sDAC_data_RNO_23Z0Z_6\
        );

    \I__7580\ : InMux
    port map (
            O => \N__37829\,
            I => \N__37826\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__37826\,
            I => \N__37823\
        );

    \I__7578\ : Span4Mux_v
    port map (
            O => \N__37823\,
            I => \N__37820\
        );

    \I__7577\ : Span4Mux_h
    port map (
            O => \N__37820\,
            I => \N__37817\
        );

    \I__7576\ : Odrv4
    port map (
            O => \N__37817\,
            I => \sDAC_data_RNO_11Z0Z_6\
        );

    \I__7575\ : InMux
    port map (
            O => \N__37814\,
            I => \N__37811\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__37811\,
            I => \sDAC_mem_28Z0Z_2\
        );

    \I__7573\ : CEMux
    port map (
            O => \N__37808\,
            I => \N__37803\
        );

    \I__7572\ : CEMux
    port map (
            O => \N__37807\,
            I => \N__37800\
        );

    \I__7571\ : CEMux
    port map (
            O => \N__37806\,
            I => \N__37797\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__37803\,
            I => \N__37793\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__37800\,
            I => \N__37790\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__37797\,
            I => \N__37786\
        );

    \I__7567\ : CEMux
    port map (
            O => \N__37796\,
            I => \N__37783\
        );

    \I__7566\ : Span4Mux_h
    port map (
            O => \N__37793\,
            I => \N__37780\
        );

    \I__7565\ : Span4Mux_v
    port map (
            O => \N__37790\,
            I => \N__37777\
        );

    \I__7564\ : CEMux
    port map (
            O => \N__37789\,
            I => \N__37774\
        );

    \I__7563\ : Span4Mux_v
    port map (
            O => \N__37786\,
            I => \N__37771\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__37783\,
            I => \N__37768\
        );

    \I__7561\ : Span4Mux_h
    port map (
            O => \N__37780\,
            I => \N__37765\
        );

    \I__7560\ : Span4Mux_h
    port map (
            O => \N__37777\,
            I => \N__37760\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__37774\,
            I => \N__37760\
        );

    \I__7558\ : Span4Mux_h
    port map (
            O => \N__37771\,
            I => \N__37755\
        );

    \I__7557\ : Span4Mux_v
    port map (
            O => \N__37768\,
            I => \N__37755\
        );

    \I__7556\ : Span4Mux_v
    port map (
            O => \N__37765\,
            I => \N__37752\
        );

    \I__7555\ : Span4Mux_v
    port map (
            O => \N__37760\,
            I => \N__37749\
        );

    \I__7554\ : Span4Mux_h
    port map (
            O => \N__37755\,
            I => \N__37746\
        );

    \I__7553\ : Odrv4
    port map (
            O => \N__37752\,
            I => \sDAC_mem_28_1_sqmuxa\
        );

    \I__7552\ : Odrv4
    port map (
            O => \N__37749\,
            I => \sDAC_mem_28_1_sqmuxa\
        );

    \I__7551\ : Odrv4
    port map (
            O => \N__37746\,
            I => \sDAC_mem_28_1_sqmuxa\
        );

    \I__7550\ : InMux
    port map (
            O => \N__37739\,
            I => \N__37736\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__37736\,
            I => \N__37733\
        );

    \I__7548\ : Span4Mux_h
    port map (
            O => \N__37733\,
            I => \N__37730\
        );

    \I__7547\ : Span4Mux_h
    port map (
            O => \N__37730\,
            I => \N__37727\
        );

    \I__7546\ : Odrv4
    port map (
            O => \N__37727\,
            I => \sDAC_mem_30Z0Z_2\
        );

    \I__7545\ : InMux
    port map (
            O => \N__37724\,
            I => \N__37721\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__37721\,
            I => \N__37718\
        );

    \I__7543\ : Span12Mux_h
    port map (
            O => \N__37718\,
            I => \N__37715\
        );

    \I__7542\ : Odrv12
    port map (
            O => \N__37715\,
            I => \sDAC_mem_31Z0Z_2\
        );

    \I__7541\ : InMux
    port map (
            O => \N__37712\,
            I => \N__37709\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__37709\,
            I => \sDAC_data_RNO_24Z0Z_5\
        );

    \I__7539\ : InMux
    port map (
            O => \N__37706\,
            I => \N__37703\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__37703\,
            I => \N__37700\
        );

    \I__7537\ : Span12Mux_h
    port map (
            O => \N__37700\,
            I => \N__37697\
        );

    \I__7536\ : Odrv12
    port map (
            O => \N__37697\,
            I => \sDAC_mem_26Z0Z_3\
        );

    \I__7535\ : InMux
    port map (
            O => \N__37694\,
            I => \N__37691\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__37691\,
            I => \N__37688\
        );

    \I__7533\ : Span4Mux_h
    port map (
            O => \N__37688\,
            I => \N__37685\
        );

    \I__7532\ : Odrv4
    port map (
            O => \N__37685\,
            I => \sDAC_mem_27Z0Z_3\
        );

    \I__7531\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37679\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__37679\,
            I => \sDAC_data_RNO_31Z0Z_6\
        );

    \I__7529\ : InMux
    port map (
            O => \N__37676\,
            I => \N__37673\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__37673\,
            I => \N__37670\
        );

    \I__7527\ : Span4Mux_h
    port map (
            O => \N__37670\,
            I => \N__37667\
        );

    \I__7526\ : Odrv4
    port map (
            O => \N__37667\,
            I => \sDAC_data_RNO_5Z0Z_3\
        );

    \I__7525\ : InMux
    port map (
            O => \N__37664\,
            I => \N__37661\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__37661\,
            I => \sDAC_data_RNO_2Z0Z_3\
        );

    \I__7523\ : CascadeMux
    port map (
            O => \N__37658\,
            I => \sDAC_data_RNO_1Z0Z_3_cascade_\
        );

    \I__7522\ : InMux
    port map (
            O => \N__37655\,
            I => \N__37652\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__37652\,
            I => \N__37649\
        );

    \I__7520\ : Span4Mux_v
    port map (
            O => \N__37649\,
            I => \N__37646\
        );

    \I__7519\ : Span4Mux_v
    port map (
            O => \N__37646\,
            I => \N__37643\
        );

    \I__7518\ : Odrv4
    port map (
            O => \N__37643\,
            I => \sEEDACZ0Z_0\
        );

    \I__7517\ : CascadeMux
    port map (
            O => \N__37640\,
            I => \sDAC_data_2_3_cascade_\
        );

    \I__7516\ : InMux
    port map (
            O => \N__37637\,
            I => \N__37624\
        );

    \I__7515\ : InMux
    port map (
            O => \N__37636\,
            I => \N__37621\
        );

    \I__7514\ : InMux
    port map (
            O => \N__37635\,
            I => \N__37618\
        );

    \I__7513\ : InMux
    port map (
            O => \N__37634\,
            I => \N__37611\
        );

    \I__7512\ : InMux
    port map (
            O => \N__37633\,
            I => \N__37611\
        );

    \I__7511\ : InMux
    port map (
            O => \N__37632\,
            I => \N__37611\
        );

    \I__7510\ : InMux
    port map (
            O => \N__37631\,
            I => \N__37608\
        );

    \I__7509\ : InMux
    port map (
            O => \N__37630\,
            I => \N__37605\
        );

    \I__7508\ : InMux
    port map (
            O => \N__37629\,
            I => \N__37602\
        );

    \I__7507\ : InMux
    port map (
            O => \N__37628\,
            I => \N__37599\
        );

    \I__7506\ : InMux
    port map (
            O => \N__37627\,
            I => \N__37596\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__37624\,
            I => \N__37593\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__37621\,
            I => \N__37590\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__37618\,
            I => \N__37585\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__37611\,
            I => \N__37585\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__37608\,
            I => \N__37579\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__37605\,
            I => \N__37576\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__37602\,
            I => \N__37573\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__37599\,
            I => \N__37564\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__37596\,
            I => \N__37564\
        );

    \I__7496\ : Span4Mux_h
    port map (
            O => \N__37593\,
            I => \N__37564\
        );

    \I__7495\ : Span4Mux_h
    port map (
            O => \N__37590\,
            I => \N__37564\
        );

    \I__7494\ : Span4Mux_v
    port map (
            O => \N__37585\,
            I => \N__37561\
        );

    \I__7493\ : InMux
    port map (
            O => \N__37584\,
            I => \N__37554\
        );

    \I__7492\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37554\
        );

    \I__7491\ : InMux
    port map (
            O => \N__37582\,
            I => \N__37554\
        );

    \I__7490\ : Span4Mux_h
    port map (
            O => \N__37579\,
            I => \N__37551\
        );

    \I__7489\ : Span4Mux_v
    port map (
            O => \N__37576\,
            I => \N__37548\
        );

    \I__7488\ : Span4Mux_v
    port map (
            O => \N__37573\,
            I => \N__37545\
        );

    \I__7487\ : Span4Mux_v
    port map (
            O => \N__37564\,
            I => \N__37542\
        );

    \I__7486\ : Span4Mux_v
    port map (
            O => \N__37561\,
            I => \N__37539\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__37554\,
            I => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\
        );

    \I__7484\ : Odrv4
    port map (
            O => \N__37551\,
            I => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\
        );

    \I__7483\ : Odrv4
    port map (
            O => \N__37548\,
            I => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\
        );

    \I__7482\ : Odrv4
    port map (
            O => \N__37545\,
            I => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\
        );

    \I__7481\ : Odrv4
    port map (
            O => \N__37542\,
            I => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\
        );

    \I__7480\ : Odrv4
    port map (
            O => \N__37539\,
            I => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\
        );

    \I__7479\ : InMux
    port map (
            O => \N__37526\,
            I => \N__37523\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__37523\,
            I => \N__37520\
        );

    \I__7477\ : Span4Mux_h
    port map (
            O => \N__37520\,
            I => \N__37517\
        );

    \I__7476\ : Span4Mux_v
    port map (
            O => \N__37517\,
            I => \N__37514\
        );

    \I__7475\ : Odrv4
    port map (
            O => \N__37514\,
            I => \sDAC_dataZ0Z_3\
        );

    \I__7474\ : InMux
    port map (
            O => \N__37511\,
            I => \N__37508\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__37508\,
            I => \N__37505\
        );

    \I__7472\ : Span4Mux_v
    port map (
            O => \N__37505\,
            I => \N__37502\
        );

    \I__7471\ : Odrv4
    port map (
            O => \N__37502\,
            I => \sDAC_data_RNO_21Z0Z_3\
        );

    \I__7470\ : InMux
    port map (
            O => \N__37499\,
            I => \N__37496\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__37496\,
            I => \N__37493\
        );

    \I__7468\ : Span4Mux_v
    port map (
            O => \N__37493\,
            I => \N__37490\
        );

    \I__7467\ : Odrv4
    port map (
            O => \N__37490\,
            I => \sDAC_data_RNO_20Z0Z_3\
        );

    \I__7466\ : CascadeMux
    port map (
            O => \N__37487\,
            I => \N__37482\
        );

    \I__7465\ : InMux
    port map (
            O => \N__37486\,
            I => \N__37478\
        );

    \I__7464\ : InMux
    port map (
            O => \N__37485\,
            I => \N__37473\
        );

    \I__7463\ : InMux
    port map (
            O => \N__37482\,
            I => \N__37473\
        );

    \I__7462\ : CascadeMux
    port map (
            O => \N__37481\,
            I => \N__37468\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__37478\,
            I => \N__37463\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__37473\,
            I => \N__37463\
        );

    \I__7459\ : CascadeMux
    port map (
            O => \N__37472\,
            I => \N__37458\
        );

    \I__7458\ : InMux
    port map (
            O => \N__37471\,
            I => \N__37449\
        );

    \I__7457\ : InMux
    port map (
            O => \N__37468\,
            I => \N__37449\
        );

    \I__7456\ : Span4Mux_v
    port map (
            O => \N__37463\,
            I => \N__37446\
        );

    \I__7455\ : InMux
    port map (
            O => \N__37462\,
            I => \N__37443\
        );

    \I__7454\ : InMux
    port map (
            O => \N__37461\,
            I => \N__37436\
        );

    \I__7453\ : InMux
    port map (
            O => \N__37458\,
            I => \N__37433\
        );

    \I__7452\ : InMux
    port map (
            O => \N__37457\,
            I => \N__37428\
        );

    \I__7451\ : InMux
    port map (
            O => \N__37456\,
            I => \N__37428\
        );

    \I__7450\ : InMux
    port map (
            O => \N__37455\,
            I => \N__37423\
        );

    \I__7449\ : InMux
    port map (
            O => \N__37454\,
            I => \N__37423\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__37449\,
            I => \N__37420\
        );

    \I__7447\ : Span4Mux_h
    port map (
            O => \N__37446\,
            I => \N__37416\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__37443\,
            I => \N__37413\
        );

    \I__7445\ : InMux
    port map (
            O => \N__37442\,
            I => \N__37408\
        );

    \I__7444\ : InMux
    port map (
            O => \N__37441\,
            I => \N__37408\
        );

    \I__7443\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37403\
        );

    \I__7442\ : InMux
    port map (
            O => \N__37439\,
            I => \N__37403\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__37436\,
            I => \N__37396\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__37433\,
            I => \N__37396\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__37428\,
            I => \N__37396\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__37423\,
            I => \N__37391\
        );

    \I__7437\ : Span4Mux_h
    port map (
            O => \N__37420\,
            I => \N__37391\
        );

    \I__7436\ : InMux
    port map (
            O => \N__37419\,
            I => \N__37387\
        );

    \I__7435\ : Sp12to4
    port map (
            O => \N__37416\,
            I => \N__37382\
        );

    \I__7434\ : Sp12to4
    port map (
            O => \N__37413\,
            I => \N__37382\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__37408\,
            I => \N__37379\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__37403\,
            I => \N__37376\
        );

    \I__7431\ : Span4Mux_v
    port map (
            O => \N__37396\,
            I => \N__37371\
        );

    \I__7430\ : Span4Mux_v
    port map (
            O => \N__37391\,
            I => \N__37371\
        );

    \I__7429\ : InMux
    port map (
            O => \N__37390\,
            I => \N__37368\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__37387\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__7427\ : Odrv12
    port map (
            O => \N__37382\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__7426\ : Odrv4
    port map (
            O => \N__37379\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__7425\ : Odrv12
    port map (
            O => \N__37376\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__7424\ : Odrv4
    port map (
            O => \N__37371\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__37368\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__7422\ : InMux
    port map (
            O => \N__37355\,
            I => \N__37352\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__37352\,
            I => \N__37348\
        );

    \I__7420\ : InMux
    port map (
            O => \N__37351\,
            I => \N__37345\
        );

    \I__7419\ : Span4Mux_v
    port map (
            O => \N__37348\,
            I => \N__37336\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__37345\,
            I => \N__37336\
        );

    \I__7417\ : InMux
    port map (
            O => \N__37344\,
            I => \N__37331\
        );

    \I__7416\ : InMux
    port map (
            O => \N__37343\,
            I => \N__37328\
        );

    \I__7415\ : InMux
    port map (
            O => \N__37342\,
            I => \N__37324\
        );

    \I__7414\ : InMux
    port map (
            O => \N__37341\,
            I => \N__37321\
        );

    \I__7413\ : Span4Mux_h
    port map (
            O => \N__37336\,
            I => \N__37318\
        );

    \I__7412\ : InMux
    port map (
            O => \N__37335\,
            I => \N__37315\
        );

    \I__7411\ : InMux
    port map (
            O => \N__37334\,
            I => \N__37312\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__37331\,
            I => \N__37309\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__37328\,
            I => \N__37306\
        );

    \I__7408\ : InMux
    port map (
            O => \N__37327\,
            I => \N__37302\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__37324\,
            I => \N__37297\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__37321\,
            I => \N__37297\
        );

    \I__7405\ : Span4Mux_h
    port map (
            O => \N__37318\,
            I => \N__37290\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__37315\,
            I => \N__37290\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__37312\,
            I => \N__37290\
        );

    \I__7402\ : Span4Mux_h
    port map (
            O => \N__37309\,
            I => \N__37285\
        );

    \I__7401\ : Span4Mux_v
    port map (
            O => \N__37306\,
            I => \N__37285\
        );

    \I__7400\ : InMux
    port map (
            O => \N__37305\,
            I => \N__37282\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__37302\,
            I => \sDAC_mem_pointerZ0Z_3\
        );

    \I__7398\ : Odrv4
    port map (
            O => \N__37297\,
            I => \sDAC_mem_pointerZ0Z_3\
        );

    \I__7397\ : Odrv4
    port map (
            O => \N__37290\,
            I => \sDAC_mem_pointerZ0Z_3\
        );

    \I__7396\ : Odrv4
    port map (
            O => \N__37285\,
            I => \sDAC_mem_pointerZ0Z_3\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__37282\,
            I => \sDAC_mem_pointerZ0Z_3\
        );

    \I__7394\ : CascadeMux
    port map (
            O => \N__37271\,
            I => \sDAC_data_RNO_10Z0Z_3_cascade_\
        );

    \I__7393\ : InMux
    port map (
            O => \N__37268\,
            I => \N__37265\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__37265\,
            I => \N__37262\
        );

    \I__7391\ : Span4Mux_h
    port map (
            O => \N__37262\,
            I => \N__37259\
        );

    \I__7390\ : Odrv4
    port map (
            O => \N__37259\,
            I => \sDAC_data_RNO_11Z0Z_3\
        );

    \I__7389\ : InMux
    port map (
            O => \N__37256\,
            I => \N__37253\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__37253\,
            I => \sDAC_data_2_41_ns_1_3\
        );

    \I__7387\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37247\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__37247\,
            I => \sDAC_data_RNO_15Z0Z_3\
        );

    \I__7385\ : InMux
    port map (
            O => \N__37244\,
            I => \N__37241\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__37241\,
            I => \sDAC_data_2_14_ns_1_3\
        );

    \I__7383\ : InMux
    port map (
            O => \N__37238\,
            I => \N__37235\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__37235\,
            I => \N__37232\
        );

    \I__7381\ : Span4Mux_v
    port map (
            O => \N__37232\,
            I => \N__37229\
        );

    \I__7380\ : Odrv4
    port map (
            O => \N__37229\,
            I => \sDAC_data_RNO_28Z0Z_3\
        );

    \I__7379\ : InMux
    port map (
            O => \N__37226\,
            I => \N__37223\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__37223\,
            I => \sDAC_data_RNO_29Z0Z_3\
        );

    \I__7377\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37217\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__37217\,
            I => \sDAC_data_2_32_ns_1_3\
        );

    \I__7375\ : InMux
    port map (
            O => \N__37214\,
            I => \N__37211\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__37211\,
            I => \N__37208\
        );

    \I__7373\ : Odrv12
    port map (
            O => \N__37208\,
            I => \sDAC_data_2_39_ns_1_5\
        );

    \I__7372\ : InMux
    port map (
            O => \N__37205\,
            I => \N__37202\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__37202\,
            I => \N__37199\
        );

    \I__7370\ : Odrv4
    port map (
            O => \N__37199\,
            I => \sDAC_data_RNO_11Z0Z_5\
        );

    \I__7369\ : InMux
    port map (
            O => \N__37196\,
            I => \N__37193\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__37193\,
            I => \N__37190\
        );

    \I__7367\ : Span4Mux_v
    port map (
            O => \N__37190\,
            I => \N__37187\
        );

    \I__7366\ : Span4Mux_v
    port map (
            O => \N__37187\,
            I => \N__37184\
        );

    \I__7365\ : Odrv4
    port map (
            O => \N__37184\,
            I => \sDAC_mem_pointerZ0Z_7\
        );

    \I__7364\ : InMux
    port map (
            O => \N__37181\,
            I => \N__37178\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__37178\,
            I => \N__37175\
        );

    \I__7362\ : Odrv12
    port map (
            O => \N__37175\,
            I => \sDAC_mem_pointerZ0Z_6\
        );

    \I__7361\ : InMux
    port map (
            O => \N__37172\,
            I => \N__37169\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__37169\,
            I => un17_sdacdyn_0
        );

    \I__7359\ : InMux
    port map (
            O => \N__37166\,
            I => \N__37163\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__37163\,
            I => \N__37160\
        );

    \I__7357\ : Span4Mux_v
    port map (
            O => \N__37160\,
            I => \N__37157\
        );

    \I__7356\ : Odrv4
    port map (
            O => \N__37157\,
            I => \sDAC_data_RNO_5Z0Z_5\
        );

    \I__7355\ : InMux
    port map (
            O => \N__37154\,
            I => \N__37151\
        );

    \I__7354\ : LocalMux
    port map (
            O => \N__37151\,
            I => \sDAC_data_RNO_2Z0Z_5\
        );

    \I__7353\ : CascadeMux
    port map (
            O => \N__37148\,
            I => \sDAC_data_RNO_1Z0Z_5_cascade_\
        );

    \I__7352\ : InMux
    port map (
            O => \N__37145\,
            I => \N__37142\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__37142\,
            I => \N__37139\
        );

    \I__7350\ : Span4Mux_v
    port map (
            O => \N__37139\,
            I => \N__37136\
        );

    \I__7349\ : Span4Mux_v
    port map (
            O => \N__37136\,
            I => \N__37133\
        );

    \I__7348\ : Odrv4
    port map (
            O => \N__37133\,
            I => \sEEDACZ0Z_2\
        );

    \I__7347\ : CascadeMux
    port map (
            O => \N__37130\,
            I => \sDAC_data_2_5_cascade_\
        );

    \I__7346\ : InMux
    port map (
            O => \N__37127\,
            I => \N__37124\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__37124\,
            I => \N__37121\
        );

    \I__7344\ : Span4Mux_h
    port map (
            O => \N__37121\,
            I => \N__37118\
        );

    \I__7343\ : Span4Mux_v
    port map (
            O => \N__37118\,
            I => \N__37115\
        );

    \I__7342\ : Span4Mux_h
    port map (
            O => \N__37115\,
            I => \N__37112\
        );

    \I__7341\ : Span4Mux_h
    port map (
            O => \N__37112\,
            I => \N__37109\
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__37109\,
            I => \sDAC_dataZ0Z_5\
        );

    \I__7339\ : InMux
    port map (
            O => \N__37106\,
            I => \N__37103\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__37103\,
            I => \sDAC_data_RNO_15Z0Z_5\
        );

    \I__7337\ : InMux
    port map (
            O => \N__37100\,
            I => \N__37097\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__37097\,
            I => \sDAC_data_2_14_ns_1_5\
        );

    \I__7335\ : InMux
    port map (
            O => \N__37094\,
            I => \N__37091\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__37091\,
            I => \sDAC_data_RNO_29Z0Z_5\
        );

    \I__7333\ : InMux
    port map (
            O => \N__37088\,
            I => \N__37085\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__37085\,
            I => \N__37082\
        );

    \I__7331\ : Span4Mux_h
    port map (
            O => \N__37082\,
            I => \N__37079\
        );

    \I__7330\ : Span4Mux_v
    port map (
            O => \N__37079\,
            I => \N__37076\
        );

    \I__7329\ : Odrv4
    port map (
            O => \N__37076\,
            I => \sDAC_data_RNO_28Z0Z_5\
        );

    \I__7328\ : InMux
    port map (
            O => \N__37073\,
            I => \N__37070\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__37070\,
            I => \N__37067\
        );

    \I__7326\ : Odrv4
    port map (
            O => \N__37067\,
            I => \sDAC_data_RNO_20Z0Z_5\
        );

    \I__7325\ : CascadeMux
    port map (
            O => \N__37064\,
            I => \sDAC_data_2_32_ns_1_5_cascade_\
        );

    \I__7324\ : InMux
    port map (
            O => \N__37061\,
            I => \N__37058\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__37058\,
            I => \N__37055\
        );

    \I__7322\ : Span4Mux_h
    port map (
            O => \N__37055\,
            I => \N__37052\
        );

    \I__7321\ : Odrv4
    port map (
            O => \N__37052\,
            I => \sDAC_data_RNO_21Z0Z_5\
        );

    \I__7320\ : CascadeMux
    port map (
            O => \N__37049\,
            I => \sDAC_data_RNO_10Z0Z_5_cascade_\
        );

    \I__7319\ : InMux
    port map (
            O => \N__37046\,
            I => \N__37043\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__37043\,
            I => \sDAC_data_2_41_ns_1_5\
        );

    \I__7317\ : InMux
    port map (
            O => \N__37040\,
            I => \N__37037\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__37037\,
            I => \N__37034\
        );

    \I__7315\ : Span4Mux_h
    port map (
            O => \N__37034\,
            I => \N__37031\
        );

    \I__7314\ : Odrv4
    port map (
            O => \N__37031\,
            I => \sDAC_mem_9Z0Z_6\
        );

    \I__7313\ : InMux
    port map (
            O => \N__37028\,
            I => \N__37025\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__37025\,
            I => \N__37022\
        );

    \I__7311\ : Span4Mux_h
    port map (
            O => \N__37022\,
            I => \N__37019\
        );

    \I__7310\ : Odrv4
    port map (
            O => \N__37019\,
            I => \sDAC_mem_9Z0Z_7\
        );

    \I__7309\ : InMux
    port map (
            O => \N__37016\,
            I => \N__37013\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__7307\ : Odrv12
    port map (
            O => \N__37010\,
            I => \sDAC_mem_15Z0Z_6\
        );

    \I__7306\ : InMux
    port map (
            O => \N__37007\,
            I => \N__37004\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__37004\,
            I => \N__37001\
        );

    \I__7304\ : Span4Mux_h
    port map (
            O => \N__37001\,
            I => \N__36998\
        );

    \I__7303\ : Span4Mux_h
    port map (
            O => \N__36998\,
            I => \N__36995\
        );

    \I__7302\ : Odrv4
    port map (
            O => \N__36995\,
            I => \sDAC_mem_14Z0Z_6\
        );

    \I__7301\ : CascadeMux
    port map (
            O => \N__36992\,
            I => \sDAC_data_RNO_18Z0Z_9_cascade_\
        );

    \I__7300\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36986\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__36986\,
            I => \sDAC_data_RNO_19Z0Z_9\
        );

    \I__7298\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36980\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__36980\,
            I => \N__36977\
        );

    \I__7296\ : Span4Mux_h
    port map (
            O => \N__36977\,
            I => \N__36974\
        );

    \I__7295\ : Odrv4
    port map (
            O => \N__36974\,
            I => \sDAC_data_2_24_ns_1_9\
        );

    \I__7294\ : InMux
    port map (
            O => \N__36971\,
            I => \N__36968\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__36968\,
            I => \sDAC_mem_12Z0Z_6\
        );

    \I__7292\ : CEMux
    port map (
            O => \N__36965\,
            I => \N__36961\
        );

    \I__7291\ : CEMux
    port map (
            O => \N__36964\,
            I => \N__36956\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__36961\,
            I => \N__36953\
        );

    \I__7289\ : CEMux
    port map (
            O => \N__36960\,
            I => \N__36949\
        );

    \I__7288\ : CEMux
    port map (
            O => \N__36959\,
            I => \N__36946\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__36956\,
            I => \N__36943\
        );

    \I__7286\ : Span4Mux_h
    port map (
            O => \N__36953\,
            I => \N__36940\
        );

    \I__7285\ : CEMux
    port map (
            O => \N__36952\,
            I => \N__36937\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__36949\,
            I => \N__36934\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__36946\,
            I => \N__36931\
        );

    \I__7282\ : Span4Mux_h
    port map (
            O => \N__36943\,
            I => \N__36924\
        );

    \I__7281\ : Span4Mux_v
    port map (
            O => \N__36940\,
            I => \N__36924\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__36937\,
            I => \N__36924\
        );

    \I__7279\ : Span4Mux_v
    port map (
            O => \N__36934\,
            I => \N__36921\
        );

    \I__7278\ : Span4Mux_h
    port map (
            O => \N__36931\,
            I => \N__36918\
        );

    \I__7277\ : Span4Mux_h
    port map (
            O => \N__36924\,
            I => \N__36915\
        );

    \I__7276\ : Span4Mux_h
    port map (
            O => \N__36921\,
            I => \N__36910\
        );

    \I__7275\ : Span4Mux_h
    port map (
            O => \N__36918\,
            I => \N__36910\
        );

    \I__7274\ : Span4Mux_h
    port map (
            O => \N__36915\,
            I => \N__36907\
        );

    \I__7273\ : Odrv4
    port map (
            O => \N__36910\,
            I => \sDAC_mem_12_1_sqmuxa\
        );

    \I__7272\ : Odrv4
    port map (
            O => \N__36907\,
            I => \sDAC_mem_12_1_sqmuxa\
        );

    \I__7271\ : CascadeMux
    port map (
            O => \N__36902\,
            I => \op_le_op_le_un15_sdacdynlt4_cascade_\
        );

    \I__7270\ : InMux
    port map (
            O => \N__36899\,
            I => \N__36896\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__36896\,
            I => \N__36893\
        );

    \I__7268\ : Span4Mux_h
    port map (
            O => \N__36893\,
            I => \N__36890\
        );

    \I__7267\ : Sp12to4
    port map (
            O => \N__36890\,
            I => \N__36887\
        );

    \I__7266\ : Odrv12
    port map (
            O => \N__36887\,
            I => un17_sdacdyn_1
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__36884\,
            I => \sDAC_data_RNO_26Z0Z_7_cascade_\
        );

    \I__7264\ : InMux
    port map (
            O => \N__36881\,
            I => \N__36878\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__36878\,
            I => \N__36875\
        );

    \I__7262\ : Span4Mux_h
    port map (
            O => \N__36875\,
            I => \N__36872\
        );

    \I__7261\ : Odrv4
    port map (
            O => \N__36872\,
            I => \sDAC_data_RNO_14Z0Z_7\
        );

    \I__7260\ : InMux
    port map (
            O => \N__36869\,
            I => \N__36866\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__36866\,
            I => \sDAC_mem_32Z0Z_4\
        );

    \I__7258\ : CascadeMux
    port map (
            O => \N__36863\,
            I => \sDAC_data_RNO_26Z0Z_8_cascade_\
        );

    \I__7257\ : CascadeMux
    port map (
            O => \N__36860\,
            I => \N__36857\
        );

    \I__7256\ : InMux
    port map (
            O => \N__36857\,
            I => \N__36854\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__36854\,
            I => \N__36851\
        );

    \I__7254\ : Span4Mux_h
    port map (
            O => \N__36851\,
            I => \N__36848\
        );

    \I__7253\ : Odrv4
    port map (
            O => \N__36848\,
            I => \sDAC_data_RNO_14Z0Z_8\
        );

    \I__7252\ : InMux
    port map (
            O => \N__36845\,
            I => \N__36842\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__36842\,
            I => \N__36839\
        );

    \I__7250\ : Span4Mux_v
    port map (
            O => \N__36839\,
            I => \N__36836\
        );

    \I__7249\ : Odrv4
    port map (
            O => \N__36836\,
            I => \sDAC_mem_9Z0Z_0\
        );

    \I__7248\ : InMux
    port map (
            O => \N__36833\,
            I => \N__36830\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__36830\,
            I => \N__36827\
        );

    \I__7246\ : Span4Mux_h
    port map (
            O => \N__36827\,
            I => \N__36824\
        );

    \I__7245\ : Odrv4
    port map (
            O => \N__36824\,
            I => \sDAC_mem_9Z0Z_1\
        );

    \I__7244\ : InMux
    port map (
            O => \N__36821\,
            I => \N__36818\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__36818\,
            I => \sDAC_mem_9Z0Z_2\
        );

    \I__7242\ : InMux
    port map (
            O => \N__36815\,
            I => \N__36812\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__36812\,
            I => \N__36809\
        );

    \I__7240\ : Span4Mux_h
    port map (
            O => \N__36809\,
            I => \N__36806\
        );

    \I__7239\ : Span4Mux_h
    port map (
            O => \N__36806\,
            I => \N__36803\
        );

    \I__7238\ : Odrv4
    port map (
            O => \N__36803\,
            I => \sDAC_mem_9Z0Z_3\
        );

    \I__7237\ : InMux
    port map (
            O => \N__36800\,
            I => \N__36797\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__36797\,
            I => \N__36794\
        );

    \I__7235\ : Sp12to4
    port map (
            O => \N__36794\,
            I => \N__36791\
        );

    \I__7234\ : Odrv12
    port map (
            O => \N__36791\,
            I => \sDAC_mem_9Z0Z_4\
        );

    \I__7233\ : InMux
    port map (
            O => \N__36788\,
            I => \N__36785\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__36785\,
            I => \N__36782\
        );

    \I__7231\ : Span4Mux_v
    port map (
            O => \N__36782\,
            I => \N__36779\
        );

    \I__7230\ : Odrv4
    port map (
            O => \N__36779\,
            I => \sDAC_mem_9Z0Z_5\
        );

    \I__7229\ : InMux
    port map (
            O => \N__36776\,
            I => \N__36773\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__36773\,
            I => \N__36770\
        );

    \I__7227\ : Span4Mux_h
    port map (
            O => \N__36770\,
            I => \N__36767\
        );

    \I__7226\ : Odrv4
    port map (
            O => \N__36767\,
            I => \sDAC_mem_23Z0Z_3\
        );

    \I__7225\ : InMux
    port map (
            O => \N__36764\,
            I => \N__36761\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__36761\,
            I => \N__36758\
        );

    \I__7223\ : Span4Mux_v
    port map (
            O => \N__36758\,
            I => \N__36755\
        );

    \I__7222\ : Span4Mux_v
    port map (
            O => \N__36755\,
            I => \N__36752\
        );

    \I__7221\ : Span4Mux_v
    port map (
            O => \N__36752\,
            I => \N__36749\
        );

    \I__7220\ : Odrv4
    port map (
            O => \N__36749\,
            I => \sDAC_mem_23Z0Z_4\
        );

    \I__7219\ : InMux
    port map (
            O => \N__36746\,
            I => \N__36743\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__36743\,
            I => \N__36740\
        );

    \I__7217\ : Span4Mux_v
    port map (
            O => \N__36740\,
            I => \N__36737\
        );

    \I__7216\ : Sp12to4
    port map (
            O => \N__36737\,
            I => \N__36734\
        );

    \I__7215\ : Span12Mux_h
    port map (
            O => \N__36734\,
            I => \N__36731\
        );

    \I__7214\ : Odrv12
    port map (
            O => \N__36731\,
            I => \sDAC_mem_23Z0Z_5\
        );

    \I__7213\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36725\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__36725\,
            I => \N__36722\
        );

    \I__7211\ : Span12Mux_v
    port map (
            O => \N__36722\,
            I => \N__36719\
        );

    \I__7210\ : Odrv12
    port map (
            O => \N__36719\,
            I => \sDAC_mem_23Z0Z_6\
        );

    \I__7209\ : InMux
    port map (
            O => \N__36716\,
            I => \N__36713\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__36713\,
            I => \N__36710\
        );

    \I__7207\ : Span4Mux_h
    port map (
            O => \N__36710\,
            I => \N__36707\
        );

    \I__7206\ : Span4Mux_v
    port map (
            O => \N__36707\,
            I => \N__36704\
        );

    \I__7205\ : Odrv4
    port map (
            O => \N__36704\,
            I => \sDAC_mem_23Z0Z_7\
        );

    \I__7204\ : CEMux
    port map (
            O => \N__36701\,
            I => \N__36698\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__36698\,
            I => \N__36695\
        );

    \I__7202\ : Span4Mux_v
    port map (
            O => \N__36695\,
            I => \N__36692\
        );

    \I__7201\ : Span4Mux_h
    port map (
            O => \N__36692\,
            I => \N__36689\
        );

    \I__7200\ : Span4Mux_h
    port map (
            O => \N__36689\,
            I => \N__36686\
        );

    \I__7199\ : Odrv4
    port map (
            O => \N__36686\,
            I => \sDAC_mem_23_1_sqmuxa\
        );

    \I__7198\ : CascadeMux
    port map (
            O => \N__36683\,
            I => \sDAC_data_RNO_26Z0Z_6_cascade_\
        );

    \I__7197\ : InMux
    port map (
            O => \N__36680\,
            I => \N__36677\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__36677\,
            I => \sDAC_mem_32Z0Z_3\
        );

    \I__7195\ : InMux
    port map (
            O => \N__36674\,
            I => \N__36671\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__36671\,
            I => \N__36668\
        );

    \I__7193\ : Span4Mux_v
    port map (
            O => \N__36668\,
            I => \N__36665\
        );

    \I__7192\ : Odrv4
    port map (
            O => \N__36665\,
            I => \sDAC_data_RNO_14Z0Z_6\
        );

    \I__7191\ : InMux
    port map (
            O => \N__36662\,
            I => \N__36659\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__36659\,
            I => \N__36656\
        );

    \I__7189\ : Odrv4
    port map (
            O => \N__36656\,
            I => \sDAC_mem_20Z0Z_4\
        );

    \I__7188\ : InMux
    port map (
            O => \N__36653\,
            I => \N__36650\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__36650\,
            I => \N__36647\
        );

    \I__7186\ : Sp12to4
    port map (
            O => \N__36647\,
            I => \N__36644\
        );

    \I__7185\ : Span12Mux_v
    port map (
            O => \N__36644\,
            I => \N__36641\
        );

    \I__7184\ : Odrv12
    port map (
            O => \N__36641\,
            I => \sDAC_mem_20Z0Z_7\
        );

    \I__7183\ : CEMux
    port map (
            O => \N__36638\,
            I => \N__36634\
        );

    \I__7182\ : CEMux
    port map (
            O => \N__36637\,
            I => \N__36631\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__36634\,
            I => \N__36628\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__36631\,
            I => \N__36625\
        );

    \I__7179\ : Span4Mux_h
    port map (
            O => \N__36628\,
            I => \N__36622\
        );

    \I__7178\ : Span12Mux_v
    port map (
            O => \N__36625\,
            I => \N__36619\
        );

    \I__7177\ : Span4Mux_v
    port map (
            O => \N__36622\,
            I => \N__36616\
        );

    \I__7176\ : Odrv12
    port map (
            O => \N__36619\,
            I => \sDAC_mem_20_1_sqmuxa\
        );

    \I__7175\ : Odrv4
    port map (
            O => \N__36616\,
            I => \sDAC_mem_20_1_sqmuxa\
        );

    \I__7174\ : InMux
    port map (
            O => \N__36611\,
            I => \N__36608\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__36608\,
            I => \N__36605\
        );

    \I__7172\ : Span4Mux_h
    port map (
            O => \N__36605\,
            I => \N__36602\
        );

    \I__7171\ : Span4Mux_v
    port map (
            O => \N__36602\,
            I => \N__36599\
        );

    \I__7170\ : Odrv4
    port map (
            O => \N__36599\,
            I => \sDAC_mem_6Z0Z_0\
        );

    \I__7169\ : InMux
    port map (
            O => \N__36596\,
            I => \N__36593\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__36593\,
            I => \N__36590\
        );

    \I__7167\ : Span4Mux_h
    port map (
            O => \N__36590\,
            I => \N__36587\
        );

    \I__7166\ : Span4Mux_v
    port map (
            O => \N__36587\,
            I => \N__36584\
        );

    \I__7165\ : Odrv4
    port map (
            O => \N__36584\,
            I => \sDAC_mem_6Z0Z_1\
        );

    \I__7164\ : InMux
    port map (
            O => \N__36581\,
            I => \N__36578\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__36578\,
            I => \N__36575\
        );

    \I__7162\ : Span4Mux_h
    port map (
            O => \N__36575\,
            I => \N__36572\
        );

    \I__7161\ : Odrv4
    port map (
            O => \N__36572\,
            I => \sDAC_mem_6Z0Z_4\
        );

    \I__7160\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36566\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__36566\,
            I => \N__36563\
        );

    \I__7158\ : Span4Mux_h
    port map (
            O => \N__36563\,
            I => \N__36560\
        );

    \I__7157\ : Span4Mux_v
    port map (
            O => \N__36560\,
            I => \N__36557\
        );

    \I__7156\ : Odrv4
    port map (
            O => \N__36557\,
            I => \sDAC_mem_6Z0Z_7\
        );

    \I__7155\ : CEMux
    port map (
            O => \N__36554\,
            I => \N__36550\
        );

    \I__7154\ : CEMux
    port map (
            O => \N__36553\,
            I => \N__36546\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__36550\,
            I => \N__36543\
        );

    \I__7152\ : CEMux
    port map (
            O => \N__36549\,
            I => \N__36540\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__36546\,
            I => \N__36537\
        );

    \I__7150\ : Span4Mux_v
    port map (
            O => \N__36543\,
            I => \N__36532\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__36540\,
            I => \N__36532\
        );

    \I__7148\ : Span4Mux_v
    port map (
            O => \N__36537\,
            I => \N__36529\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__36532\,
            I => \N__36526\
        );

    \I__7146\ : Span4Mux_h
    port map (
            O => \N__36529\,
            I => \N__36523\
        );

    \I__7145\ : Span4Mux_h
    port map (
            O => \N__36526\,
            I => \N__36520\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__36523\,
            I => \sDAC_mem_6_1_sqmuxa\
        );

    \I__7143\ : Odrv4
    port map (
            O => \N__36520\,
            I => \sDAC_mem_6_1_sqmuxa\
        );

    \I__7142\ : InMux
    port map (
            O => \N__36515\,
            I => \N__36512\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__36512\,
            I => \N__36509\
        );

    \I__7140\ : Span4Mux_h
    port map (
            O => \N__36509\,
            I => \N__36506\
        );

    \I__7139\ : Odrv4
    port map (
            O => \N__36506\,
            I => \sDAC_mem_23Z0Z_0\
        );

    \I__7138\ : InMux
    port map (
            O => \N__36503\,
            I => \N__36500\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__36500\,
            I => \N__36497\
        );

    \I__7136\ : Span4Mux_v
    port map (
            O => \N__36497\,
            I => \N__36494\
        );

    \I__7135\ : Odrv4
    port map (
            O => \N__36494\,
            I => \sDAC_mem_23Z0Z_1\
        );

    \I__7134\ : InMux
    port map (
            O => \N__36491\,
            I => \N__36488\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__36488\,
            I => \N__36485\
        );

    \I__7132\ : Span4Mux_h
    port map (
            O => \N__36485\,
            I => \N__36482\
        );

    \I__7131\ : Odrv4
    port map (
            O => \N__36482\,
            I => \sDAC_mem_23Z0Z_2\
        );

    \I__7130\ : CascadeMux
    port map (
            O => \N__36479\,
            I => \N__36476\
        );

    \I__7129\ : InMux
    port map (
            O => \N__36476\,
            I => \N__36473\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__36473\,
            I => \N__36470\
        );

    \I__7127\ : Span4Mux_h
    port map (
            O => \N__36470\,
            I => \N__36467\
        );

    \I__7126\ : Span4Mux_v
    port map (
            O => \N__36467\,
            I => \N__36464\
        );

    \I__7125\ : Odrv4
    port map (
            O => \N__36464\,
            I => \sDAC_mem_4Z0Z_5\
        );

    \I__7124\ : InMux
    port map (
            O => \N__36461\,
            I => \N__36458\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__36458\,
            I => \N__36455\
        );

    \I__7122\ : Sp12to4
    port map (
            O => \N__36455\,
            I => \N__36452\
        );

    \I__7121\ : Odrv12
    port map (
            O => \N__36452\,
            I => \sDAC_mem_4Z0Z_7\
        );

    \I__7120\ : InMux
    port map (
            O => \N__36449\,
            I => \N__36446\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__36446\,
            I => \N__36443\
        );

    \I__7118\ : Span4Mux_v
    port map (
            O => \N__36443\,
            I => \N__36440\
        );

    \I__7117\ : Odrv4
    port map (
            O => \N__36440\,
            I => \sDAC_mem_20Z0Z_0\
        );

    \I__7116\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36434\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__36434\,
            I => \N__36431\
        );

    \I__7114\ : Span4Mux_v
    port map (
            O => \N__36431\,
            I => \N__36428\
        );

    \I__7113\ : Odrv4
    port map (
            O => \N__36428\,
            I => \sDAC_mem_20Z0Z_1\
        );

    \I__7112\ : InMux
    port map (
            O => \N__36425\,
            I => \N__36422\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__36422\,
            I => \N__36419\
        );

    \I__7110\ : Span4Mux_h
    port map (
            O => \N__36419\,
            I => \N__36416\
        );

    \I__7109\ : Odrv4
    port map (
            O => \N__36416\,
            I => \sDAC_mem_20Z0Z_2\
        );

    \I__7108\ : InMux
    port map (
            O => \N__36413\,
            I => \N__36410\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__36410\,
            I => \N__36407\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__36407\,
            I => \sDAC_mem_20Z0Z_3\
        );

    \I__7105\ : InMux
    port map (
            O => \N__36404\,
            I => \N__36401\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__36401\,
            I => \N__36398\
        );

    \I__7103\ : Span4Mux_h
    port map (
            O => \N__36398\,
            I => \N__36395\
        );

    \I__7102\ : Sp12to4
    port map (
            O => \N__36395\,
            I => \N__36392\
        );

    \I__7101\ : Span12Mux_v
    port map (
            O => \N__36392\,
            I => \N__36389\
        );

    \I__7100\ : Span12Mux_h
    port map (
            O => \N__36389\,
            I => \N__36385\
        );

    \I__7099\ : InMux
    port map (
            O => \N__36388\,
            I => \N__36382\
        );

    \I__7098\ : Odrv12
    port map (
            O => \N__36385\,
            I => \sRAM_pointer_writeZ0Z_17\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__36382\,
            I => \sRAM_pointer_writeZ0Z_17\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__36377\,
            I => \N__36374\
        );

    \I__7095\ : InMux
    port map (
            O => \N__36374\,
            I => \N__36371\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__36371\,
            I => \N__36368\
        );

    \I__7093\ : Span4Mux_h
    port map (
            O => \N__36368\,
            I => \N__36364\
        );

    \I__7092\ : InMux
    port map (
            O => \N__36367\,
            I => \N__36361\
        );

    \I__7091\ : Odrv4
    port map (
            O => \N__36364\,
            I => \sRAM_pointer_readZ0Z_17\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__36361\,
            I => \sRAM_pointer_readZ0Z_17\
        );

    \I__7089\ : IoInMux
    port map (
            O => \N__36356\,
            I => \N__36353\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__36353\,
            I => \N__36350\
        );

    \I__7087\ : IoSpan4Mux
    port map (
            O => \N__36350\,
            I => \N__36347\
        );

    \I__7086\ : Span4Mux_s3_h
    port map (
            O => \N__36347\,
            I => \N__36344\
        );

    \I__7085\ : Sp12to4
    port map (
            O => \N__36344\,
            I => \N__36341\
        );

    \I__7084\ : Odrv12
    port map (
            O => \N__36341\,
            I => \RAM_ADD_c_17\
        );

    \I__7083\ : InMux
    port map (
            O => \N__36338\,
            I => \N__36335\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__36335\,
            I => \N__36332\
        );

    \I__7081\ : Span4Mux_v
    port map (
            O => \N__36332\,
            I => \N__36329\
        );

    \I__7080\ : Span4Mux_v
    port map (
            O => \N__36329\,
            I => \N__36326\
        );

    \I__7079\ : Sp12to4
    port map (
            O => \N__36326\,
            I => \N__36323\
        );

    \I__7078\ : Span12Mux_h
    port map (
            O => \N__36323\,
            I => \N__36319\
        );

    \I__7077\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36316\
        );

    \I__7076\ : Odrv12
    port map (
            O => \N__36319\,
            I => \sRAM_pointer_writeZ0Z_18\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__36316\,
            I => \sRAM_pointer_writeZ0Z_18\
        );

    \I__7074\ : CascadeMux
    port map (
            O => \N__36311\,
            I => \N__36308\
        );

    \I__7073\ : InMux
    port map (
            O => \N__36308\,
            I => \N__36305\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__36305\,
            I => \N__36302\
        );

    \I__7071\ : Span12Mux_h
    port map (
            O => \N__36302\,
            I => \N__36298\
        );

    \I__7070\ : InMux
    port map (
            O => \N__36301\,
            I => \N__36295\
        );

    \I__7069\ : Odrv12
    port map (
            O => \N__36298\,
            I => \sRAM_pointer_readZ0Z_18\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__36295\,
            I => \sRAM_pointer_readZ0Z_18\
        );

    \I__7067\ : IoInMux
    port map (
            O => \N__36290\,
            I => \N__36287\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__36287\,
            I => \N__36284\
        );

    \I__7065\ : IoSpan4Mux
    port map (
            O => \N__36284\,
            I => \N__36281\
        );

    \I__7064\ : Span4Mux_s1_h
    port map (
            O => \N__36281\,
            I => \N__36278\
        );

    \I__7063\ : Sp12to4
    port map (
            O => \N__36278\,
            I => \N__36275\
        );

    \I__7062\ : Span12Mux_h
    port map (
            O => \N__36275\,
            I => \N__36272\
        );

    \I__7061\ : Span12Mux_v
    port map (
            O => \N__36272\,
            I => \N__36269\
        );

    \I__7060\ : Odrv12
    port map (
            O => \N__36269\,
            I => \RAM_ADD_c_18\
        );

    \I__7059\ : InMux
    port map (
            O => \N__36266\,
            I => \N__36263\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__36263\,
            I => \N__36260\
        );

    \I__7057\ : Span4Mux_v
    port map (
            O => \N__36260\,
            I => \N__36257\
        );

    \I__7056\ : Span4Mux_h
    port map (
            O => \N__36257\,
            I => \N__36254\
        );

    \I__7055\ : Sp12to4
    port map (
            O => \N__36254\,
            I => \N__36251\
        );

    \I__7054\ : Span12Mux_h
    port map (
            O => \N__36251\,
            I => \N__36247\
        );

    \I__7053\ : InMux
    port map (
            O => \N__36250\,
            I => \N__36244\
        );

    \I__7052\ : Odrv12
    port map (
            O => \N__36247\,
            I => \sRAM_pointer_writeZ0Z_9\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__36244\,
            I => \sRAM_pointer_writeZ0Z_9\
        );

    \I__7050\ : CascadeMux
    port map (
            O => \N__36239\,
            I => \N__36236\
        );

    \I__7049\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36233\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__36233\,
            I => \N__36230\
        );

    \I__7047\ : Span4Mux_v
    port map (
            O => \N__36230\,
            I => \N__36226\
        );

    \I__7046\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36223\
        );

    \I__7045\ : Odrv4
    port map (
            O => \N__36226\,
            I => \sRAM_pointer_readZ0Z_9\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__36223\,
            I => \sRAM_pointer_readZ0Z_9\
        );

    \I__7043\ : IoInMux
    port map (
            O => \N__36218\,
            I => \N__36215\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__36215\,
            I => \N__36212\
        );

    \I__7041\ : Span4Mux_s3_h
    port map (
            O => \N__36212\,
            I => \N__36209\
        );

    \I__7040\ : Span4Mux_h
    port map (
            O => \N__36209\,
            I => \N__36206\
        );

    \I__7039\ : Span4Mux_h
    port map (
            O => \N__36206\,
            I => \N__36203\
        );

    \I__7038\ : Span4Mux_v
    port map (
            O => \N__36203\,
            I => \N__36200\
        );

    \I__7037\ : Odrv4
    port map (
            O => \N__36200\,
            I => \RAM_ADD_c_9\
        );

    \I__7036\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36194\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__36194\,
            I => \N__36191\
        );

    \I__7034\ : Span4Mux_h
    port map (
            O => \N__36191\,
            I => \N__36188\
        );

    \I__7033\ : Span4Mux_h
    port map (
            O => \N__36188\,
            I => \N__36185\
        );

    \I__7032\ : Sp12to4
    port map (
            O => \N__36185\,
            I => \N__36182\
        );

    \I__7031\ : Span12Mux_v
    port map (
            O => \N__36182\,
            I => \N__36178\
        );

    \I__7030\ : InMux
    port map (
            O => \N__36181\,
            I => \N__36175\
        );

    \I__7029\ : Odrv12
    port map (
            O => \N__36178\,
            I => \sRAM_pointer_writeZ0Z_7\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__36175\,
            I => \sRAM_pointer_writeZ0Z_7\
        );

    \I__7027\ : CascadeMux
    port map (
            O => \N__36170\,
            I => \N__36167\
        );

    \I__7026\ : InMux
    port map (
            O => \N__36167\,
            I => \N__36164\
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__36164\,
            I => \N__36160\
        );

    \I__7024\ : InMux
    port map (
            O => \N__36163\,
            I => \N__36157\
        );

    \I__7023\ : Odrv12
    port map (
            O => \N__36160\,
            I => \sRAM_pointer_readZ0Z_7\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__36157\,
            I => \sRAM_pointer_readZ0Z_7\
        );

    \I__7021\ : IoInMux
    port map (
            O => \N__36152\,
            I => \N__36149\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__36149\,
            I => \N__36146\
        );

    \I__7019\ : Span4Mux_s0_h
    port map (
            O => \N__36146\,
            I => \N__36143\
        );

    \I__7018\ : Sp12to4
    port map (
            O => \N__36143\,
            I => \N__36140\
        );

    \I__7017\ : Span12Mux_s8_v
    port map (
            O => \N__36140\,
            I => \N__36137\
        );

    \I__7016\ : Odrv12
    port map (
            O => \N__36137\,
            I => \RAM_ADD_c_7\
        );

    \I__7015\ : InMux
    port map (
            O => \N__36134\,
            I => \N__36131\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__36131\,
            I => \N__36127\
        );

    \I__7013\ : InMux
    port map (
            O => \N__36130\,
            I => \N__36124\
        );

    \I__7012\ : Odrv4
    port map (
            O => \N__36127\,
            I => \sRAM_pointer_readZ0Z_2\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__36124\,
            I => \sRAM_pointer_readZ0Z_2\
        );

    \I__7010\ : CascadeMux
    port map (
            O => \N__36119\,
            I => \N__36116\
        );

    \I__7009\ : InMux
    port map (
            O => \N__36116\,
            I => \N__36113\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__36113\,
            I => \N__36110\
        );

    \I__7007\ : Span4Mux_v
    port map (
            O => \N__36110\,
            I => \N__36107\
        );

    \I__7006\ : Span4Mux_h
    port map (
            O => \N__36107\,
            I => \N__36104\
        );

    \I__7005\ : Sp12to4
    port map (
            O => \N__36104\,
            I => \N__36101\
        );

    \I__7004\ : Span12Mux_h
    port map (
            O => \N__36101\,
            I => \N__36097\
        );

    \I__7003\ : InMux
    port map (
            O => \N__36100\,
            I => \N__36094\
        );

    \I__7002\ : Odrv12
    port map (
            O => \N__36097\,
            I => \sRAM_pointer_writeZ0Z_2\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__36094\,
            I => \sRAM_pointer_writeZ0Z_2\
        );

    \I__7000\ : IoInMux
    port map (
            O => \N__36089\,
            I => \N__36086\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__36086\,
            I => \N__36083\
        );

    \I__6998\ : Span4Mux_s2_v
    port map (
            O => \N__36083\,
            I => \N__36080\
        );

    \I__6997\ : Span4Mux_v
    port map (
            O => \N__36080\,
            I => \N__36077\
        );

    \I__6996\ : Odrv4
    port map (
            O => \N__36077\,
            I => \RAM_ADD_c_2\
        );

    \I__6995\ : InMux
    port map (
            O => \N__36074\,
            I => \N__36071\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__36071\,
            I => \N__36068\
        );

    \I__6993\ : Span4Mux_v
    port map (
            O => \N__36068\,
            I => \N__36065\
        );

    \I__6992\ : Span4Mux_h
    port map (
            O => \N__36065\,
            I => \N__36062\
        );

    \I__6991\ : Sp12to4
    port map (
            O => \N__36062\,
            I => \N__36059\
        );

    \I__6990\ : Span12Mux_h
    port map (
            O => \N__36059\,
            I => \N__36055\
        );

    \I__6989\ : InMux
    port map (
            O => \N__36058\,
            I => \N__36052\
        );

    \I__6988\ : Odrv12
    port map (
            O => \N__36055\,
            I => \sRAM_pointer_writeZ0Z_1\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__36052\,
            I => \sRAM_pointer_writeZ0Z_1\
        );

    \I__6986\ : CascadeMux
    port map (
            O => \N__36047\,
            I => \N__36044\
        );

    \I__6985\ : InMux
    port map (
            O => \N__36044\,
            I => \N__36041\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__36041\,
            I => \N__36037\
        );

    \I__6983\ : InMux
    port map (
            O => \N__36040\,
            I => \N__36034\
        );

    \I__6982\ : Odrv4
    port map (
            O => \N__36037\,
            I => \sRAM_pointer_readZ0Z_1\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__36034\,
            I => \sRAM_pointer_readZ0Z_1\
        );

    \I__6980\ : IoInMux
    port map (
            O => \N__36029\,
            I => \N__36026\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__36026\,
            I => \N__36023\
        );

    \I__6978\ : Span12Mux_s2_v
    port map (
            O => \N__36023\,
            I => \N__36020\
        );

    \I__6977\ : Odrv12
    port map (
            O => \N__36020\,
            I => \RAM_ADD_c_1\
        );

    \I__6976\ : InMux
    port map (
            O => \N__36017\,
            I => \N__36014\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__36014\,
            I => \N__36011\
        );

    \I__6974\ : Span4Mux_v
    port map (
            O => \N__36011\,
            I => \N__36008\
        );

    \I__6973\ : Span4Mux_h
    port map (
            O => \N__36008\,
            I => \N__36005\
        );

    \I__6972\ : Span4Mux_v
    port map (
            O => \N__36005\,
            I => \N__36002\
        );

    \I__6971\ : Sp12to4
    port map (
            O => \N__36002\,
            I => \N__35998\
        );

    \I__6970\ : InMux
    port map (
            O => \N__36001\,
            I => \N__35995\
        );

    \I__6969\ : Odrv12
    port map (
            O => \N__35998\,
            I => \sRAM_pointer_writeZ0Z_6\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__35995\,
            I => \sRAM_pointer_writeZ0Z_6\
        );

    \I__6967\ : CascadeMux
    port map (
            O => \N__35990\,
            I => \N__35987\
        );

    \I__6966\ : InMux
    port map (
            O => \N__35987\,
            I => \N__35984\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__35984\,
            I => \N__35980\
        );

    \I__6964\ : InMux
    port map (
            O => \N__35983\,
            I => \N__35977\
        );

    \I__6963\ : Odrv12
    port map (
            O => \N__35980\,
            I => \sRAM_pointer_readZ0Z_6\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__35977\,
            I => \sRAM_pointer_readZ0Z_6\
        );

    \I__6961\ : IoInMux
    port map (
            O => \N__35972\,
            I => \N__35969\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__35969\,
            I => \N__35966\
        );

    \I__6959\ : IoSpan4Mux
    port map (
            O => \N__35966\,
            I => \N__35963\
        );

    \I__6958\ : Span4Mux_s3_h
    port map (
            O => \N__35963\,
            I => \N__35960\
        );

    \I__6957\ : Span4Mux_h
    port map (
            O => \N__35960\,
            I => \N__35957\
        );

    \I__6956\ : Span4Mux_h
    port map (
            O => \N__35957\,
            I => \N__35954\
        );

    \I__6955\ : Odrv4
    port map (
            O => \N__35954\,
            I => \RAM_ADD_c_6\
        );

    \I__6954\ : InMux
    port map (
            O => \N__35951\,
            I => \N__35948\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__35948\,
            I => \N__35945\
        );

    \I__6952\ : Span4Mux_v
    port map (
            O => \N__35945\,
            I => \N__35942\
        );

    \I__6951\ : Span4Mux_h
    port map (
            O => \N__35942\,
            I => \N__35939\
        );

    \I__6950\ : Sp12to4
    port map (
            O => \N__35939\,
            I => \N__35936\
        );

    \I__6949\ : Span12Mux_h
    port map (
            O => \N__35936\,
            I => \N__35933\
        );

    \I__6948\ : Odrv12
    port map (
            O => \N__35933\,
            I => \ADC4_c\
        );

    \I__6947\ : IoInMux
    port map (
            O => \N__35930\,
            I => \N__35927\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__35927\,
            I => \N__35924\
        );

    \I__6945\ : Span4Mux_s2_v
    port map (
            O => \N__35924\,
            I => \N__35921\
        );

    \I__6944\ : Span4Mux_h
    port map (
            O => \N__35921\,
            I => \N__35918\
        );

    \I__6943\ : Span4Mux_h
    port map (
            O => \N__35918\,
            I => \N__35915\
        );

    \I__6942\ : Span4Mux_v
    port map (
            O => \N__35915\,
            I => \N__35912\
        );

    \I__6941\ : Odrv4
    port map (
            O => \N__35912\,
            I => \RAM_DATA_1Z0Z_4\
        );

    \I__6940\ : InMux
    port map (
            O => \N__35909\,
            I => \N__35906\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__35906\,
            I => \N__35903\
        );

    \I__6938\ : Span4Mux_v
    port map (
            O => \N__35903\,
            I => \N__35899\
        );

    \I__6937\ : InMux
    port map (
            O => \N__35902\,
            I => \N__35896\
        );

    \I__6936\ : Odrv4
    port map (
            O => \N__35899\,
            I => \sRAM_pointer_readZ0Z_0\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__35896\,
            I => \sRAM_pointer_readZ0Z_0\
        );

    \I__6934\ : CascadeMux
    port map (
            O => \N__35891\,
            I => \N__35888\
        );

    \I__6933\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35885\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__35885\,
            I => \N__35882\
        );

    \I__6931\ : Span4Mux_h
    port map (
            O => \N__35882\,
            I => \N__35879\
        );

    \I__6930\ : Sp12to4
    port map (
            O => \N__35879\,
            I => \N__35876\
        );

    \I__6929\ : Span12Mux_s7_v
    port map (
            O => \N__35876\,
            I => \N__35873\
        );

    \I__6928\ : Span12Mux_h
    port map (
            O => \N__35873\,
            I => \N__35869\
        );

    \I__6927\ : InMux
    port map (
            O => \N__35872\,
            I => \N__35866\
        );

    \I__6926\ : Odrv12
    port map (
            O => \N__35869\,
            I => \sRAM_pointer_writeZ0Z_0\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__35866\,
            I => \sRAM_pointer_writeZ0Z_0\
        );

    \I__6924\ : IoInMux
    port map (
            O => \N__35861\,
            I => \N__35858\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__35858\,
            I => \N__35855\
        );

    \I__6922\ : IoSpan4Mux
    port map (
            O => \N__35855\,
            I => \N__35852\
        );

    \I__6921\ : Sp12to4
    port map (
            O => \N__35852\,
            I => \N__35849\
        );

    \I__6920\ : Odrv12
    port map (
            O => \N__35849\,
            I => \RAM_ADD_c_0\
        );

    \I__6919\ : InMux
    port map (
            O => \N__35846\,
            I => \N__35843\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__35843\,
            I => \N__35840\
        );

    \I__6917\ : Span4Mux_v
    port map (
            O => \N__35840\,
            I => \N__35836\
        );

    \I__6916\ : InMux
    port map (
            O => \N__35839\,
            I => \N__35833\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__35836\,
            I => \sRAM_pointer_readZ0Z_10\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__35833\,
            I => \sRAM_pointer_readZ0Z_10\
        );

    \I__6913\ : InMux
    port map (
            O => \N__35828\,
            I => \N__35825\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__35825\,
            I => \N__35822\
        );

    \I__6911\ : Span4Mux_v
    port map (
            O => \N__35822\,
            I => \N__35819\
        );

    \I__6910\ : Span4Mux_h
    port map (
            O => \N__35819\,
            I => \N__35816\
        );

    \I__6909\ : Span4Mux_h
    port map (
            O => \N__35816\,
            I => \N__35813\
        );

    \I__6908\ : Span4Mux_h
    port map (
            O => \N__35813\,
            I => \N__35810\
        );

    \I__6907\ : Span4Mux_h
    port map (
            O => \N__35810\,
            I => \N__35806\
        );

    \I__6906\ : InMux
    port map (
            O => \N__35809\,
            I => \N__35803\
        );

    \I__6905\ : Odrv4
    port map (
            O => \N__35806\,
            I => \sRAM_pointer_writeZ0Z_10\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__35803\,
            I => \sRAM_pointer_writeZ0Z_10\
        );

    \I__6903\ : IoInMux
    port map (
            O => \N__35798\,
            I => \N__35795\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__35795\,
            I => \N__35792\
        );

    \I__6901\ : IoSpan4Mux
    port map (
            O => \N__35792\,
            I => \N__35789\
        );

    \I__6900\ : Span4Mux_s1_h
    port map (
            O => \N__35789\,
            I => \N__35786\
        );

    \I__6899\ : Sp12to4
    port map (
            O => \N__35786\,
            I => \N__35783\
        );

    \I__6898\ : Span12Mux_h
    port map (
            O => \N__35783\,
            I => \N__35780\
        );

    \I__6897\ : Span12Mux_v
    port map (
            O => \N__35780\,
            I => \N__35777\
        );

    \I__6896\ : Odrv12
    port map (
            O => \N__35777\,
            I => \RAM_ADD_c_10\
        );

    \I__6895\ : InMux
    port map (
            O => \N__35774\,
            I => \N__35771\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__35771\,
            I => \N__35768\
        );

    \I__6893\ : Span4Mux_v
    port map (
            O => \N__35768\,
            I => \N__35764\
        );

    \I__6892\ : InMux
    port map (
            O => \N__35767\,
            I => \N__35761\
        );

    \I__6891\ : Odrv4
    port map (
            O => \N__35764\,
            I => \sRAM_pointer_readZ0Z_11\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__35761\,
            I => \sRAM_pointer_readZ0Z_11\
        );

    \I__6889\ : CascadeMux
    port map (
            O => \N__35756\,
            I => \N__35753\
        );

    \I__6888\ : InMux
    port map (
            O => \N__35753\,
            I => \N__35750\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__35750\,
            I => \N__35747\
        );

    \I__6886\ : Span4Mux_v
    port map (
            O => \N__35747\,
            I => \N__35744\
        );

    \I__6885\ : Span4Mux_h
    port map (
            O => \N__35744\,
            I => \N__35741\
        );

    \I__6884\ : Sp12to4
    port map (
            O => \N__35741\,
            I => \N__35738\
        );

    \I__6883\ : Span12Mux_h
    port map (
            O => \N__35738\,
            I => \N__35734\
        );

    \I__6882\ : InMux
    port map (
            O => \N__35737\,
            I => \N__35731\
        );

    \I__6881\ : Odrv12
    port map (
            O => \N__35734\,
            I => \sRAM_pointer_writeZ0Z_11\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__35731\,
            I => \sRAM_pointer_writeZ0Z_11\
        );

    \I__6879\ : IoInMux
    port map (
            O => \N__35726\,
            I => \N__35723\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__35723\,
            I => \N__35720\
        );

    \I__6877\ : Span4Mux_s0_h
    port map (
            O => \N__35720\,
            I => \N__35717\
        );

    \I__6876\ : Sp12to4
    port map (
            O => \N__35717\,
            I => \N__35714\
        );

    \I__6875\ : Span12Mux_v
    port map (
            O => \N__35714\,
            I => \N__35711\
        );

    \I__6874\ : Span12Mux_h
    port map (
            O => \N__35711\,
            I => \N__35708\
        );

    \I__6873\ : Odrv12
    port map (
            O => \N__35708\,
            I => \RAM_ADD_c_11\
        );

    \I__6872\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35702\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__35702\,
            I => \N__35699\
        );

    \I__6870\ : Span4Mux_v
    port map (
            O => \N__35699\,
            I => \N__35696\
        );

    \I__6869\ : Span4Mux_h
    port map (
            O => \N__35696\,
            I => \N__35693\
        );

    \I__6868\ : Sp12to4
    port map (
            O => \N__35693\,
            I => \N__35690\
        );

    \I__6867\ : Span12Mux_v
    port map (
            O => \N__35690\,
            I => \N__35686\
        );

    \I__6866\ : InMux
    port map (
            O => \N__35689\,
            I => \N__35683\
        );

    \I__6865\ : Odrv12
    port map (
            O => \N__35686\,
            I => \sRAM_pointer_writeZ0Z_12\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__35683\,
            I => \sRAM_pointer_writeZ0Z_12\
        );

    \I__6863\ : InMux
    port map (
            O => \N__35678\,
            I => \N__35675\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__35675\,
            I => \N__35672\
        );

    \I__6861\ : Span4Mux_v
    port map (
            O => \N__35672\,
            I => \N__35668\
        );

    \I__6860\ : InMux
    port map (
            O => \N__35671\,
            I => \N__35665\
        );

    \I__6859\ : Odrv4
    port map (
            O => \N__35668\,
            I => \sRAM_pointer_readZ0Z_12\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__35665\,
            I => \sRAM_pointer_readZ0Z_12\
        );

    \I__6857\ : IoInMux
    port map (
            O => \N__35660\,
            I => \N__35657\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__35657\,
            I => \N__35654\
        );

    \I__6855\ : Span4Mux_s0_h
    port map (
            O => \N__35654\,
            I => \N__35651\
        );

    \I__6854\ : Sp12to4
    port map (
            O => \N__35651\,
            I => \N__35648\
        );

    \I__6853\ : Span12Mux_v
    port map (
            O => \N__35648\,
            I => \N__35645\
        );

    \I__6852\ : Span12Mux_h
    port map (
            O => \N__35645\,
            I => \N__35642\
        );

    \I__6851\ : Odrv12
    port map (
            O => \N__35642\,
            I => \RAM_ADD_c_12\
        );

    \I__6850\ : InMux
    port map (
            O => \N__35639\,
            I => \N__35636\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__35636\,
            I => \N__35633\
        );

    \I__6848\ : Span4Mux_h
    port map (
            O => \N__35633\,
            I => \N__35629\
        );

    \I__6847\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35626\
        );

    \I__6846\ : Odrv4
    port map (
            O => \N__35629\,
            I => \sRAM_pointer_readZ0Z_13\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__35626\,
            I => \sRAM_pointer_readZ0Z_13\
        );

    \I__6844\ : CascadeMux
    port map (
            O => \N__35621\,
            I => \N__35618\
        );

    \I__6843\ : InMux
    port map (
            O => \N__35618\,
            I => \N__35615\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__35615\,
            I => \N__35612\
        );

    \I__6841\ : Span4Mux_h
    port map (
            O => \N__35612\,
            I => \N__35609\
        );

    \I__6840\ : Sp12to4
    port map (
            O => \N__35609\,
            I => \N__35606\
        );

    \I__6839\ : Span12Mux_h
    port map (
            O => \N__35606\,
            I => \N__35602\
        );

    \I__6838\ : InMux
    port map (
            O => \N__35605\,
            I => \N__35599\
        );

    \I__6837\ : Odrv12
    port map (
            O => \N__35602\,
            I => \sRAM_pointer_writeZ0Z_13\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__35599\,
            I => \sRAM_pointer_writeZ0Z_13\
        );

    \I__6835\ : IoInMux
    port map (
            O => \N__35594\,
            I => \N__35591\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__35591\,
            I => \N__35588\
        );

    \I__6833\ : Sp12to4
    port map (
            O => \N__35588\,
            I => \N__35585\
        );

    \I__6832\ : Span12Mux_h
    port map (
            O => \N__35585\,
            I => \N__35582\
        );

    \I__6831\ : Span12Mux_v
    port map (
            O => \N__35582\,
            I => \N__35579\
        );

    \I__6830\ : Odrv12
    port map (
            O => \N__35579\,
            I => \RAM_ADD_c_13\
        );

    \I__6829\ : InMux
    port map (
            O => \N__35576\,
            I => \N__35573\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__35573\,
            I => \N__35570\
        );

    \I__6827\ : Span4Mux_v
    port map (
            O => \N__35570\,
            I => \N__35567\
        );

    \I__6826\ : Span4Mux_h
    port map (
            O => \N__35567\,
            I => \N__35564\
        );

    \I__6825\ : Sp12to4
    port map (
            O => \N__35564\,
            I => \N__35561\
        );

    \I__6824\ : Span12Mux_h
    port map (
            O => \N__35561\,
            I => \N__35557\
        );

    \I__6823\ : InMux
    port map (
            O => \N__35560\,
            I => \N__35554\
        );

    \I__6822\ : Odrv12
    port map (
            O => \N__35557\,
            I => \sRAM_pointer_writeZ0Z_14\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__35554\,
            I => \sRAM_pointer_writeZ0Z_14\
        );

    \I__6820\ : InMux
    port map (
            O => \N__35549\,
            I => \N__35546\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__35546\,
            I => \N__35543\
        );

    \I__6818\ : Span4Mux_h
    port map (
            O => \N__35543\,
            I => \N__35540\
        );

    \I__6817\ : Span4Mux_h
    port map (
            O => \N__35540\,
            I => \N__35536\
        );

    \I__6816\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35533\
        );

    \I__6815\ : Odrv4
    port map (
            O => \N__35536\,
            I => \sRAM_pointer_readZ0Z_14\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__35533\,
            I => \sRAM_pointer_readZ0Z_14\
        );

    \I__6813\ : IoInMux
    port map (
            O => \N__35528\,
            I => \N__35525\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__35525\,
            I => \N__35522\
        );

    \I__6811\ : IoSpan4Mux
    port map (
            O => \N__35522\,
            I => \N__35519\
        );

    \I__6810\ : Span4Mux_s1_h
    port map (
            O => \N__35519\,
            I => \N__35516\
        );

    \I__6809\ : Sp12to4
    port map (
            O => \N__35516\,
            I => \N__35513\
        );

    \I__6808\ : Span12Mux_h
    port map (
            O => \N__35513\,
            I => \N__35510\
        );

    \I__6807\ : Span12Mux_v
    port map (
            O => \N__35510\,
            I => \N__35507\
        );

    \I__6806\ : Odrv12
    port map (
            O => \N__35507\,
            I => \RAM_ADD_c_14\
        );

    \I__6805\ : InMux
    port map (
            O => \N__35504\,
            I => \N__35501\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__35501\,
            I => \N__35498\
        );

    \I__6803\ : Span4Mux_h
    port map (
            O => \N__35498\,
            I => \N__35494\
        );

    \I__6802\ : InMux
    port map (
            O => \N__35497\,
            I => \N__35491\
        );

    \I__6801\ : Odrv4
    port map (
            O => \N__35494\,
            I => \sRAM_pointer_readZ0Z_15\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__35491\,
            I => \sRAM_pointer_readZ0Z_15\
        );

    \I__6799\ : CascadeMux
    port map (
            O => \N__35486\,
            I => \N__35483\
        );

    \I__6798\ : InMux
    port map (
            O => \N__35483\,
            I => \N__35480\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__35480\,
            I => \N__35477\
        );

    \I__6796\ : Span4Mux_v
    port map (
            O => \N__35477\,
            I => \N__35474\
        );

    \I__6795\ : Span4Mux_h
    port map (
            O => \N__35474\,
            I => \N__35471\
        );

    \I__6794\ : Span4Mux_h
    port map (
            O => \N__35471\,
            I => \N__35468\
        );

    \I__6793\ : Sp12to4
    port map (
            O => \N__35468\,
            I => \N__35465\
        );

    \I__6792\ : Span12Mux_h
    port map (
            O => \N__35465\,
            I => \N__35461\
        );

    \I__6791\ : InMux
    port map (
            O => \N__35464\,
            I => \N__35458\
        );

    \I__6790\ : Odrv12
    port map (
            O => \N__35461\,
            I => \sRAM_pointer_writeZ0Z_15\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__35458\,
            I => \sRAM_pointer_writeZ0Z_15\
        );

    \I__6788\ : IoInMux
    port map (
            O => \N__35453\,
            I => \N__35450\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__35450\,
            I => \N__35447\
        );

    \I__6786\ : IoSpan4Mux
    port map (
            O => \N__35447\,
            I => \N__35444\
        );

    \I__6785\ : Span4Mux_s2_h
    port map (
            O => \N__35444\,
            I => \N__35441\
        );

    \I__6784\ : Span4Mux_h
    port map (
            O => \N__35441\,
            I => \N__35438\
        );

    \I__6783\ : Span4Mux_h
    port map (
            O => \N__35438\,
            I => \N__35435\
        );

    \I__6782\ : Odrv4
    port map (
            O => \N__35435\,
            I => \RAM_ADD_c_15\
        );

    \I__6781\ : InMux
    port map (
            O => \N__35432\,
            I => \N__35429\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__35429\,
            I => \N__35426\
        );

    \I__6779\ : Span4Mux_h
    port map (
            O => \N__35426\,
            I => \N__35422\
        );

    \I__6778\ : InMux
    port map (
            O => \N__35425\,
            I => \N__35419\
        );

    \I__6777\ : Odrv4
    port map (
            O => \N__35422\,
            I => \sRAM_pointer_readZ0Z_16\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__35419\,
            I => \sRAM_pointer_readZ0Z_16\
        );

    \I__6775\ : CascadeMux
    port map (
            O => \N__35414\,
            I => \N__35411\
        );

    \I__6774\ : InMux
    port map (
            O => \N__35411\,
            I => \N__35408\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__35408\,
            I => \N__35405\
        );

    \I__6772\ : Span4Mux_v
    port map (
            O => \N__35405\,
            I => \N__35402\
        );

    \I__6771\ : Span4Mux_h
    port map (
            O => \N__35402\,
            I => \N__35399\
        );

    \I__6770\ : Span4Mux_h
    port map (
            O => \N__35399\,
            I => \N__35396\
        );

    \I__6769\ : Span4Mux_h
    port map (
            O => \N__35396\,
            I => \N__35392\
        );

    \I__6768\ : InMux
    port map (
            O => \N__35395\,
            I => \N__35389\
        );

    \I__6767\ : Span4Mux_h
    port map (
            O => \N__35392\,
            I => \N__35386\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__35389\,
            I => \sRAM_pointer_writeZ0Z_16\
        );

    \I__6765\ : Odrv4
    port map (
            O => \N__35386\,
            I => \sRAM_pointer_writeZ0Z_16\
        );

    \I__6764\ : IoInMux
    port map (
            O => \N__35381\,
            I => \N__35378\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__35378\,
            I => \N__35375\
        );

    \I__6762\ : IoSpan4Mux
    port map (
            O => \N__35375\,
            I => \N__35372\
        );

    \I__6761\ : Span4Mux_s1_h
    port map (
            O => \N__35372\,
            I => \N__35369\
        );

    \I__6760\ : Span4Mux_h
    port map (
            O => \N__35369\,
            I => \N__35366\
        );

    \I__6759\ : Span4Mux_h
    port map (
            O => \N__35366\,
            I => \N__35363\
        );

    \I__6758\ : Odrv4
    port map (
            O => \N__35363\,
            I => \RAM_ADD_c_16\
        );

    \I__6757\ : InMux
    port map (
            O => \N__35360\,
            I => \N__35356\
        );

    \I__6756\ : InMux
    port map (
            O => \N__35359\,
            I => \N__35353\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__35356\,
            I => \button_debounce_counterZ0Z_19\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__35353\,
            I => \button_debounce_counterZ0Z_19\
        );

    \I__6753\ : InMux
    port map (
            O => \N__35348\,
            I => un1_button_debounce_counter_cry_18
        );

    \I__6752\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35341\
        );

    \I__6751\ : InMux
    port map (
            O => \N__35344\,
            I => \N__35338\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__35341\,
            I => \button_debounce_counterZ0Z_20\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__35338\,
            I => \button_debounce_counterZ0Z_20\
        );

    \I__6748\ : InMux
    port map (
            O => \N__35333\,
            I => un1_button_debounce_counter_cry_19
        );

    \I__6747\ : CascadeMux
    port map (
            O => \N__35330\,
            I => \N__35326\
        );

    \I__6746\ : InMux
    port map (
            O => \N__35329\,
            I => \N__35323\
        );

    \I__6745\ : InMux
    port map (
            O => \N__35326\,
            I => \N__35320\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__35323\,
            I => \button_debounce_counterZ0Z_21\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__35320\,
            I => \button_debounce_counterZ0Z_21\
        );

    \I__6742\ : InMux
    port map (
            O => \N__35315\,
            I => un1_button_debounce_counter_cry_20
        );

    \I__6741\ : InMux
    port map (
            O => \N__35312\,
            I => \N__35309\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__35309\,
            I => \N__35306\
        );

    \I__6739\ : Span4Mux_v
    port map (
            O => \N__35306\,
            I => \N__35302\
        );

    \I__6738\ : InMux
    port map (
            O => \N__35305\,
            I => \N__35299\
        );

    \I__6737\ : Span4Mux_h
    port map (
            O => \N__35302\,
            I => \N__35296\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__35299\,
            I => \button_debounce_counterZ0Z_22\
        );

    \I__6735\ : Odrv4
    port map (
            O => \N__35296\,
            I => \button_debounce_counterZ0Z_22\
        );

    \I__6734\ : InMux
    port map (
            O => \N__35291\,
            I => un1_button_debounce_counter_cry_21
        );

    \I__6733\ : InMux
    port map (
            O => \N__35288\,
            I => \bfn_16_16_0_\
        );

    \I__6732\ : CascadeMux
    port map (
            O => \N__35285\,
            I => \N__35281\
        );

    \I__6731\ : InMux
    port map (
            O => \N__35284\,
            I => \N__35278\
        );

    \I__6730\ : InMux
    port map (
            O => \N__35281\,
            I => \N__35275\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__35278\,
            I => \button_debounce_counterZ0Z_23\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__35275\,
            I => \button_debounce_counterZ0Z_23\
        );

    \I__6727\ : CEMux
    port map (
            O => \N__35270\,
            I => \N__35267\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__35267\,
            I => \N__35264\
        );

    \I__6725\ : Span4Mux_h
    port map (
            O => \N__35264\,
            I => \N__35261\
        );

    \I__6724\ : Span4Mux_v
    port map (
            O => \N__35261\,
            I => \N__35258\
        );

    \I__6723\ : Odrv4
    port map (
            O => \N__35258\,
            I => \LED3_c_0\
        );

    \I__6722\ : InMux
    port map (
            O => \N__35255\,
            I => \N__35252\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__35252\,
            I => \N__35249\
        );

    \I__6720\ : Span4Mux_h
    port map (
            O => \N__35249\,
            I => \N__35245\
        );

    \I__6719\ : InMux
    port map (
            O => \N__35248\,
            I => \N__35242\
        );

    \I__6718\ : Odrv4
    port map (
            O => \N__35245\,
            I => \sRAM_pointer_readZ0Z_5\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__35242\,
            I => \sRAM_pointer_readZ0Z_5\
        );

    \I__6716\ : InMux
    port map (
            O => \N__35237\,
            I => \N__35234\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__35234\,
            I => \N__35231\
        );

    \I__6714\ : Span12Mux_v
    port map (
            O => \N__35231\,
            I => \N__35228\
        );

    \I__6713\ : Span12Mux_h
    port map (
            O => \N__35228\,
            I => \N__35224\
        );

    \I__6712\ : InMux
    port map (
            O => \N__35227\,
            I => \N__35221\
        );

    \I__6711\ : Odrv12
    port map (
            O => \N__35224\,
            I => \sRAM_pointer_writeZ0Z_5\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__35221\,
            I => \sRAM_pointer_writeZ0Z_5\
        );

    \I__6709\ : IoInMux
    port map (
            O => \N__35216\,
            I => \N__35213\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__35213\,
            I => \N__35210\
        );

    \I__6707\ : Span4Mux_s3_h
    port map (
            O => \N__35210\,
            I => \N__35207\
        );

    \I__6706\ : Span4Mux_h
    port map (
            O => \N__35207\,
            I => \N__35204\
        );

    \I__6705\ : Span4Mux_h
    port map (
            O => \N__35204\,
            I => \N__35201\
        );

    \I__6704\ : Span4Mux_v
    port map (
            O => \N__35201\,
            I => \N__35198\
        );

    \I__6703\ : Odrv4
    port map (
            O => \N__35198\,
            I => \RAM_ADD_c_5\
        );

    \I__6702\ : InMux
    port map (
            O => \N__35195\,
            I => un1_button_debounce_counter_cry_9
        );

    \I__6701\ : InMux
    port map (
            O => \N__35192\,
            I => un1_button_debounce_counter_cry_10
        );

    \I__6700\ : InMux
    port map (
            O => \N__35189\,
            I => un1_button_debounce_counter_cry_11
        );

    \I__6699\ : InMux
    port map (
            O => \N__35186\,
            I => un1_button_debounce_counter_cry_12
        );

    \I__6698\ : InMux
    port map (
            O => \N__35183\,
            I => un1_button_debounce_counter_cry_13
        );

    \I__6697\ : InMux
    port map (
            O => \N__35180\,
            I => \N__35176\
        );

    \I__6696\ : InMux
    port map (
            O => \N__35179\,
            I => \N__35173\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__35176\,
            I => \N__35170\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__35173\,
            I => \button_debounce_counterZ0Z_15\
        );

    \I__6693\ : Odrv4
    port map (
            O => \N__35170\,
            I => \button_debounce_counterZ0Z_15\
        );

    \I__6692\ : InMux
    port map (
            O => \N__35165\,
            I => un1_button_debounce_counter_cry_14
        );

    \I__6691\ : InMux
    port map (
            O => \N__35162\,
            I => \N__35159\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__35159\,
            I => \N__35155\
        );

    \I__6689\ : InMux
    port map (
            O => \N__35158\,
            I => \N__35152\
        );

    \I__6688\ : Span4Mux_h
    port map (
            O => \N__35155\,
            I => \N__35149\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__35152\,
            I => \button_debounce_counterZ0Z_16\
        );

    \I__6686\ : Odrv4
    port map (
            O => \N__35149\,
            I => \button_debounce_counterZ0Z_16\
        );

    \I__6685\ : InMux
    port map (
            O => \N__35144\,
            I => un1_button_debounce_counter_cry_15
        );

    \I__6684\ : InMux
    port map (
            O => \N__35141\,
            I => \N__35137\
        );

    \I__6683\ : InMux
    port map (
            O => \N__35140\,
            I => \N__35134\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__35137\,
            I => \N__35131\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__35134\,
            I => \button_debounce_counterZ0Z_17\
        );

    \I__6680\ : Odrv4
    port map (
            O => \N__35131\,
            I => \button_debounce_counterZ0Z_17\
        );

    \I__6679\ : InMux
    port map (
            O => \N__35126\,
            I => \bfn_16_15_0_\
        );

    \I__6678\ : InMux
    port map (
            O => \N__35123\,
            I => \N__35119\
        );

    \I__6677\ : InMux
    port map (
            O => \N__35122\,
            I => \N__35116\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__35119\,
            I => \button_debounce_counterZ0Z_18\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__35116\,
            I => \button_debounce_counterZ0Z_18\
        );

    \I__6674\ : InMux
    port map (
            O => \N__35111\,
            I => un1_button_debounce_counter_cry_17
        );

    \I__6673\ : CascadeMux
    port map (
            O => \N__35108\,
            I => \N__35105\
        );

    \I__6672\ : InMux
    port map (
            O => \N__35105\,
            I => \N__35102\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__35102\,
            I => \N__35098\
        );

    \I__6670\ : InMux
    port map (
            O => \N__35101\,
            I => \N__35095\
        );

    \I__6669\ : Odrv12
    port map (
            O => \N__35098\,
            I => \button_debounce_counterZ0Z_2\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__35095\,
            I => \button_debounce_counterZ0Z_2\
        );

    \I__6667\ : InMux
    port map (
            O => \N__35090\,
            I => un1_button_debounce_counter_cry_1
        );

    \I__6666\ : InMux
    port map (
            O => \N__35087\,
            I => \N__35083\
        );

    \I__6665\ : InMux
    port map (
            O => \N__35086\,
            I => \N__35080\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__35083\,
            I => \button_debounce_counterZ0Z_3\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__35080\,
            I => \button_debounce_counterZ0Z_3\
        );

    \I__6662\ : InMux
    port map (
            O => \N__35075\,
            I => un1_button_debounce_counter_cry_2
        );

    \I__6661\ : InMux
    port map (
            O => \N__35072\,
            I => \N__35068\
        );

    \I__6660\ : InMux
    port map (
            O => \N__35071\,
            I => \N__35065\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__35068\,
            I => \button_debounce_counterZ0Z_4\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__35065\,
            I => \button_debounce_counterZ0Z_4\
        );

    \I__6657\ : InMux
    port map (
            O => \N__35060\,
            I => un1_button_debounce_counter_cry_3
        );

    \I__6656\ : CascadeMux
    port map (
            O => \N__35057\,
            I => \N__35054\
        );

    \I__6655\ : InMux
    port map (
            O => \N__35054\,
            I => \N__35050\
        );

    \I__6654\ : InMux
    port map (
            O => \N__35053\,
            I => \N__35047\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__35050\,
            I => \button_debounce_counterZ0Z_5\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__35047\,
            I => \button_debounce_counterZ0Z_5\
        );

    \I__6651\ : InMux
    port map (
            O => \N__35042\,
            I => un1_button_debounce_counter_cry_4
        );

    \I__6650\ : InMux
    port map (
            O => \N__35039\,
            I => \N__35036\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__35036\,
            I => \N__35032\
        );

    \I__6648\ : InMux
    port map (
            O => \N__35035\,
            I => \N__35029\
        );

    \I__6647\ : Odrv4
    port map (
            O => \N__35032\,
            I => \button_debounce_counterZ0Z_6\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__35029\,
            I => \button_debounce_counterZ0Z_6\
        );

    \I__6645\ : InMux
    port map (
            O => \N__35024\,
            I => un1_button_debounce_counter_cry_5
        );

    \I__6644\ : InMux
    port map (
            O => \N__35021\,
            I => un1_button_debounce_counter_cry_6
        );

    \I__6643\ : InMux
    port map (
            O => \N__35018\,
            I => un1_button_debounce_counter_cry_7
        );

    \I__6642\ : InMux
    port map (
            O => \N__35015\,
            I => \bfn_16_14_0_\
        );

    \I__6641\ : InMux
    port map (
            O => \N__35012\,
            I => \N__35009\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__35009\,
            I => \N__35006\
        );

    \I__6639\ : Span4Mux_h
    port map (
            O => \N__35006\,
            I => \N__35003\
        );

    \I__6638\ : Span4Mux_v
    port map (
            O => \N__35003\,
            I => \N__35000\
        );

    \I__6637\ : Odrv4
    port map (
            O => \N__35000\,
            I => \sDAC_mem_19Z0Z_3\
        );

    \I__6636\ : CEMux
    port map (
            O => \N__34997\,
            I => \N__34994\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__34994\,
            I => \N__34991\
        );

    \I__6634\ : Span4Mux_v
    port map (
            O => \N__34991\,
            I => \N__34987\
        );

    \I__6633\ : CEMux
    port map (
            O => \N__34990\,
            I => \N__34984\
        );

    \I__6632\ : Span4Mux_v
    port map (
            O => \N__34987\,
            I => \N__34979\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__34984\,
            I => \N__34979\
        );

    \I__6630\ : Odrv4
    port map (
            O => \N__34979\,
            I => \sDAC_mem_19_1_sqmuxa\
        );

    \I__6629\ : InMux
    port map (
            O => \N__34976\,
            I => \N__34973\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__34973\,
            I => \N__34970\
        );

    \I__6627\ : Span12Mux_v
    port map (
            O => \N__34970\,
            I => \N__34967\
        );

    \I__6626\ : Odrv12
    port map (
            O => \N__34967\,
            I => \sDAC_mem_35Z0Z_7\
        );

    \I__6625\ : InMux
    port map (
            O => \N__34964\,
            I => \N__34961\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__34961\,
            I => \sDAC_data_2_6_bm_1_10\
        );

    \I__6623\ : CascadeMux
    port map (
            O => \N__34958\,
            I => \sDAC_data_RNO_15Z0Z_10_cascade_\
        );

    \I__6622\ : InMux
    port map (
            O => \N__34955\,
            I => \N__34952\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__34952\,
            I => \N__34949\
        );

    \I__6620\ : Odrv4
    port map (
            O => \N__34949\,
            I => \sDAC_data_RNO_5Z0Z_10\
        );

    \I__6619\ : CascadeMux
    port map (
            O => \N__34946\,
            I => \sDAC_data_2_14_ns_1_10_cascade_\
        );

    \I__6618\ : InMux
    port map (
            O => \N__34943\,
            I => \N__34940\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__34940\,
            I => \sDAC_data_RNO_1Z0Z_10\
        );

    \I__6616\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34934\
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__34934\,
            I => \N__34931\
        );

    \I__6614\ : Span4Mux_h
    port map (
            O => \N__34931\,
            I => \N__34928\
        );

    \I__6613\ : Span4Mux_v
    port map (
            O => \N__34928\,
            I => \N__34925\
        );

    \I__6612\ : Span4Mux_v
    port map (
            O => \N__34925\,
            I => \N__34922\
        );

    \I__6611\ : Odrv4
    port map (
            O => \N__34922\,
            I => \sDAC_mem_36Z0Z_7\
        );

    \I__6610\ : CascadeMux
    port map (
            O => \N__34919\,
            I => \sDAC_data_2_13_am_1_10_cascade_\
        );

    \I__6609\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34913\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__34913\,
            I => \sDAC_data_RNO_4Z0Z_10\
        );

    \I__6607\ : InMux
    port map (
            O => \N__34910\,
            I => \N__34907\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__34907\,
            I => \sDAC_data_RNO_26Z0Z_10\
        );

    \I__6605\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34901\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__34901\,
            I => \sDAC_data_RNO_14Z0Z_10\
        );

    \I__6603\ : CascadeMux
    port map (
            O => \N__34898\,
            I => \sDAC_data_2_20_am_1_3_cascade_\
        );

    \I__6602\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34892\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__34892\,
            I => \N__34889\
        );

    \I__6600\ : Span4Mux_h
    port map (
            O => \N__34889\,
            I => \N__34886\
        );

    \I__6599\ : Odrv4
    port map (
            O => \N__34886\,
            I => \sDAC_data_2_24_ns_1_3\
        );

    \I__6598\ : CascadeMux
    port map (
            O => \N__34883\,
            I => \sDAC_data_RNO_7Z0Z_3_cascade_\
        );

    \I__6597\ : InMux
    port map (
            O => \N__34880\,
            I => \N__34877\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__34877\,
            I => \sDAC_data_RNO_8Z0Z_3\
        );

    \I__6595\ : InMux
    port map (
            O => \N__34874\,
            I => \N__34871\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__34871\,
            I => \N__34868\
        );

    \I__6593\ : Span4Mux_v
    port map (
            O => \N__34868\,
            I => \N__34863\
        );

    \I__6592\ : InMux
    port map (
            O => \N__34867\,
            I => \N__34860\
        );

    \I__6591\ : CascadeMux
    port map (
            O => \N__34866\,
            I => \N__34854\
        );

    \I__6590\ : Span4Mux_h
    port map (
            O => \N__34863\,
            I => \N__34850\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__34860\,
            I => \N__34847\
        );

    \I__6588\ : InMux
    port map (
            O => \N__34859\,
            I => \N__34836\
        );

    \I__6587\ : InMux
    port map (
            O => \N__34858\,
            I => \N__34836\
        );

    \I__6586\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34836\
        );

    \I__6585\ : InMux
    port map (
            O => \N__34854\,
            I => \N__34836\
        );

    \I__6584\ : InMux
    port map (
            O => \N__34853\,
            I => \N__34836\
        );

    \I__6583\ : Odrv4
    port map (
            O => \N__34850\,
            I => \N_333\
        );

    \I__6582\ : Odrv12
    port map (
            O => \N__34847\,
            I => \N_333\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__34836\,
            I => \N_333\
        );

    \I__6580\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34826\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__34826\,
            I => \sDAC_mem_19Z0Z_0\
        );

    \I__6578\ : InMux
    port map (
            O => \N__34823\,
            I => \N__34820\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__34820\,
            I => \N__34817\
        );

    \I__6576\ : Span4Mux_h
    port map (
            O => \N__34817\,
            I => \N__34814\
        );

    \I__6575\ : Span4Mux_h
    port map (
            O => \N__34814\,
            I => \N__34811\
        );

    \I__6574\ : Odrv4
    port map (
            O => \N__34811\,
            I => \sDAC_mem_18Z0Z_0\
        );

    \I__6573\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34805\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__34805\,
            I => \sDAC_mem_19Z0Z_1\
        );

    \I__6571\ : InMux
    port map (
            O => \N__34802\,
            I => \N__34799\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__34799\,
            I => \N__34796\
        );

    \I__6569\ : Span4Mux_h
    port map (
            O => \N__34796\,
            I => \N__34793\
        );

    \I__6568\ : Span4Mux_h
    port map (
            O => \N__34793\,
            I => \N__34790\
        );

    \I__6567\ : Odrv4
    port map (
            O => \N__34790\,
            I => \sDAC_mem_18Z0Z_1\
        );

    \I__6566\ : InMux
    port map (
            O => \N__34787\,
            I => \N__34784\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__34784\,
            I => \N__34781\
        );

    \I__6564\ : Span4Mux_v
    port map (
            O => \N__34781\,
            I => \N__34778\
        );

    \I__6563\ : Odrv4
    port map (
            O => \N__34778\,
            I => \sDAC_data_RNO_29Z0Z_4\
        );

    \I__6562\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34772\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__34772\,
            I => \sDAC_mem_19Z0Z_2\
        );

    \I__6560\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34766\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__34766\,
            I => \N__34763\
        );

    \I__6558\ : Span12Mux_v
    port map (
            O => \N__34763\,
            I => \N__34760\
        );

    \I__6557\ : Odrv12
    port map (
            O => \N__34760\,
            I => \sDAC_mem_18Z0Z_2\
        );

    \I__6556\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34754\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__34754\,
            I => \N__34751\
        );

    \I__6554\ : Span4Mux_v
    port map (
            O => \N__34751\,
            I => \N__34748\
        );

    \I__6553\ : Span4Mux_v
    port map (
            O => \N__34748\,
            I => \N__34745\
        );

    \I__6552\ : Odrv4
    port map (
            O => \N__34745\,
            I => \sDAC_mem_40Z0Z_2\
        );

    \I__6551\ : InMux
    port map (
            O => \N__34742\,
            I => \N__34739\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__34739\,
            I => \N__34736\
        );

    \I__6549\ : Span4Mux_v
    port map (
            O => \N__34736\,
            I => \N__34733\
        );

    \I__6548\ : Span4Mux_h
    port map (
            O => \N__34733\,
            I => \N__34730\
        );

    \I__6547\ : Odrv4
    port map (
            O => \N__34730\,
            I => \sDAC_mem_8Z0Z_2\
        );

    \I__6546\ : CascadeMux
    port map (
            O => \N__34727\,
            I => \sDAC_data_2_20_am_1_5_cascade_\
        );

    \I__6545\ : InMux
    port map (
            O => \N__34724\,
            I => \N__34721\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__34721\,
            I => \N__34718\
        );

    \I__6543\ : Odrv4
    port map (
            O => \N__34718\,
            I => \sDAC_data_2_24_ns_1_5\
        );

    \I__6542\ : CascadeMux
    port map (
            O => \N__34715\,
            I => \sDAC_data_RNO_7Z0Z_5_cascade_\
        );

    \I__6541\ : InMux
    port map (
            O => \N__34712\,
            I => \N__34709\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__34709\,
            I => \sDAC_data_RNO_8Z0Z_5\
        );

    \I__6539\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34703\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__34703\,
            I => \N__34700\
        );

    \I__6537\ : Span4Mux_h
    port map (
            O => \N__34700\,
            I => \N__34697\
        );

    \I__6536\ : Odrv4
    port map (
            O => \N__34697\,
            I => \sDAC_mem_34Z0Z_0\
        );

    \I__6535\ : InMux
    port map (
            O => \N__34694\,
            I => \N__34691\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__34691\,
            I => \N__34688\
        );

    \I__6533\ : Span4Mux_v
    port map (
            O => \N__34688\,
            I => \N__34685\
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__34685\,
            I => \sDAC_mem_2Z0Z_0\
        );

    \I__6531\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34679\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__34679\,
            I => \N__34676\
        );

    \I__6529\ : Span4Mux_h
    port map (
            O => \N__34676\,
            I => \N__34673\
        );

    \I__6528\ : Span4Mux_v
    port map (
            O => \N__34673\,
            I => \N__34670\
        );

    \I__6527\ : Span4Mux_h
    port map (
            O => \N__34670\,
            I => \N__34667\
        );

    \I__6526\ : Odrv4
    port map (
            O => \N__34667\,
            I => \sDAC_mem_35Z0Z_0\
        );

    \I__6525\ : CascadeMux
    port map (
            O => \N__34664\,
            I => \sDAC_data_2_6_bm_1_3_cascade_\
        );

    \I__6524\ : InMux
    port map (
            O => \N__34661\,
            I => \N__34658\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__34658\,
            I => \sDAC_mem_3Z0Z_0\
        );

    \I__6522\ : InMux
    port map (
            O => \N__34655\,
            I => \N__34652\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__34652\,
            I => \N__34649\
        );

    \I__6520\ : Span4Mux_h
    port map (
            O => \N__34649\,
            I => \N__34646\
        );

    \I__6519\ : Span4Mux_h
    port map (
            O => \N__34646\,
            I => \N__34643\
        );

    \I__6518\ : Span4Mux_v
    port map (
            O => \N__34643\,
            I => \N__34640\
        );

    \I__6517\ : Odrv4
    port map (
            O => \N__34640\,
            I => \sDAC_mem_42Z0Z_0\
        );

    \I__6516\ : InMux
    port map (
            O => \N__34637\,
            I => \N__34634\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__34634\,
            I => \N__34631\
        );

    \I__6514\ : Sp12to4
    port map (
            O => \N__34631\,
            I => \N__34628\
        );

    \I__6513\ : Span12Mux_v
    port map (
            O => \N__34628\,
            I => \N__34625\
        );

    \I__6512\ : Odrv12
    port map (
            O => \N__34625\,
            I => \sDAC_mem_10Z0Z_0\
        );

    \I__6511\ : CascadeMux
    port map (
            O => \N__34622\,
            I => \sDAC_data_RNO_17Z0Z_3_cascade_\
        );

    \I__6510\ : InMux
    port map (
            O => \N__34619\,
            I => \N__34616\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__34616\,
            I => \N__34613\
        );

    \I__6508\ : Span12Mux_v
    port map (
            O => \N__34613\,
            I => \N__34610\
        );

    \I__6507\ : Odrv12
    port map (
            O => \N__34610\,
            I => \sDAC_mem_11Z0Z_0\
        );

    \I__6506\ : InMux
    port map (
            O => \N__34607\,
            I => \N__34604\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__34604\,
            I => \N__34601\
        );

    \I__6504\ : Span4Mux_v
    port map (
            O => \N__34601\,
            I => \N__34598\
        );

    \I__6503\ : Span4Mux_v
    port map (
            O => \N__34598\,
            I => \N__34595\
        );

    \I__6502\ : Odrv4
    port map (
            O => \N__34595\,
            I => \sDAC_mem_40Z0Z_0\
        );

    \I__6501\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34589\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__34589\,
            I => \N__34586\
        );

    \I__6499\ : Span4Mux_v
    port map (
            O => \N__34586\,
            I => \N__34583\
        );

    \I__6498\ : Span4Mux_h
    port map (
            O => \N__34583\,
            I => \N__34580\
        );

    \I__6497\ : Odrv4
    port map (
            O => \N__34580\,
            I => \sDAC_mem_8Z0Z_0\
        );

    \I__6496\ : InMux
    port map (
            O => \N__34577\,
            I => \sDAC_mem_pointer_0_cry_1\
        );

    \I__6495\ : InMux
    port map (
            O => \N__34574\,
            I => \sDAC_mem_pointer_0_cry_2\
        );

    \I__6494\ : InMux
    port map (
            O => \N__34571\,
            I => \sDAC_mem_pointer_0_cry_3\
        );

    \I__6493\ : InMux
    port map (
            O => \N__34568\,
            I => \sDAC_mem_pointer_0_cry_4\
        );

    \I__6492\ : InMux
    port map (
            O => \N__34565\,
            I => \N__34562\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__34562\,
            I => \N__34559\
        );

    \I__6490\ : Span4Mux_h
    port map (
            O => \N__34559\,
            I => \N__34556\
        );

    \I__6489\ : Odrv4
    port map (
            O => \N__34556\,
            I => \sDAC_mem_34Z0Z_2\
        );

    \I__6488\ : InMux
    port map (
            O => \N__34553\,
            I => \N__34550\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__34550\,
            I => \N__34547\
        );

    \I__6486\ : Span4Mux_h
    port map (
            O => \N__34547\,
            I => \N__34544\
        );

    \I__6485\ : Odrv4
    port map (
            O => \N__34544\,
            I => \sDAC_mem_2Z0Z_2\
        );

    \I__6484\ : InMux
    port map (
            O => \N__34541\,
            I => \N__34538\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__34538\,
            I => \N__34535\
        );

    \I__6482\ : Span4Mux_h
    port map (
            O => \N__34535\,
            I => \N__34532\
        );

    \I__6481\ : Span4Mux_h
    port map (
            O => \N__34532\,
            I => \N__34529\
        );

    \I__6480\ : Span4Mux_h
    port map (
            O => \N__34529\,
            I => \N__34526\
        );

    \I__6479\ : Odrv4
    port map (
            O => \N__34526\,
            I => \sDAC_mem_35Z0Z_2\
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__34523\,
            I => \sDAC_data_2_6_bm_1_5_cascade_\
        );

    \I__6477\ : InMux
    port map (
            O => \N__34520\,
            I => \N__34517\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__34517\,
            I => \sDAC_mem_3Z0Z_2\
        );

    \I__6475\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34511\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__34511\,
            I => \N__34508\
        );

    \I__6473\ : Span12Mux_v
    port map (
            O => \N__34508\,
            I => \N__34505\
        );

    \I__6472\ : Odrv12
    port map (
            O => \N__34505\,
            I => \sDAC_mem_42Z0Z_2\
        );

    \I__6471\ : InMux
    port map (
            O => \N__34502\,
            I => \N__34499\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__34499\,
            I => \N__34496\
        );

    \I__6469\ : Span4Mux_v
    port map (
            O => \N__34496\,
            I => \N__34493\
        );

    \I__6468\ : Span4Mux_h
    port map (
            O => \N__34493\,
            I => \N__34490\
        );

    \I__6467\ : Odrv4
    port map (
            O => \N__34490\,
            I => \sDAC_mem_10Z0Z_2\
        );

    \I__6466\ : CascadeMux
    port map (
            O => \N__34487\,
            I => \sDAC_data_RNO_17Z0Z_5_cascade_\
        );

    \I__6465\ : InMux
    port map (
            O => \N__34484\,
            I => \N__34481\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__34481\,
            I => \N__34478\
        );

    \I__6463\ : Span4Mux_h
    port map (
            O => \N__34478\,
            I => \N__34475\
        );

    \I__6462\ : Span4Mux_h
    port map (
            O => \N__34475\,
            I => \N__34472\
        );

    \I__6461\ : Odrv4
    port map (
            O => \N__34472\,
            I => \sDAC_mem_11Z0Z_2\
        );

    \I__6460\ : CascadeMux
    port map (
            O => \N__34469\,
            I => \sDAC_data_RNO_26Z0Z_9_cascade_\
        );

    \I__6459\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34463\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__34463\,
            I => \sDAC_mem_32Z0Z_6\
        );

    \I__6457\ : InMux
    port map (
            O => \N__34460\,
            I => \N__34457\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__34457\,
            I => \sDAC_data_RNO_14Z0Z_9\
        );

    \I__6455\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34451\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__34451\,
            I => \N__34448\
        );

    \I__6453\ : Odrv12
    port map (
            O => \N__34448\,
            I => \sDAC_mem_21Z0Z_0\
        );

    \I__6452\ : InMux
    port map (
            O => \N__34445\,
            I => \N__34442\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__34442\,
            I => \N__34439\
        );

    \I__6450\ : Odrv12
    port map (
            O => \N__34439\,
            I => \sDAC_mem_21Z0Z_1\
        );

    \I__6449\ : InMux
    port map (
            O => \N__34436\,
            I => \N__34433\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__34433\,
            I => \N__34430\
        );

    \I__6447\ : Span4Mux_v
    port map (
            O => \N__34430\,
            I => \N__34427\
        );

    \I__6446\ : Odrv4
    port map (
            O => \N__34427\,
            I => \sDAC_data_RNO_20Z0Z_4\
        );

    \I__6445\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34421\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__34421\,
            I => \N__34418\
        );

    \I__6443\ : Odrv4
    port map (
            O => \N__34418\,
            I => \sDAC_mem_21Z0Z_2\
        );

    \I__6442\ : InMux
    port map (
            O => \N__34415\,
            I => \N__34412\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__34412\,
            I => \N__34409\
        );

    \I__6440\ : Odrv4
    port map (
            O => \N__34409\,
            I => \sDAC_mem_21Z0Z_3\
        );

    \I__6439\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34403\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__34403\,
            I => \N__34400\
        );

    \I__6437\ : Span4Mux_h
    port map (
            O => \N__34400\,
            I => \N__34397\
        );

    \I__6436\ : Odrv4
    port map (
            O => \N__34397\,
            I => \sDAC_data_RNO_20Z0Z_6\
        );

    \I__6435\ : InMux
    port map (
            O => \N__34394\,
            I => \N__34391\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__34391\,
            I => \N__34388\
        );

    \I__6433\ : Odrv4
    port map (
            O => \N__34388\,
            I => \sDAC_mem_21Z0Z_4\
        );

    \I__6432\ : InMux
    port map (
            O => \N__34385\,
            I => \N__34382\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__34382\,
            I => \N__34379\
        );

    \I__6430\ : Odrv4
    port map (
            O => \N__34379\,
            I => \sDAC_data_RNO_20Z0Z_7\
        );

    \I__6429\ : InMux
    port map (
            O => \N__34376\,
            I => \N__34373\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__34373\,
            I => \N__34370\
        );

    \I__6427\ : Span4Mux_h
    port map (
            O => \N__34370\,
            I => \N__34367\
        );

    \I__6426\ : Odrv4
    port map (
            O => \N__34367\,
            I => \sDAC_mem_34Z0Z_6\
        );

    \I__6425\ : InMux
    port map (
            O => \N__34364\,
            I => \N__34361\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__34361\,
            I => \N__34358\
        );

    \I__6423\ : Odrv12
    port map (
            O => \N__34358\,
            I => \sDAC_mem_2Z0Z_6\
        );

    \I__6422\ : InMux
    port map (
            O => \N__34355\,
            I => \N__34352\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__34352\,
            I => \N__34349\
        );

    \I__6420\ : Odrv12
    port map (
            O => \N__34349\,
            I => \sDAC_mem_35Z0Z_6\
        );

    \I__6419\ : CascadeMux
    port map (
            O => \N__34346\,
            I => \sDAC_data_2_6_bm_1_9_cascade_\
        );

    \I__6418\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34340\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__34340\,
            I => \sDAC_mem_3Z0Z_6\
        );

    \I__6416\ : InMux
    port map (
            O => \N__34337\,
            I => \N__34334\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__34334\,
            I => \sDAC_data_RNO_15Z0Z_9\
        );

    \I__6414\ : InMux
    port map (
            O => \N__34331\,
            I => \N__34328\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__34328\,
            I => \N__34325\
        );

    \I__6412\ : Span4Mux_h
    port map (
            O => \N__34325\,
            I => \N__34322\
        );

    \I__6411\ : Span4Mux_h
    port map (
            O => \N__34322\,
            I => \N__34319\
        );

    \I__6410\ : Odrv4
    port map (
            O => \N__34319\,
            I => \sDAC_mem_42Z0Z_6\
        );

    \I__6409\ : InMux
    port map (
            O => \N__34316\,
            I => \N__34313\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__34313\,
            I => \N__34310\
        );

    \I__6407\ : Span4Mux_h
    port map (
            O => \N__34310\,
            I => \N__34307\
        );

    \I__6406\ : Span4Mux_h
    port map (
            O => \N__34307\,
            I => \N__34304\
        );

    \I__6405\ : Odrv4
    port map (
            O => \N__34304\,
            I => \sDAC_mem_10Z0Z_6\
        );

    \I__6404\ : CascadeMux
    port map (
            O => \N__34301\,
            I => \sDAC_data_RNO_17Z0Z_9_cascade_\
        );

    \I__6403\ : InMux
    port map (
            O => \N__34298\,
            I => \N__34295\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__34295\,
            I => \N__34292\
        );

    \I__6401\ : Odrv12
    port map (
            O => \N__34292\,
            I => \sDAC_mem_11Z0Z_6\
        );

    \I__6400\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34286\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__34286\,
            I => \N__34283\
        );

    \I__6398\ : Span4Mux_h
    port map (
            O => \N__34283\,
            I => \N__34280\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__34280\,
            I => \sDAC_mem_40Z0Z_6\
        );

    \I__6396\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34274\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__34274\,
            I => \N__34271\
        );

    \I__6394\ : Span4Mux_h
    port map (
            O => \N__34271\,
            I => \N__34268\
        );

    \I__6393\ : Odrv4
    port map (
            O => \N__34268\,
            I => \sDAC_mem_8Z0Z_6\
        );

    \I__6392\ : CascadeMux
    port map (
            O => \N__34265\,
            I => \sDAC_data_2_20_am_1_9_cascade_\
        );

    \I__6391\ : CascadeMux
    port map (
            O => \N__34262\,
            I => \sDAC_data_RNO_7Z0Z_9_cascade_\
        );

    \I__6390\ : InMux
    port map (
            O => \N__34259\,
            I => \N__34256\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__34256\,
            I => \sDAC_data_RNO_8Z0Z_9\
        );

    \I__6388\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34250\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__34250\,
            I => \sDAC_data_RNO_2Z0Z_9\
        );

    \I__6386\ : CEMux
    port map (
            O => \N__34247\,
            I => \N__34244\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__34244\,
            I => \N__34241\
        );

    \I__6384\ : Span4Mux_h
    port map (
            O => \N__34241\,
            I => \N__34238\
        );

    \I__6383\ : Odrv4
    port map (
            O => \N__34238\,
            I => \sDAC_mem_21_1_sqmuxa\
        );

    \I__6382\ : InMux
    port map (
            O => \N__34235\,
            I => \N__34232\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__34232\,
            I => \N__34229\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__34229\,
            I => \N__34226\
        );

    \I__6379\ : Odrv4
    port map (
            O => \N__34226\,
            I => \sDAC_mem_34Z0Z_4\
        );

    \I__6378\ : InMux
    port map (
            O => \N__34223\,
            I => \N__34220\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__34220\,
            I => \N__34217\
        );

    \I__6376\ : Span4Mux_h
    port map (
            O => \N__34217\,
            I => \N__34214\
        );

    \I__6375\ : Odrv4
    port map (
            O => \N__34214\,
            I => \sDAC_mem_2Z0Z_4\
        );

    \I__6374\ : InMux
    port map (
            O => \N__34211\,
            I => \N__34208\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__34208\,
            I => \N__34205\
        );

    \I__6372\ : Span4Mux_v
    port map (
            O => \N__34205\,
            I => \N__34202\
        );

    \I__6371\ : Sp12to4
    port map (
            O => \N__34202\,
            I => \N__34199\
        );

    \I__6370\ : Odrv12
    port map (
            O => \N__34199\,
            I => \sDAC_mem_35Z0Z_4\
        );

    \I__6369\ : CascadeMux
    port map (
            O => \N__34196\,
            I => \sDAC_data_2_6_bm_1_7_cascade_\
        );

    \I__6368\ : InMux
    port map (
            O => \N__34193\,
            I => \N__34190\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__34190\,
            I => \sDAC_mem_3Z0Z_4\
        );

    \I__6366\ : InMux
    port map (
            O => \N__34187\,
            I => \N__34184\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__34184\,
            I => \sDAC_data_RNO_15Z0Z_7\
        );

    \I__6364\ : InMux
    port map (
            O => \N__34181\,
            I => \N__34178\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__34178\,
            I => \N__34175\
        );

    \I__6362\ : Span4Mux_h
    port map (
            O => \N__34175\,
            I => \N__34172\
        );

    \I__6361\ : Odrv4
    port map (
            O => \N__34172\,
            I => \sDAC_mem_40Z0Z_4\
        );

    \I__6360\ : InMux
    port map (
            O => \N__34169\,
            I => \N__34166\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__34166\,
            I => \N__34163\
        );

    \I__6358\ : Span12Mux_v
    port map (
            O => \N__34163\,
            I => \N__34160\
        );

    \I__6357\ : Odrv12
    port map (
            O => \N__34160\,
            I => \sDAC_mem_8Z0Z_4\
        );

    \I__6356\ : CascadeMux
    port map (
            O => \N__34157\,
            I => \sDAC_data_2_20_am_1_7_cascade_\
        );

    \I__6355\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34151\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__34151\,
            I => \N__34148\
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__34148\,
            I => \sDAC_data_2_24_ns_1_7\
        );

    \I__6352\ : CascadeMux
    port map (
            O => \N__34145\,
            I => \sDAC_data_RNO_7Z0Z_7_cascade_\
        );

    \I__6351\ : InMux
    port map (
            O => \N__34142\,
            I => \N__34139\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__34139\,
            I => \sDAC_data_RNO_2Z0Z_7\
        );

    \I__6349\ : InMux
    port map (
            O => \N__34136\,
            I => \N__34133\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__34133\,
            I => \N__34130\
        );

    \I__6347\ : Span4Mux_h
    port map (
            O => \N__34130\,
            I => \N__34127\
        );

    \I__6346\ : Span4Mux_h
    port map (
            O => \N__34127\,
            I => \N__34124\
        );

    \I__6345\ : Odrv4
    port map (
            O => \N__34124\,
            I => \sDAC_mem_11Z0Z_4\
        );

    \I__6344\ : InMux
    port map (
            O => \N__34121\,
            I => \N__34118\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__34118\,
            I => \sDAC_data_RNO_8Z0Z_7\
        );

    \I__6342\ : InMux
    port map (
            O => \N__34115\,
            I => \N__34112\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__34112\,
            I => \N__34109\
        );

    \I__6340\ : Odrv12
    port map (
            O => \N__34109\,
            I => \sDAC_mem_42Z0Z_4\
        );

    \I__6339\ : InMux
    port map (
            O => \N__34106\,
            I => \N__34103\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__34103\,
            I => \N__34100\
        );

    \I__6337\ : Odrv12
    port map (
            O => \N__34100\,
            I => \sDAC_mem_10Z0Z_4\
        );

    \I__6336\ : InMux
    port map (
            O => \N__34097\,
            I => \N__34094\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__34094\,
            I => \sDAC_data_RNO_17Z0Z_7\
        );

    \I__6334\ : InMux
    port map (
            O => \N__34091\,
            I => \N__34088\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__34088\,
            I => \N__34085\
        );

    \I__6332\ : Span4Mux_h
    port map (
            O => \N__34085\,
            I => \N__34082\
        );

    \I__6331\ : Odrv4
    port map (
            O => \N__34082\,
            I => \sDAC_mem_19Z0Z_6\
        );

    \I__6330\ : InMux
    port map (
            O => \N__34079\,
            I => \N__34076\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__34076\,
            I => \N__34073\
        );

    \I__6328\ : Sp12to4
    port map (
            O => \N__34073\,
            I => \N__34070\
        );

    \I__6327\ : Odrv12
    port map (
            O => \N__34070\,
            I => \sDAC_mem_19Z0Z_7\
        );

    \I__6326\ : InMux
    port map (
            O => \N__34067\,
            I => \N__34064\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__34064\,
            I => \N__34061\
        );

    \I__6324\ : Odrv4
    port map (
            O => \N__34061\,
            I => \sDAC_mem_21Z0Z_5\
        );

    \I__6323\ : InMux
    port map (
            O => \N__34058\,
            I => \N__34055\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__34055\,
            I => \N__34052\
        );

    \I__6321\ : Span4Mux_h
    port map (
            O => \N__34052\,
            I => \N__34049\
        );

    \I__6320\ : Odrv4
    port map (
            O => \N__34049\,
            I => \sDAC_mem_21Z0Z_6\
        );

    \I__6319\ : InMux
    port map (
            O => \N__34046\,
            I => \N__34043\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__34043\,
            I => \N__34040\
        );

    \I__6317\ : Span4Mux_v
    port map (
            O => \N__34040\,
            I => \N__34037\
        );

    \I__6316\ : Span4Mux_v
    port map (
            O => \N__34037\,
            I => \N__34034\
        );

    \I__6315\ : Odrv4
    port map (
            O => \N__34034\,
            I => \sDAC_mem_21Z0Z_7\
        );

    \I__6314\ : CascadeMux
    port map (
            O => \N__34031\,
            I => \sRead_data_RNOZ0Z_0_cascade_\
        );

    \I__6313\ : IoInMux
    port map (
            O => \N__34028\,
            I => \N__34025\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__34025\,
            I => \N__34022\
        );

    \I__6311\ : IoSpan4Mux
    port map (
            O => \N__34022\,
            I => \N__34019\
        );

    \I__6310\ : IoSpan4Mux
    port map (
            O => \N__34019\,
            I => \N__34016\
        );

    \I__6309\ : Span4Mux_s3_v
    port map (
            O => \N__34016\,
            I => \N__34010\
        );

    \I__6308\ : InMux
    port map (
            O => \N__34015\,
            I => \N__34007\
        );

    \I__6307\ : InMux
    port map (
            O => \N__34014\,
            I => \N__34001\
        );

    \I__6306\ : InMux
    port map (
            O => \N__34013\,
            I => \N__34001\
        );

    \I__6305\ : Span4Mux_v
    port map (
            O => \N__34010\,
            I => \N__33996\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__34007\,
            I => \N__33996\
        );

    \I__6303\ : InMux
    port map (
            O => \N__34006\,
            I => \N__33993\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__34001\,
            I => \N__33990\
        );

    \I__6301\ : Odrv4
    port map (
            O => \N__33996\,
            I => \ADC_clk_c\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__33993\,
            I => \ADC_clk_c\
        );

    \I__6299\ : Odrv4
    port map (
            O => \N__33990\,
            I => \ADC_clk_c\
        );

    \I__6298\ : InMux
    port map (
            O => \N__33983\,
            I => \N__33979\
        );

    \I__6297\ : InMux
    port map (
            O => \N__33982\,
            I => \N__33976\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__33979\,
            I => \sRead_dataZ0\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__33976\,
            I => \sRead_dataZ0\
        );

    \I__6294\ : InMux
    port map (
            O => \N__33971\,
            I => \N__33968\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__33968\,
            I => spi_data_miso_0_sqmuxa_2_i_o2_4
        );

    \I__6292\ : InMux
    port map (
            O => \N__33965\,
            I => \N__33962\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__33962\,
            I => spi_data_miso_0_sqmuxa_2_i_o2_5
        );

    \I__6290\ : InMux
    port map (
            O => \N__33959\,
            I => \N__33956\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__33956\,
            I => \N__33953\
        );

    \I__6288\ : Span12Mux_v
    port map (
            O => \N__33953\,
            I => \N__33950\
        );

    \I__6287\ : Span12Mux_h
    port map (
            O => \N__33950\,
            I => \N__33947\
        );

    \I__6286\ : Odrv12
    port map (
            O => \N__33947\,
            I => \ADC3_c\
        );

    \I__6285\ : IoInMux
    port map (
            O => \N__33944\,
            I => \N__33941\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__33941\,
            I => \N__33938\
        );

    \I__6283\ : Span4Mux_s2_v
    port map (
            O => \N__33938\,
            I => \N__33935\
        );

    \I__6282\ : Span4Mux_h
    port map (
            O => \N__33935\,
            I => \N__33932\
        );

    \I__6281\ : Span4Mux_h
    port map (
            O => \N__33932\,
            I => \N__33929\
        );

    \I__6280\ : Span4Mux_v
    port map (
            O => \N__33929\,
            I => \N__33926\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__33926\,
            I => \RAM_DATA_1Z0Z_3\
        );

    \I__6278\ : InMux
    port map (
            O => \N__33923\,
            I => \N__33920\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__33920\,
            I => \N__33917\
        );

    \I__6276\ : Span4Mux_h
    port map (
            O => \N__33917\,
            I => \N__33914\
        );

    \I__6275\ : Odrv4
    port map (
            O => \N__33914\,
            I => \sDAC_mem_19Z0Z_4\
        );

    \I__6274\ : InMux
    port map (
            O => \N__33911\,
            I => \N__33908\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__33908\,
            I => \N__33905\
        );

    \I__6272\ : Span4Mux_h
    port map (
            O => \N__33905\,
            I => \N__33902\
        );

    \I__6271\ : Odrv4
    port map (
            O => \N__33902\,
            I => \sDAC_mem_19Z0Z_5\
        );

    \I__6270\ : InMux
    port map (
            O => \N__33899\,
            I => \N__33896\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__33896\,
            I => \sDAC_mem_22Z0Z_6\
        );

    \I__6268\ : CEMux
    port map (
            O => \N__33893\,
            I => \N__33890\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__33890\,
            I => \N__33887\
        );

    \I__6266\ : Span4Mux_v
    port map (
            O => \N__33887\,
            I => \N__33884\
        );

    \I__6265\ : Span4Mux_v
    port map (
            O => \N__33884\,
            I => \N__33880\
        );

    \I__6264\ : CEMux
    port map (
            O => \N__33883\,
            I => \N__33877\
        );

    \I__6263\ : Span4Mux_h
    port map (
            O => \N__33880\,
            I => \N__33872\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__33877\,
            I => \N__33872\
        );

    \I__6261\ : Odrv4
    port map (
            O => \N__33872\,
            I => \sDAC_mem_22_1_sqmuxa\
        );

    \I__6260\ : InMux
    port map (
            O => \N__33869\,
            I => \N__33866\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__33866\,
            I => \N__33863\
        );

    \I__6258\ : Odrv12
    port map (
            O => \N__33863\,
            I => \sDAC_mem_29Z0Z_0\
        );

    \I__6257\ : InMux
    port map (
            O => \N__33860\,
            I => \N__33857\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__33857\,
            I => \N__33854\
        );

    \I__6255\ : Span4Mux_v
    port map (
            O => \N__33854\,
            I => \N__33851\
        );

    \I__6254\ : Span4Mux_h
    port map (
            O => \N__33851\,
            I => \N__33848\
        );

    \I__6253\ : Odrv4
    port map (
            O => \N__33848\,
            I => \sDAC_mem_28Z0Z_0\
        );

    \I__6252\ : InMux
    port map (
            O => \N__33845\,
            I => \N__33842\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__33842\,
            I => \sDAC_data_RNO_23Z0Z_3\
        );

    \I__6250\ : InMux
    port map (
            O => \N__33839\,
            I => \N__33836\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__33836\,
            I => \N__33833\
        );

    \I__6248\ : Span4Mux_h
    port map (
            O => \N__33833\,
            I => \N__33830\
        );

    \I__6247\ : Odrv4
    port map (
            O => \N__33830\,
            I => \sDAC_mem_29Z0Z_3\
        );

    \I__6246\ : InMux
    port map (
            O => \N__33827\,
            I => \N__33824\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__33824\,
            I => \N__33821\
        );

    \I__6244\ : Span4Mux_h
    port map (
            O => \N__33821\,
            I => \N__33818\
        );

    \I__6243\ : Span4Mux_h
    port map (
            O => \N__33818\,
            I => \N__33815\
        );

    \I__6242\ : Odrv4
    port map (
            O => \N__33815\,
            I => \sDAC_mem_28Z0Z_3\
        );

    \I__6241\ : CascadeMux
    port map (
            O => \N__33812\,
            I => \sbuttonModeStatus_0_sqmuxa_14_cascade_\
        );

    \I__6240\ : InMux
    port map (
            O => \N__33809\,
            I => \N__33806\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__33806\,
            I => \sbuttonModeStatus_0_sqmuxa_13\
        );

    \I__6238\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33800\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__33800\,
            I => \N__33797\
        );

    \I__6236\ : Span4Mux_h
    port map (
            O => \N__33797\,
            I => \N__33794\
        );

    \I__6235\ : Odrv4
    port map (
            O => \N__33794\,
            I => \sbuttonModeStatus_0_sqmuxa_22\
        );

    \I__6234\ : InMux
    port map (
            O => \N__33791\,
            I => \N__33788\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__33788\,
            I => \N__33785\
        );

    \I__6232\ : Span4Mux_h
    port map (
            O => \N__33785\,
            I => \N__33782\
        );

    \I__6231\ : Span4Mux_h
    port map (
            O => \N__33782\,
            I => \N__33779\
        );

    \I__6230\ : Span4Mux_v
    port map (
            O => \N__33779\,
            I => \N__33776\
        );

    \I__6229\ : Odrv4
    port map (
            O => \N__33776\,
            I => \sEEPonPoff_1_sqmuxa_0_a3_0_a2_1\
        );

    \I__6228\ : InMux
    port map (
            O => \N__33773\,
            I => \N__33770\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__33770\,
            I => \N__33765\
        );

    \I__6226\ : InMux
    port map (
            O => \N__33769\,
            I => \N__33762\
        );

    \I__6225\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33759\
        );

    \I__6224\ : Span4Mux_v
    port map (
            O => \N__33765\,
            I => \N__33756\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__33762\,
            I => \N__33751\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__33759\,
            I => \N__33748\
        );

    \I__6221\ : Span4Mux_h
    port map (
            O => \N__33756\,
            I => \N__33740\
        );

    \I__6220\ : InMux
    port map (
            O => \N__33755\,
            I => \N__33734\
        );

    \I__6219\ : InMux
    port map (
            O => \N__33754\,
            I => \N__33734\
        );

    \I__6218\ : Span12Mux_v
    port map (
            O => \N__33751\,
            I => \N__33729\
        );

    \I__6217\ : Span4Mux_v
    port map (
            O => \N__33748\,
            I => \N__33726\
        );

    \I__6216\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33723\
        );

    \I__6215\ : InMux
    port map (
            O => \N__33746\,
            I => \N__33718\
        );

    \I__6214\ : InMux
    port map (
            O => \N__33745\,
            I => \N__33718\
        );

    \I__6213\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33715\
        );

    \I__6212\ : InMux
    port map (
            O => \N__33743\,
            I => \N__33712\
        );

    \I__6211\ : Span4Mux_h
    port map (
            O => \N__33740\,
            I => \N__33709\
        );

    \I__6210\ : InMux
    port map (
            O => \N__33739\,
            I => \N__33706\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__33734\,
            I => \N__33703\
        );

    \I__6208\ : InMux
    port map (
            O => \N__33733\,
            I => \N__33698\
        );

    \I__6207\ : InMux
    port map (
            O => \N__33732\,
            I => \N__33698\
        );

    \I__6206\ : Odrv12
    port map (
            O => \N__33729\,
            I => \sPointer_RNI5LBD1Z0Z_0\
        );

    \I__6205\ : Odrv4
    port map (
            O => \N__33726\,
            I => \sPointer_RNI5LBD1Z0Z_0\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__33723\,
            I => \sPointer_RNI5LBD1Z0Z_0\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__33718\,
            I => \sPointer_RNI5LBD1Z0Z_0\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__33715\,
            I => \sPointer_RNI5LBD1Z0Z_0\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__33712\,
            I => \sPointer_RNI5LBD1Z0Z_0\
        );

    \I__6200\ : Odrv4
    port map (
            O => \N__33709\,
            I => \sPointer_RNI5LBD1Z0Z_0\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__33706\,
            I => \sPointer_RNI5LBD1Z0Z_0\
        );

    \I__6198\ : Odrv4
    port map (
            O => \N__33703\,
            I => \sPointer_RNI5LBD1Z0Z_0\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__33698\,
            I => \sPointer_RNI5LBD1Z0Z_0\
        );

    \I__6196\ : CEMux
    port map (
            O => \N__33677\,
            I => \N__33674\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__33674\,
            I => \sEEPonPoff_1_sqmuxa\
        );

    \I__6194\ : IoInMux
    port map (
            O => \N__33671\,
            I => \N__33668\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__33668\,
            I => \N__33665\
        );

    \I__6192\ : IoSpan4Mux
    port map (
            O => \N__33665\,
            I => \N__33662\
        );

    \I__6191\ : IoSpan4Mux
    port map (
            O => \N__33662\,
            I => \N__33659\
        );

    \I__6190\ : Span4Mux_s2_h
    port map (
            O => \N__33659\,
            I => \N__33656\
        );

    \I__6189\ : Sp12to4
    port map (
            O => \N__33656\,
            I => \N__33653\
        );

    \I__6188\ : Odrv12
    port map (
            O => \N__33653\,
            I => \RAM_nWE_0_i\
        );

    \I__6187\ : InMux
    port map (
            O => \N__33650\,
            I => \N__33647\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__33647\,
            I => \sDAC_mem_27Z0Z_0\
        );

    \I__6185\ : InMux
    port map (
            O => \N__33644\,
            I => \N__33641\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__33641\,
            I => \N__33638\
        );

    \I__6183\ : Odrv12
    port map (
            O => \N__33638\,
            I => \sDAC_mem_26Z0Z_0\
        );

    \I__6182\ : InMux
    port map (
            O => \N__33635\,
            I => \N__33632\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__33632\,
            I => \N__33629\
        );

    \I__6180\ : Span4Mux_v
    port map (
            O => \N__33629\,
            I => \N__33626\
        );

    \I__6179\ : Span4Mux_h
    port map (
            O => \N__33626\,
            I => \N__33623\
        );

    \I__6178\ : Odrv4
    port map (
            O => \N__33623\,
            I => \sDAC_mem_24Z0Z_0\
        );

    \I__6177\ : CascadeMux
    port map (
            O => \N__33620\,
            I => \sDAC_data_RNO_30Z0Z_3_cascade_\
        );

    \I__6176\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33614\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__33614\,
            I => \sDAC_data_RNO_31Z0Z_3\
        );

    \I__6174\ : InMux
    port map (
            O => \N__33611\,
            I => \N__33608\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__33608\,
            I => \sDAC_data_RNO_24Z0Z_3\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__33605\,
            I => \sDAC_data_2_39_ns_1_3_cascade_\
        );

    \I__6171\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33599\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__33599\,
            I => \N__33596\
        );

    \I__6169\ : Span4Mux_v
    port map (
            O => \N__33596\,
            I => \N__33593\
        );

    \I__6168\ : Span4Mux_v
    port map (
            O => \N__33593\,
            I => \N__33590\
        );

    \I__6167\ : Odrv4
    port map (
            O => \N__33590\,
            I => \sDAC_data_RNO_21Z0Z_7\
        );

    \I__6166\ : InMux
    port map (
            O => \N__33587\,
            I => \N__33584\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__33584\,
            I => \sDAC_mem_22Z0Z_4\
        );

    \I__6164\ : InMux
    port map (
            O => \N__33581\,
            I => \N__33578\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__33578\,
            I => \N__33575\
        );

    \I__6162\ : Span4Mux_h
    port map (
            O => \N__33575\,
            I => \N__33572\
        );

    \I__6161\ : Span4Mux_v
    port map (
            O => \N__33572\,
            I => \N__33569\
        );

    \I__6160\ : Odrv4
    port map (
            O => \N__33569\,
            I => \sDAC_data_RNO_21Z0Z_8\
        );

    \I__6159\ : InMux
    port map (
            O => \N__33566\,
            I => \N__33563\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__33563\,
            I => \sDAC_mem_22Z0Z_5\
        );

    \I__6157\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33557\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__33557\,
            I => \N__33554\
        );

    \I__6155\ : Span12Mux_v
    port map (
            O => \N__33554\,
            I => \N__33551\
        );

    \I__6154\ : Odrv12
    port map (
            O => \N__33551\,
            I => \sDAC_data_RNO_21Z0Z_9\
        );

    \I__6153\ : InMux
    port map (
            O => \N__33548\,
            I => \N__33545\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__33545\,
            I => \sDAC_data_RNO_20Z0Z_10\
        );

    \I__6151\ : CascadeMux
    port map (
            O => \N__33542\,
            I => \N__33539\
        );

    \I__6150\ : InMux
    port map (
            O => \N__33539\,
            I => \N__33536\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__33536\,
            I => \N__33533\
        );

    \I__6148\ : Span4Mux_v
    port map (
            O => \N__33533\,
            I => \N__33530\
        );

    \I__6147\ : Span4Mux_h
    port map (
            O => \N__33530\,
            I => \N__33527\
        );

    \I__6146\ : Odrv4
    port map (
            O => \N__33527\,
            I => \sDAC_mem_18Z0Z_7\
        );

    \I__6145\ : InMux
    port map (
            O => \N__33524\,
            I => \N__33521\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__33521\,
            I => \sDAC_data_RNO_29Z0Z_10\
        );

    \I__6143\ : InMux
    port map (
            O => \N__33518\,
            I => \N__33515\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__33515\,
            I => \sDAC_mem_16Z0Z_7\
        );

    \I__6141\ : CEMux
    port map (
            O => \N__33512\,
            I => \N__33509\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__33509\,
            I => \N__33505\
        );

    \I__6139\ : CEMux
    port map (
            O => \N__33508\,
            I => \N__33501\
        );

    \I__6138\ : Span4Mux_h
    port map (
            O => \N__33505\,
            I => \N__33498\
        );

    \I__6137\ : CEMux
    port map (
            O => \N__33504\,
            I => \N__33495\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__33501\,
            I => \N__33492\
        );

    \I__6135\ : Span4Mux_h
    port map (
            O => \N__33498\,
            I => \N__33487\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__33495\,
            I => \N__33487\
        );

    \I__6133\ : Span4Mux_v
    port map (
            O => \N__33492\,
            I => \N__33484\
        );

    \I__6132\ : Span4Mux_v
    port map (
            O => \N__33487\,
            I => \N__33481\
        );

    \I__6131\ : Span4Mux_h
    port map (
            O => \N__33484\,
            I => \N__33478\
        );

    \I__6130\ : Span4Mux_h
    port map (
            O => \N__33481\,
            I => \N__33475\
        );

    \I__6129\ : Odrv4
    port map (
            O => \N__33478\,
            I => \sDAC_mem_16_1_sqmuxa\
        );

    \I__6128\ : Odrv4
    port map (
            O => \N__33475\,
            I => \sDAC_mem_16_1_sqmuxa\
        );

    \I__6127\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33467\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__33467\,
            I => \sDAC_data_RNO_31Z0Z_10\
        );

    \I__6125\ : InMux
    port map (
            O => \N__33464\,
            I => \N__33461\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__33461\,
            I => \sDAC_data_RNO_30Z0Z_10\
        );

    \I__6123\ : InMux
    port map (
            O => \N__33458\,
            I => \N__33455\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__33455\,
            I => \N__33452\
        );

    \I__6121\ : Odrv12
    port map (
            O => \N__33452\,
            I => \sDAC_mem_31Z0Z_7\
        );

    \I__6120\ : InMux
    port map (
            O => \N__33449\,
            I => \N__33446\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__33446\,
            I => \N__33443\
        );

    \I__6118\ : Span4Mux_h
    port map (
            O => \N__33443\,
            I => \N__33440\
        );

    \I__6117\ : Span4Mux_h
    port map (
            O => \N__33440\,
            I => \N__33437\
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__33437\,
            I => \sDAC_mem_30Z0Z_7\
        );

    \I__6115\ : InMux
    port map (
            O => \N__33434\,
            I => \N__33431\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__33431\,
            I => \N__33428\
        );

    \I__6113\ : Span4Mux_h
    port map (
            O => \N__33428\,
            I => \N__33425\
        );

    \I__6112\ : Span4Mux_h
    port map (
            O => \N__33425\,
            I => \N__33422\
        );

    \I__6111\ : Odrv4
    port map (
            O => \N__33422\,
            I => \sDAC_mem_29Z0Z_7\
        );

    \I__6110\ : InMux
    port map (
            O => \N__33419\,
            I => \N__33416\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__33416\,
            I => \sDAC_data_RNO_24Z0Z_10\
        );

    \I__6108\ : CascadeMux
    port map (
            O => \N__33413\,
            I => \sDAC_data_RNO_23Z0Z_10_cascade_\
        );

    \I__6107\ : InMux
    port map (
            O => \N__33410\,
            I => \N__33407\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__33407\,
            I => \sDAC_data_2_39_ns_1_10\
        );

    \I__6105\ : InMux
    port map (
            O => \N__33404\,
            I => \N__33401\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__33401\,
            I => \N__33398\
        );

    \I__6103\ : Odrv4
    port map (
            O => \N__33398\,
            I => \sDAC_data_RNO_11Z0Z_10\
        );

    \I__6102\ : InMux
    port map (
            O => \N__33395\,
            I => \N__33392\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__33392\,
            I => \sDAC_mem_28Z0Z_7\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__33389\,
            I => \N__33385\
        );

    \I__6099\ : CascadeMux
    port map (
            O => \N__33388\,
            I => \N__33382\
        );

    \I__6098\ : InMux
    port map (
            O => \N__33385\,
            I => \N__33377\
        );

    \I__6097\ : InMux
    port map (
            O => \N__33382\,
            I => \N__33370\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__33381\,
            I => \N__33367\
        );

    \I__6095\ : CascadeMux
    port map (
            O => \N__33380\,
            I => \N__33363\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__33377\,
            I => \N__33359\
        );

    \I__6093\ : InMux
    port map (
            O => \N__33376\,
            I => \N__33356\
        );

    \I__6092\ : InMux
    port map (
            O => \N__33375\,
            I => \N__33353\
        );

    \I__6091\ : InMux
    port map (
            O => \N__33374\,
            I => \N__33350\
        );

    \I__6090\ : InMux
    port map (
            O => \N__33373\,
            I => \N__33347\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__33370\,
            I => \N__33344\
        );

    \I__6088\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33339\
        );

    \I__6087\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33339\
        );

    \I__6086\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33336\
        );

    \I__6085\ : InMux
    port map (
            O => \N__33362\,
            I => \N__33333\
        );

    \I__6084\ : Span4Mux_v
    port map (
            O => \N__33359\,
            I => \N__33326\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__33356\,
            I => \N__33326\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__33353\,
            I => \N__33321\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__33350\,
            I => \N__33321\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__33347\,
            I => \N__33318\
        );

    \I__6079\ : Span4Mux_h
    port map (
            O => \N__33344\,
            I => \N__33313\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__33339\,
            I => \N__33313\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__33336\,
            I => \N__33310\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__33333\,
            I => \N__33307\
        );

    \I__6075\ : InMux
    port map (
            O => \N__33332\,
            I => \N__33304\
        );

    \I__6074\ : InMux
    port map (
            O => \N__33331\,
            I => \N__33301\
        );

    \I__6073\ : Span4Mux_v
    port map (
            O => \N__33326\,
            I => \N__33294\
        );

    \I__6072\ : Span4Mux_h
    port map (
            O => \N__33321\,
            I => \N__33294\
        );

    \I__6071\ : Span4Mux_v
    port map (
            O => \N__33318\,
            I => \N__33294\
        );

    \I__6070\ : Span4Mux_v
    port map (
            O => \N__33313\,
            I => \N__33287\
        );

    \I__6069\ : Span4Mux_v
    port map (
            O => \N__33310\,
            I => \N__33287\
        );

    \I__6068\ : Span4Mux_h
    port map (
            O => \N__33307\,
            I => \N__33287\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__33304\,
            I => un7_spon_20
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__33301\,
            I => un7_spon_20
        );

    \I__6065\ : Odrv4
    port map (
            O => \N__33294\,
            I => un7_spon_20
        );

    \I__6064\ : Odrv4
    port map (
            O => \N__33287\,
            I => un7_spon_20
        );

    \I__6063\ : CascadeMux
    port map (
            O => \N__33278\,
            I => \N__33270\
        );

    \I__6062\ : InMux
    port map (
            O => \N__33277\,
            I => \N__33267\
        );

    \I__6061\ : CascadeMux
    port map (
            O => \N__33276\,
            I => \N__33264\
        );

    \I__6060\ : CascadeMux
    port map (
            O => \N__33275\,
            I => \N__33261\
        );

    \I__6059\ : CascadeMux
    port map (
            O => \N__33274\,
            I => \N__33258\
        );

    \I__6058\ : InMux
    port map (
            O => \N__33273\,
            I => \N__33254\
        );

    \I__6057\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33250\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__33267\,
            I => \N__33246\
        );

    \I__6055\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33241\
        );

    \I__6054\ : InMux
    port map (
            O => \N__33261\,
            I => \N__33241\
        );

    \I__6053\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33238\
        );

    \I__6052\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33235\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__33254\,
            I => \N__33232\
        );

    \I__6050\ : InMux
    port map (
            O => \N__33253\,
            I => \N__33229\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__33250\,
            I => \N__33226\
        );

    \I__6048\ : InMux
    port map (
            O => \N__33249\,
            I => \N__33220\
        );

    \I__6047\ : Span4Mux_v
    port map (
            O => \N__33246\,
            I => \N__33215\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__33241\,
            I => \N__33215\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__33238\,
            I => \N__33210\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__33235\,
            I => \N__33210\
        );

    \I__6043\ : Span4Mux_v
    port map (
            O => \N__33232\,
            I => \N__33205\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__33229\,
            I => \N__33205\
        );

    \I__6041\ : Span4Mux_h
    port map (
            O => \N__33226\,
            I => \N__33202\
        );

    \I__6040\ : InMux
    port map (
            O => \N__33225\,
            I => \N__33199\
        );

    \I__6039\ : InMux
    port map (
            O => \N__33224\,
            I => \N__33196\
        );

    \I__6038\ : InMux
    port map (
            O => \N__33223\,
            I => \N__33193\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__33220\,
            I => \N__33190\
        );

    \I__6036\ : Span4Mux_v
    port map (
            O => \N__33215\,
            I => \N__33181\
        );

    \I__6035\ : Span4Mux_h
    port map (
            O => \N__33210\,
            I => \N__33181\
        );

    \I__6034\ : Span4Mux_v
    port map (
            O => \N__33205\,
            I => \N__33181\
        );

    \I__6033\ : Span4Mux_v
    port map (
            O => \N__33202\,
            I => \N__33181\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__33199\,
            I => un7_spon_19
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__33196\,
            I => un7_spon_19
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__33193\,
            I => un7_spon_19
        );

    \I__6029\ : Odrv12
    port map (
            O => \N__33190\,
            I => un7_spon_19
        );

    \I__6028\ : Odrv4
    port map (
            O => \N__33181\,
            I => un7_spon_19
        );

    \I__6027\ : InMux
    port map (
            O => \N__33170\,
            I => \N__33162\
        );

    \I__6026\ : CascadeMux
    port map (
            O => \N__33169\,
            I => \N__33158\
        );

    \I__6025\ : CascadeMux
    port map (
            O => \N__33168\,
            I => \N__33155\
        );

    \I__6024\ : InMux
    port map (
            O => \N__33167\,
            I => \N__33151\
        );

    \I__6023\ : CascadeMux
    port map (
            O => \N__33166\,
            I => \N__33147\
        );

    \I__6022\ : CascadeMux
    port map (
            O => \N__33165\,
            I => \N__33144\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__33162\,
            I => \N__33141\
        );

    \I__6020\ : InMux
    port map (
            O => \N__33161\,
            I => \N__33138\
        );

    \I__6019\ : InMux
    port map (
            O => \N__33158\,
            I => \N__33135\
        );

    \I__6018\ : InMux
    port map (
            O => \N__33155\,
            I => \N__33132\
        );

    \I__6017\ : InMux
    port map (
            O => \N__33154\,
            I => \N__33129\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__33151\,
            I => \N__33126\
        );

    \I__6015\ : InMux
    port map (
            O => \N__33150\,
            I => \N__33123\
        );

    \I__6014\ : InMux
    port map (
            O => \N__33147\,
            I => \N__33120\
        );

    \I__6013\ : InMux
    port map (
            O => \N__33144\,
            I => \N__33117\
        );

    \I__6012\ : Span4Mux_v
    port map (
            O => \N__33141\,
            I => \N__33110\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__33138\,
            I => \N__33110\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__33135\,
            I => \N__33105\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__33132\,
            I => \N__33105\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__33129\,
            I => \N__33102\
        );

    \I__6007\ : Span4Mux_h
    port map (
            O => \N__33126\,
            I => \N__33097\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__33123\,
            I => \N__33097\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__33120\,
            I => \N__33094\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__33117\,
            I => \N__33091\
        );

    \I__6003\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33088\
        );

    \I__6002\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33085\
        );

    \I__6001\ : Span4Mux_v
    port map (
            O => \N__33110\,
            I => \N__33078\
        );

    \I__6000\ : Span4Mux_h
    port map (
            O => \N__33105\,
            I => \N__33078\
        );

    \I__5999\ : Span4Mux_v
    port map (
            O => \N__33102\,
            I => \N__33078\
        );

    \I__5998\ : Span4Mux_v
    port map (
            O => \N__33097\,
            I => \N__33071\
        );

    \I__5997\ : Span4Mux_v
    port map (
            O => \N__33094\,
            I => \N__33071\
        );

    \I__5996\ : Span4Mux_h
    port map (
            O => \N__33091\,
            I => \N__33071\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__33088\,
            I => un7_spon_21
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__33085\,
            I => un7_spon_21
        );

    \I__5993\ : Odrv4
    port map (
            O => \N__33078\,
            I => un7_spon_21
        );

    \I__5992\ : Odrv4
    port map (
            O => \N__33071\,
            I => un7_spon_21
        );

    \I__5991\ : CascadeMux
    port map (
            O => \N__33062\,
            I => \N__33059\
        );

    \I__5990\ : InMux
    port map (
            O => \N__33059\,
            I => \N__33054\
        );

    \I__5989\ : InMux
    port map (
            O => \N__33058\,
            I => \N__33049\
        );

    \I__5988\ : CascadeMux
    port map (
            O => \N__33057\,
            I => \N__33043\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__33054\,
            I => \N__33040\
        );

    \I__5986\ : InMux
    port map (
            O => \N__33053\,
            I => \N__33036\
        );

    \I__5985\ : InMux
    port map (
            O => \N__33052\,
            I => \N__33033\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__33049\,
            I => \N__33030\
        );

    \I__5983\ : InMux
    port map (
            O => \N__33048\,
            I => \N__33027\
        );

    \I__5982\ : InMux
    port map (
            O => \N__33047\,
            I => \N__33024\
        );

    \I__5981\ : CascadeMux
    port map (
            O => \N__33046\,
            I => \N__33021\
        );

    \I__5980\ : InMux
    port map (
            O => \N__33043\,
            I => \N__33018\
        );

    \I__5979\ : Span4Mux_v
    port map (
            O => \N__33040\,
            I => \N__33014\
        );

    \I__5978\ : InMux
    port map (
            O => \N__33039\,
            I => \N__33011\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__33036\,
            I => \N__33008\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__33033\,
            I => \N__33005\
        );

    \I__5975\ : Span4Mux_v
    port map (
            O => \N__33030\,
            I => \N__33000\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__33027\,
            I => \N__33000\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__33024\,
            I => \N__32997\
        );

    \I__5972\ : InMux
    port map (
            O => \N__33021\,
            I => \N__32994\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__33018\,
            I => \N__32991\
        );

    \I__5970\ : InMux
    port map (
            O => \N__33017\,
            I => \N__32987\
        );

    \I__5969\ : Span4Mux_v
    port map (
            O => \N__33014\,
            I => \N__32976\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__33011\,
            I => \N__32976\
        );

    \I__5967\ : Span4Mux_h
    port map (
            O => \N__33008\,
            I => \N__32976\
        );

    \I__5966\ : Span4Mux_h
    port map (
            O => \N__33005\,
            I => \N__32976\
        );

    \I__5965\ : Span4Mux_v
    port map (
            O => \N__33000\,
            I => \N__32976\
        );

    \I__5964\ : Span4Mux_h
    port map (
            O => \N__32997\,
            I => \N__32973\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__32994\,
            I => \N__32970\
        );

    \I__5962\ : Span4Mux_h
    port map (
            O => \N__32991\,
            I => \N__32967\
        );

    \I__5961\ : InMux
    port map (
            O => \N__32990\,
            I => \N__32964\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__32987\,
            I => un7_spon_11
        );

    \I__5959\ : Odrv4
    port map (
            O => \N__32976\,
            I => un7_spon_11
        );

    \I__5958\ : Odrv4
    port map (
            O => \N__32973\,
            I => un7_spon_11
        );

    \I__5957\ : Odrv12
    port map (
            O => \N__32970\,
            I => un7_spon_11
        );

    \I__5956\ : Odrv4
    port map (
            O => \N__32967\,
            I => un7_spon_11
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__32964\,
            I => un7_spon_11
        );

    \I__5954\ : CascadeMux
    port map (
            O => \N__32951\,
            I => \N__32948\
        );

    \I__5953\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32945\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__32945\,
            I => \N__32942\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__32942\,
            I => \N__32939\
        );

    \I__5950\ : Odrv4
    port map (
            O => \N__32939\,
            I => g0_12
        );

    \I__5949\ : InMux
    port map (
            O => \N__32936\,
            I => \N__32933\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__32933\,
            I => \sDAC_data_RNO_2Z0Z_10\
        );

    \I__5947\ : CascadeMux
    port map (
            O => \N__32930\,
            I => \sDAC_data_2_41_ns_1_10_cascade_\
        );

    \I__5946\ : InMux
    port map (
            O => \N__32927\,
            I => \N__32924\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__32924\,
            I => \sDAC_data_2_10\
        );

    \I__5944\ : InMux
    port map (
            O => \N__32921\,
            I => \N__32918\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__32918\,
            I => \N__32915\
        );

    \I__5942\ : Span4Mux_v
    port map (
            O => \N__32915\,
            I => \N__32912\
        );

    \I__5941\ : Odrv4
    port map (
            O => \N__32912\,
            I => \sbuttonModeStatus_0_sqmuxa_17\
        );

    \I__5940\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32906\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__32906\,
            I => \N__32903\
        );

    \I__5938\ : Span4Mux_v
    port map (
            O => \N__32903\,
            I => \N__32900\
        );

    \I__5937\ : Span4Mux_h
    port map (
            O => \N__32900\,
            I => \N__32897\
        );

    \I__5936\ : Span4Mux_h
    port map (
            O => \N__32897\,
            I => \N__32894\
        );

    \I__5935\ : Odrv4
    port map (
            O => \N__32894\,
            I => \sDAC_mem_22Z0Z_7\
        );

    \I__5934\ : CascadeMux
    port map (
            O => \N__32891\,
            I => \sDAC_data_RNO_28Z0Z_10_cascade_\
        );

    \I__5933\ : InMux
    port map (
            O => \N__32888\,
            I => \N__32885\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__32885\,
            I => \sDAC_data_RNO_21Z0Z_10\
        );

    \I__5931\ : CascadeMux
    port map (
            O => \N__32882\,
            I => \sDAC_data_2_32_ns_1_10_cascade_\
        );

    \I__5930\ : InMux
    port map (
            O => \N__32879\,
            I => \N__32876\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__32876\,
            I => \sDAC_data_RNO_10Z0Z_10\
        );

    \I__5928\ : InMux
    port map (
            O => \N__32873\,
            I => \N__32870\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__32870\,
            I => \N__32867\
        );

    \I__5926\ : Span4Mux_h
    port map (
            O => \N__32867\,
            I => \N__32864\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__32864\,
            I => \sDAC_mem_34Z0Z_7\
        );

    \I__5924\ : InMux
    port map (
            O => \N__32861\,
            I => \N__32858\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__32858\,
            I => \sDAC_mem_2Z0Z_7\
        );

    \I__5922\ : CEMux
    port map (
            O => \N__32855\,
            I => \N__32852\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__32852\,
            I => \N__32848\
        );

    \I__5920\ : CEMux
    port map (
            O => \N__32851\,
            I => \N__32845\
        );

    \I__5919\ : Span4Mux_v
    port map (
            O => \N__32848\,
            I => \N__32842\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__32845\,
            I => \N__32839\
        );

    \I__5917\ : Span4Mux_h
    port map (
            O => \N__32842\,
            I => \N__32836\
        );

    \I__5916\ : Span4Mux_h
    port map (
            O => \N__32839\,
            I => \N__32833\
        );

    \I__5915\ : Odrv4
    port map (
            O => \N__32836\,
            I => \sDAC_mem_2_1_sqmuxa\
        );

    \I__5914\ : Odrv4
    port map (
            O => \N__32833\,
            I => \sDAC_mem_2_1_sqmuxa\
        );

    \I__5913\ : InMux
    port map (
            O => \N__32828\,
            I => \N__32825\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__32825\,
            I => \N__32822\
        );

    \I__5911\ : Sp12to4
    port map (
            O => \N__32822\,
            I => \N__32819\
        );

    \I__5910\ : Span12Mux_h
    port map (
            O => \N__32819\,
            I => \N__32816\
        );

    \I__5909\ : Odrv12
    port map (
            O => \N__32816\,
            I => \sDAC_mem_12Z0Z_7\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__32813\,
            I => \sDAC_data_RNO_18Z0Z_10_cascade_\
        );

    \I__5907\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32807\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__32807\,
            I => \N__32804\
        );

    \I__5905\ : Span4Mux_v
    port map (
            O => \N__32804\,
            I => \N__32801\
        );

    \I__5904\ : Span4Mux_h
    port map (
            O => \N__32801\,
            I => \N__32798\
        );

    \I__5903\ : Odrv4
    port map (
            O => \N__32798\,
            I => \sDAC_mem_15Z0Z_7\
        );

    \I__5902\ : InMux
    port map (
            O => \N__32795\,
            I => \N__32792\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__32792\,
            I => \N__32789\
        );

    \I__5900\ : Span4Mux_v
    port map (
            O => \N__32789\,
            I => \N__32786\
        );

    \I__5899\ : Span4Mux_h
    port map (
            O => \N__32786\,
            I => \N__32783\
        );

    \I__5898\ : Odrv4
    port map (
            O => \N__32783\,
            I => \sDAC_mem_14Z0Z_7\
        );

    \I__5897\ : InMux
    port map (
            O => \N__32780\,
            I => \N__32777\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__32777\,
            I => \sDAC_data_RNO_19Z0Z_10\
        );

    \I__5895\ : InMux
    port map (
            O => \N__32774\,
            I => \N__32771\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__32771\,
            I => \N__32768\
        );

    \I__5893\ : Span4Mux_v
    port map (
            O => \N__32768\,
            I => \N__32765\
        );

    \I__5892\ : Span4Mux_h
    port map (
            O => \N__32765\,
            I => \N__32762\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__32762\,
            I => \sDAC_mem_42Z0Z_7\
        );

    \I__5890\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32756\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__32756\,
            I => \N__32753\
        );

    \I__5888\ : Span4Mux_h
    port map (
            O => \N__32753\,
            I => \N__32750\
        );

    \I__5887\ : Span4Mux_h
    port map (
            O => \N__32750\,
            I => \N__32747\
        );

    \I__5886\ : Span4Mux_v
    port map (
            O => \N__32747\,
            I => \N__32744\
        );

    \I__5885\ : Odrv4
    port map (
            O => \N__32744\,
            I => \sDAC_mem_10Z0Z_7\
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__32741\,
            I => \sDAC_data_RNO_17Z0Z_10_cascade_\
        );

    \I__5883\ : InMux
    port map (
            O => \N__32738\,
            I => \N__32735\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__32735\,
            I => \N__32732\
        );

    \I__5881\ : Span4Mux_v
    port map (
            O => \N__32732\,
            I => \N__32729\
        );

    \I__5880\ : Span4Mux_h
    port map (
            O => \N__32729\,
            I => \N__32726\
        );

    \I__5879\ : Span4Mux_h
    port map (
            O => \N__32726\,
            I => \N__32723\
        );

    \I__5878\ : Odrv4
    port map (
            O => \N__32723\,
            I => \sDAC_mem_11Z0Z_7\
        );

    \I__5877\ : InMux
    port map (
            O => \N__32720\,
            I => \N__32717\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__32717\,
            I => \sDAC_data_2_24_ns_1_10\
        );

    \I__5875\ : CascadeMux
    port map (
            O => \N__32714\,
            I => \sDAC_data_RNO_8Z0Z_10_cascade_\
        );

    \I__5874\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32708\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__32708\,
            I => \N__32705\
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__32705\,
            I => \sDAC_data_RNO_7Z0Z_10\
        );

    \I__5871\ : CascadeMux
    port map (
            O => \N__32702\,
            I => \sDAC_data_2_20_am_1_10_cascade_\
        );

    \I__5870\ : InMux
    port map (
            O => \N__32699\,
            I => \N__32696\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__32696\,
            I => \N__32693\
        );

    \I__5868\ : Span4Mux_v
    port map (
            O => \N__32693\,
            I => \N__32690\
        );

    \I__5867\ : Odrv4
    port map (
            O => \N__32690\,
            I => \sDAC_mem_36Z0Z_6\
        );

    \I__5866\ : CascadeMux
    port map (
            O => \N__32687\,
            I => \sDAC_data_2_13_am_1_9_cascade_\
        );

    \I__5865\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32681\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__32681\,
            I => \N__32678\
        );

    \I__5863\ : Span4Mux_h
    port map (
            O => \N__32678\,
            I => \N__32675\
        );

    \I__5862\ : Odrv4
    port map (
            O => \N__32675\,
            I => \sDAC_data_RNO_4Z0Z_9\
        );

    \I__5861\ : CascadeMux
    port map (
            O => \N__32672\,
            I => \N__32669\
        );

    \I__5860\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32666\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__32666\,
            I => \sDAC_mem_4Z0Z_6\
        );

    \I__5858\ : InMux
    port map (
            O => \N__32663\,
            I => \N__32660\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__32660\,
            I => \N__32657\
        );

    \I__5856\ : Span4Mux_h
    port map (
            O => \N__32657\,
            I => \N__32654\
        );

    \I__5855\ : Span4Mux_v
    port map (
            O => \N__32654\,
            I => \N__32651\
        );

    \I__5854\ : Odrv4
    port map (
            O => \N__32651\,
            I => \sDAC_mem_38Z0Z_7\
        );

    \I__5853\ : InMux
    port map (
            O => \N__32648\,
            I => \N__32645\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__32645\,
            I => \N__32642\
        );

    \I__5851\ : Span4Mux_v
    port map (
            O => \N__32642\,
            I => \N__32639\
        );

    \I__5850\ : Odrv4
    port map (
            O => \N__32639\,
            I => \sDAC_mem_39Z0Z_7\
        );

    \I__5849\ : CascadeMux
    port map (
            O => \N__32636\,
            I => \sDAC_data_2_13_bm_1_10_cascade_\
        );

    \I__5848\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32630\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__32630\,
            I => \N__32627\
        );

    \I__5846\ : Span4Mux_h
    port map (
            O => \N__32627\,
            I => \N__32624\
        );

    \I__5845\ : Odrv4
    port map (
            O => \N__32624\,
            I => \sDAC_mem_7Z0Z_7\
        );

    \I__5844\ : InMux
    port map (
            O => \N__32621\,
            I => \N__32618\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__32618\,
            I => \N__32615\
        );

    \I__5842\ : Span4Mux_h
    port map (
            O => \N__32615\,
            I => \N__32612\
        );

    \I__5841\ : Span4Mux_v
    port map (
            O => \N__32612\,
            I => \N__32609\
        );

    \I__5840\ : Odrv4
    port map (
            O => \N__32609\,
            I => \sDAC_mem_38Z0Z_0\
        );

    \I__5839\ : InMux
    port map (
            O => \N__32606\,
            I => \N__32603\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__32603\,
            I => \N__32600\
        );

    \I__5837\ : Span4Mux_v
    port map (
            O => \N__32600\,
            I => \N__32597\
        );

    \I__5836\ : Odrv4
    port map (
            O => \N__32597\,
            I => \sDAC_mem_39Z0Z_0\
        );

    \I__5835\ : CascadeMux
    port map (
            O => \N__32594\,
            I => \sDAC_data_2_13_bm_1_3_cascade_\
        );

    \I__5834\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32588\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__32588\,
            I => \N__32585\
        );

    \I__5832\ : Span12Mux_h
    port map (
            O => \N__32585\,
            I => \N__32582\
        );

    \I__5831\ : Odrv12
    port map (
            O => \N__32582\,
            I => \sDAC_mem_7Z0Z_0\
        );

    \I__5830\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32576\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__32576\,
            I => \N__32573\
        );

    \I__5828\ : Span4Mux_h
    port map (
            O => \N__32573\,
            I => \N__32570\
        );

    \I__5827\ : Span4Mux_v
    port map (
            O => \N__32570\,
            I => \N__32567\
        );

    \I__5826\ : Odrv4
    port map (
            O => \N__32567\,
            I => \sDAC_mem_38Z0Z_1\
        );

    \I__5825\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32561\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__32561\,
            I => \N__32558\
        );

    \I__5823\ : Span4Mux_h
    port map (
            O => \N__32558\,
            I => \N__32555\
        );

    \I__5822\ : Odrv4
    port map (
            O => \N__32555\,
            I => \sDAC_data_2_13_bm_1_4\
        );

    \I__5821\ : CascadeMux
    port map (
            O => \N__32552\,
            I => \sDAC_data_2_13_am_1_8_cascade_\
        );

    \I__5820\ : InMux
    port map (
            O => \N__32549\,
            I => \N__32546\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__32546\,
            I => \N__32543\
        );

    \I__5818\ : Span4Mux_h
    port map (
            O => \N__32543\,
            I => \N__32540\
        );

    \I__5817\ : Odrv4
    port map (
            O => \N__32540\,
            I => \sDAC_data_RNO_4Z0Z_8\
        );

    \I__5816\ : InMux
    port map (
            O => \N__32537\,
            I => \N__32534\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__32534\,
            I => \N__32531\
        );

    \I__5814\ : Span4Mux_h
    port map (
            O => \N__32531\,
            I => \N__32528\
        );

    \I__5813\ : Span4Mux_h
    port map (
            O => \N__32528\,
            I => \N__32525\
        );

    \I__5812\ : Odrv4
    port map (
            O => \N__32525\,
            I => \sDAC_mem_38Z0Z_5\
        );

    \I__5811\ : InMux
    port map (
            O => \N__32522\,
            I => \N__32519\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__32519\,
            I => \N__32516\
        );

    \I__5809\ : Odrv4
    port map (
            O => \N__32516\,
            I => \sDAC_mem_39Z0Z_5\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__32513\,
            I => \sDAC_data_2_13_bm_1_8_cascade_\
        );

    \I__5807\ : InMux
    port map (
            O => \N__32510\,
            I => \N__32507\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__32507\,
            I => \N__32504\
        );

    \I__5805\ : Span4Mux_h
    port map (
            O => \N__32504\,
            I => \N__32501\
        );

    \I__5804\ : Odrv4
    port map (
            O => \N__32501\,
            I => \sDAC_mem_7Z0Z_5\
        );

    \I__5803\ : InMux
    port map (
            O => \N__32498\,
            I => \N__32495\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__32495\,
            I => \N__32492\
        );

    \I__5801\ : Span4Mux_v
    port map (
            O => \N__32492\,
            I => \N__32489\
        );

    \I__5800\ : Odrv4
    port map (
            O => \N__32489\,
            I => \sDAC_data_RNO_5Z0Z_8\
        );

    \I__5799\ : InMux
    port map (
            O => \N__32486\,
            I => \N__32483\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__32483\,
            I => \sDAC_mem_6Z0Z_5\
        );

    \I__5797\ : InMux
    port map (
            O => \N__32480\,
            I => \N__32477\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__32477\,
            I => \N__32474\
        );

    \I__5795\ : Span4Mux_h
    port map (
            O => \N__32474\,
            I => \N__32471\
        );

    \I__5794\ : Span4Mux_h
    port map (
            O => \N__32471\,
            I => \N__32468\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__32468\,
            I => \sDAC_mem_38Z0Z_6\
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__32465\,
            I => \sDAC_data_2_13_bm_1_9_cascade_\
        );

    \I__5791\ : InMux
    port map (
            O => \N__32462\,
            I => \N__32459\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__32459\,
            I => \N__32456\
        );

    \I__5789\ : Odrv12
    port map (
            O => \N__32456\,
            I => \sDAC_mem_39Z0Z_6\
        );

    \I__5788\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32450\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__32450\,
            I => \N__32447\
        );

    \I__5786\ : Odrv4
    port map (
            O => \N__32447\,
            I => \sDAC_data_RNO_5Z0Z_9\
        );

    \I__5785\ : InMux
    port map (
            O => \N__32444\,
            I => \N__32441\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__32441\,
            I => \sDAC_mem_6Z0Z_6\
        );

    \I__5783\ : InMux
    port map (
            O => \N__32438\,
            I => \N__32435\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__32435\,
            I => \N__32432\
        );

    \I__5781\ : Span4Mux_h
    port map (
            O => \N__32432\,
            I => \N__32429\
        );

    \I__5780\ : Span4Mux_v
    port map (
            O => \N__32429\,
            I => \N__32426\
        );

    \I__5779\ : Odrv4
    port map (
            O => \N__32426\,
            I => \sDAC_mem_40Z0Z_7\
        );

    \I__5778\ : InMux
    port map (
            O => \N__32423\,
            I => \N__32420\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__32420\,
            I => \N__32417\
        );

    \I__5776\ : Span4Mux_v
    port map (
            O => \N__32417\,
            I => \N__32414\
        );

    \I__5775\ : Span4Mux_h
    port map (
            O => \N__32414\,
            I => \N__32411\
        );

    \I__5774\ : Odrv4
    port map (
            O => \N__32411\,
            I => \sDAC_mem_8Z0Z_7\
        );

    \I__5773\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32405\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__32405\,
            I => \N__32402\
        );

    \I__5771\ : Sp12to4
    port map (
            O => \N__32402\,
            I => \N__32399\
        );

    \I__5770\ : Odrv12
    port map (
            O => \N__32399\,
            I => \sDAC_mem_22Z0Z_0\
        );

    \I__5769\ : InMux
    port map (
            O => \N__32396\,
            I => \N__32393\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__32393\,
            I => \N__32390\
        );

    \I__5767\ : Sp12to4
    port map (
            O => \N__32390\,
            I => \N__32387\
        );

    \I__5766\ : Odrv12
    port map (
            O => \N__32387\,
            I => \sDAC_mem_22Z0Z_1\
        );

    \I__5765\ : InMux
    port map (
            O => \N__32384\,
            I => \N__32381\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__32381\,
            I => \sDAC_data_RNO_21Z0Z_4\
        );

    \I__5763\ : InMux
    port map (
            O => \N__32378\,
            I => \N__32375\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__32375\,
            I => \N__32372\
        );

    \I__5761\ : Span12Mux_h
    port map (
            O => \N__32372\,
            I => \N__32369\
        );

    \I__5760\ : Odrv12
    port map (
            O => \N__32369\,
            I => \sDAC_mem_22Z0Z_2\
        );

    \I__5759\ : InMux
    port map (
            O => \N__32366\,
            I => \N__32363\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__32363\,
            I => \N__32360\
        );

    \I__5757\ : Span12Mux_h
    port map (
            O => \N__32360\,
            I => \N__32357\
        );

    \I__5756\ : Odrv12
    port map (
            O => \N__32357\,
            I => \sDAC_mem_22Z0Z_3\
        );

    \I__5755\ : InMux
    port map (
            O => \N__32354\,
            I => \N__32351\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__32351\,
            I => \N__32348\
        );

    \I__5753\ : Span4Mux_h
    port map (
            O => \N__32348\,
            I => \N__32345\
        );

    \I__5752\ : Odrv4
    port map (
            O => \N__32345\,
            I => \sDAC_data_RNO_21Z0Z_6\
        );

    \I__5751\ : InMux
    port map (
            O => \N__32342\,
            I => \N__32339\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__32339\,
            I => \N__32336\
        );

    \I__5749\ : Span4Mux_v
    port map (
            O => \N__32336\,
            I => \N__32333\
        );

    \I__5748\ : Odrv4
    port map (
            O => \N__32333\,
            I => \sDAC_mem_36Z0Z_4\
        );

    \I__5747\ : CascadeMux
    port map (
            O => \N__32330\,
            I => \sDAC_data_2_13_am_1_7_cascade_\
        );

    \I__5746\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32324\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__32324\,
            I => \N__32321\
        );

    \I__5744\ : Odrv4
    port map (
            O => \N__32321\,
            I => \sDAC_data_RNO_4Z0Z_7\
        );

    \I__5743\ : InMux
    port map (
            O => \N__32318\,
            I => \N__32315\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__32315\,
            I => \sDAC_mem_4Z0Z_4\
        );

    \I__5741\ : InMux
    port map (
            O => \N__32312\,
            I => \N__32309\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__32309\,
            I => \N__32306\
        );

    \I__5739\ : Span4Mux_v
    port map (
            O => \N__32306\,
            I => \N__32303\
        );

    \I__5738\ : Odrv4
    port map (
            O => \N__32303\,
            I => \sDAC_mem_36Z0Z_5\
        );

    \I__5737\ : InMux
    port map (
            O => \N__32300\,
            I => \N__32297\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__32297\,
            I => \N__32294\
        );

    \I__5735\ : Odrv4
    port map (
            O => \N__32294\,
            I => \sEEDACZ0Z_6\
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__32291\,
            I => \sDAC_data_2_9_cascade_\
        );

    \I__5733\ : InMux
    port map (
            O => \N__32288\,
            I => \N__32285\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__32285\,
            I => \N__32282\
        );

    \I__5731\ : Odrv4
    port map (
            O => \N__32282\,
            I => \sDAC_dataZ0Z_9\
        );

    \I__5730\ : InMux
    port map (
            O => \N__32279\,
            I => \N__32276\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__32276\,
            I => \sDAC_data_2_14_ns_1_9\
        );

    \I__5728\ : InMux
    port map (
            O => \N__32273\,
            I => \N__32270\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__32270\,
            I => \N__32267\
        );

    \I__5726\ : Odrv4
    port map (
            O => \N__32267\,
            I => \sDAC_data_RNO_29Z0Z_9\
        );

    \I__5725\ : InMux
    port map (
            O => \N__32264\,
            I => \N__32261\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__32261\,
            I => \sDAC_data_RNO_28Z0Z_9\
        );

    \I__5723\ : CascadeMux
    port map (
            O => \N__32258\,
            I => \sDAC_data_2_32_ns_1_9_cascade_\
        );

    \I__5722\ : CascadeMux
    port map (
            O => \N__32255\,
            I => \sDAC_data_RNO_10Z0Z_9_cascade_\
        );

    \I__5721\ : InMux
    port map (
            O => \N__32252\,
            I => \N__32249\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__32249\,
            I => \N__32246\
        );

    \I__5719\ : Span4Mux_h
    port map (
            O => \N__32246\,
            I => \N__32243\
        );

    \I__5718\ : Span4Mux_v
    port map (
            O => \N__32243\,
            I => \N__32240\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__32240\,
            I => \sDAC_data_RNO_11Z0Z_9\
        );

    \I__5716\ : InMux
    port map (
            O => \N__32237\,
            I => \N__32234\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__32234\,
            I => \sDAC_data_2_41_ns_1_9\
        );

    \I__5714\ : InMux
    port map (
            O => \N__32231\,
            I => \N__32228\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__32228\,
            I => \N__32225\
        );

    \I__5712\ : Odrv4
    port map (
            O => \N__32225\,
            I => \sDAC_data_RNO_20Z0Z_8\
        );

    \I__5711\ : InMux
    port map (
            O => \N__32222\,
            I => \N__32219\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__32219\,
            I => \sDAC_mem_20Z0Z_5\
        );

    \I__5709\ : InMux
    port map (
            O => \N__32216\,
            I => \N__32213\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__32213\,
            I => \sDAC_data_RNO_20Z0Z_9\
        );

    \I__5707\ : InMux
    port map (
            O => \N__32210\,
            I => \N__32207\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__32207\,
            I => \sDAC_mem_20Z0Z_6\
        );

    \I__5705\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32201\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__32201\,
            I => \sDAC_data_RNO_29Z0Z_7\
        );

    \I__5703\ : InMux
    port map (
            O => \N__32198\,
            I => \N__32195\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__32195\,
            I => \N__32192\
        );

    \I__5701\ : Odrv4
    port map (
            O => \N__32192\,
            I => \sDAC_data_RNO_28Z0Z_7\
        );

    \I__5700\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32186\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__32186\,
            I => \sDAC_data_2_32_ns_1_7\
        );

    \I__5698\ : CascadeMux
    port map (
            O => \N__32183\,
            I => \sDAC_data_2_14_ns_1_7_cascade_\
        );

    \I__5697\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32177\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__32177\,
            I => \sDAC_data_RNO_5Z0Z_7\
        );

    \I__5695\ : InMux
    port map (
            O => \N__32174\,
            I => \N__32171\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__32171\,
            I => \N__32168\
        );

    \I__5693\ : Span4Mux_v
    port map (
            O => \N__32168\,
            I => \N__32165\
        );

    \I__5692\ : Span4Mux_v
    port map (
            O => \N__32165\,
            I => \N__32162\
        );

    \I__5691\ : Odrv4
    port map (
            O => \N__32162\,
            I => \sDAC_data_RNO_11Z0Z_7\
        );

    \I__5690\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32156\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__32156\,
            I => \sDAC_data_RNO_10Z0Z_7\
        );

    \I__5688\ : CascadeMux
    port map (
            O => \N__32153\,
            I => \sDAC_data_2_41_ns_1_7_cascade_\
        );

    \I__5687\ : InMux
    port map (
            O => \N__32150\,
            I => \N__32147\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__32147\,
            I => \sDAC_data_RNO_1Z0Z_7\
        );

    \I__5685\ : InMux
    port map (
            O => \N__32144\,
            I => \N__32141\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__32141\,
            I => \N__32138\
        );

    \I__5683\ : Odrv4
    port map (
            O => \N__32138\,
            I => \sEEDACZ0Z_4\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__32135\,
            I => \sDAC_data_2_7_cascade_\
        );

    \I__5681\ : InMux
    port map (
            O => \N__32132\,
            I => \N__32129\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__32129\,
            I => \N__32126\
        );

    \I__5679\ : Odrv4
    port map (
            O => \N__32126\,
            I => \sDAC_dataZ0Z_7\
        );

    \I__5678\ : CascadeMux
    port map (
            O => \N__32123\,
            I => \sDAC_data_RNO_1Z0Z_9_cascade_\
        );

    \I__5677\ : InMux
    port map (
            O => \N__32120\,
            I => \N__32117\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__32117\,
            I => \N__32114\
        );

    \I__5675\ : Odrv4
    port map (
            O => \N__32114\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_9\
        );

    \I__5674\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32108\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__32108\,
            I => \N__32105\
        );

    \I__5672\ : Span4Mux_v
    port map (
            O => \N__32105\,
            I => \N__32102\
        );

    \I__5671\ : Odrv4
    port map (
            O => \N__32102\,
            I => \sEEDACZ0Z_1\
        );

    \I__5670\ : InMux
    port map (
            O => \N__32099\,
            I => \N__32096\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__32096\,
            I => \N__32093\
        );

    \I__5668\ : Span4Mux_h
    port map (
            O => \N__32093\,
            I => \N__32090\
        );

    \I__5667\ : Odrv4
    port map (
            O => \N__32090\,
            I => \sEEDACZ0Z_3\
        );

    \I__5666\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32084\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__32084\,
            I => \N__32081\
        );

    \I__5664\ : Span4Mux_v
    port map (
            O => \N__32081\,
            I => \N__32078\
        );

    \I__5663\ : Span4Mux_h
    port map (
            O => \N__32078\,
            I => \N__32075\
        );

    \I__5662\ : Odrv4
    port map (
            O => \N__32075\,
            I => \sEEDACZ0Z_5\
        );

    \I__5661\ : InMux
    port map (
            O => \N__32072\,
            I => \N__32069\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__32069\,
            I => \N__32066\
        );

    \I__5659\ : Span4Mux_v
    port map (
            O => \N__32066\,
            I => \N__32063\
        );

    \I__5658\ : Span4Mux_v
    port map (
            O => \N__32063\,
            I => \N__32060\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__32060\,
            I => \sEEDACZ0Z_7\
        );

    \I__5656\ : CEMux
    port map (
            O => \N__32057\,
            I => \N__32054\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__32054\,
            I => \N__32051\
        );

    \I__5654\ : Odrv4
    port map (
            O => \N__32051\,
            I => \sEEDAC_1_sqmuxa\
        );

    \I__5653\ : CascadeMux
    port map (
            O => \N__32048\,
            I => \N__32042\
        );

    \I__5652\ : CascadeMux
    port map (
            O => \N__32047\,
            I => \N__32038\
        );

    \I__5651\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32034\
        );

    \I__5650\ : InMux
    port map (
            O => \N__32045\,
            I => \N__32031\
        );

    \I__5649\ : InMux
    port map (
            O => \N__32042\,
            I => \N__32028\
        );

    \I__5648\ : CascadeMux
    port map (
            O => \N__32041\,
            I => \N__32024\
        );

    \I__5647\ : InMux
    port map (
            O => \N__32038\,
            I => \N__32021\
        );

    \I__5646\ : InMux
    port map (
            O => \N__32037\,
            I => \N__32015\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__32034\,
            I => \N__32010\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__32031\,
            I => \N__32010\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__32028\,
            I => \N__32007\
        );

    \I__5642\ : InMux
    port map (
            O => \N__32027\,
            I => \N__32004\
        );

    \I__5641\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32001\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__32021\,
            I => \N__31998\
        );

    \I__5639\ : InMux
    port map (
            O => \N__32020\,
            I => \N__31995\
        );

    \I__5638\ : InMux
    port map (
            O => \N__32019\,
            I => \N__31992\
        );

    \I__5637\ : InMux
    port map (
            O => \N__32018\,
            I => \N__31987\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__32015\,
            I => \N__31984\
        );

    \I__5635\ : Span4Mux_v
    port map (
            O => \N__32010\,
            I => \N__31981\
        );

    \I__5634\ : Span4Mux_v
    port map (
            O => \N__32007\,
            I => \N__31976\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__32004\,
            I => \N__31976\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__32001\,
            I => \N__31973\
        );

    \I__5631\ : Span4Mux_h
    port map (
            O => \N__31998\,
            I => \N__31966\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__31995\,
            I => \N__31966\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__31992\,
            I => \N__31966\
        );

    \I__5628\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31963\
        );

    \I__5627\ : InMux
    port map (
            O => \N__31990\,
            I => \N__31960\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__31987\,
            I => \N__31951\
        );

    \I__5625\ : Span4Mux_h
    port map (
            O => \N__31984\,
            I => \N__31951\
        );

    \I__5624\ : Span4Mux_h
    port map (
            O => \N__31981\,
            I => \N__31951\
        );

    \I__5623\ : Span4Mux_v
    port map (
            O => \N__31976\,
            I => \N__31951\
        );

    \I__5622\ : Span4Mux_v
    port map (
            O => \N__31973\,
            I => \N__31946\
        );

    \I__5621\ : Span4Mux_v
    port map (
            O => \N__31966\,
            I => \N__31946\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__31963\,
            I => un7_spon_22
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__31960\,
            I => un7_spon_22
        );

    \I__5618\ : Odrv4
    port map (
            O => \N__31951\,
            I => un7_spon_22
        );

    \I__5617\ : Odrv4
    port map (
            O => \N__31946\,
            I => un7_spon_22
        );

    \I__5616\ : CascadeMux
    port map (
            O => \N__31937\,
            I => \N__31931\
        );

    \I__5615\ : CascadeMux
    port map (
            O => \N__31936\,
            I => \N__31926\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__31935\,
            I => \N__31923\
        );

    \I__5613\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31920\
        );

    \I__5612\ : InMux
    port map (
            O => \N__31931\,
            I => \N__31917\
        );

    \I__5611\ : CascadeMux
    port map (
            O => \N__31930\,
            I => \N__31914\
        );

    \I__5610\ : InMux
    port map (
            O => \N__31929\,
            I => \N__31910\
        );

    \I__5609\ : InMux
    port map (
            O => \N__31926\,
            I => \N__31906\
        );

    \I__5608\ : InMux
    port map (
            O => \N__31923\,
            I => \N__31902\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__31920\,
            I => \N__31899\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__31917\,
            I => \N__31896\
        );

    \I__5605\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31893\
        );

    \I__5604\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31890\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__31910\,
            I => \N__31887\
        );

    \I__5602\ : InMux
    port map (
            O => \N__31909\,
            I => \N__31884\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__31906\,
            I => \N__31879\
        );

    \I__5600\ : CascadeMux
    port map (
            O => \N__31905\,
            I => \N__31876\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__31902\,
            I => \N__31873\
        );

    \I__5598\ : Span4Mux_v
    port map (
            O => \N__31899\,
            I => \N__31866\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__31896\,
            I => \N__31866\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__31893\,
            I => \N__31866\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__31890\,
            I => \N__31863\
        );

    \I__5594\ : Span4Mux_h
    port map (
            O => \N__31887\,
            I => \N__31858\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__31884\,
            I => \N__31858\
        );

    \I__5592\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31855\
        );

    \I__5591\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31852\
        );

    \I__5590\ : Span4Mux_h
    port map (
            O => \N__31879\,
            I => \N__31849\
        );

    \I__5589\ : InMux
    port map (
            O => \N__31876\,
            I => \N__31846\
        );

    \I__5588\ : Span4Mux_v
    port map (
            O => \N__31873\,
            I => \N__31843\
        );

    \I__5587\ : Span4Mux_v
    port map (
            O => \N__31866\,
            I => \N__31838\
        );

    \I__5586\ : Span4Mux_v
    port map (
            O => \N__31863\,
            I => \N__31838\
        );

    \I__5585\ : Span4Mux_v
    port map (
            O => \N__31858\,
            I => \N__31835\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__31855\,
            I => un7_spon_23
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__31852\,
            I => un7_spon_23
        );

    \I__5582\ : Odrv4
    port map (
            O => \N__31849\,
            I => un7_spon_23
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__31846\,
            I => un7_spon_23
        );

    \I__5580\ : Odrv4
    port map (
            O => \N__31843\,
            I => un7_spon_23
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__31838\,
            I => un7_spon_23
        );

    \I__5578\ : Odrv4
    port map (
            O => \N__31835\,
            I => un7_spon_23
        );

    \I__5577\ : InMux
    port map (
            O => \N__31820\,
            I => \bfn_14_20_0_\
        );

    \I__5576\ : InMux
    port map (
            O => \N__31817\,
            I => \N__31814\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__31814\,
            I => \N__31811\
        );

    \I__5574\ : Span4Mux_v
    port map (
            O => \N__31811\,
            I => \N__31808\
        );

    \I__5573\ : Span4Mux_v
    port map (
            O => \N__31808\,
            I => \N__31805\
        );

    \I__5572\ : Odrv4
    port map (
            O => \N__31805\,
            I => \un4_spoff_cry_23_THRU_CO\
        );

    \I__5571\ : InMux
    port map (
            O => \N__31802\,
            I => \N__31799\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__31799\,
            I => \N__31796\
        );

    \I__5569\ : Odrv12
    port map (
            O => \N__31796\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_3\
        );

    \I__5568\ : InMux
    port map (
            O => \N__31793\,
            I => \N__31790\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__31790\,
            I => \N__31787\
        );

    \I__5566\ : Span4Mux_h
    port map (
            O => \N__31787\,
            I => \N__31784\
        );

    \I__5565\ : Span4Mux_v
    port map (
            O => \N__31784\,
            I => \N__31781\
        );

    \I__5564\ : Odrv4
    port map (
            O => \N__31781\,
            I => \sDAC_dataZ0Z_4\
        );

    \I__5563\ : InMux
    port map (
            O => \N__31778\,
            I => \N__31775\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__31775\,
            I => \N__31772\
        );

    \I__5561\ : Odrv12
    port map (
            O => \N__31772\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_4\
        );

    \I__5560\ : InMux
    port map (
            O => \N__31769\,
            I => \N__31766\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__31766\,
            I => \N__31763\
        );

    \I__5558\ : Odrv4
    port map (
            O => \N__31763\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_7\
        );

    \I__5557\ : InMux
    port map (
            O => \N__31760\,
            I => \N__31757\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__31757\,
            I => \N__31754\
        );

    \I__5555\ : Span4Mux_h
    port map (
            O => \N__31754\,
            I => \N__31751\
        );

    \I__5554\ : Odrv4
    port map (
            O => \N__31751\,
            I => \sDAC_dataZ0Z_8\
        );

    \I__5553\ : CascadeMux
    port map (
            O => \N__31748\,
            I => \N__31744\
        );

    \I__5552\ : InMux
    port map (
            O => \N__31747\,
            I => \N__31740\
        );

    \I__5551\ : InMux
    port map (
            O => \N__31744\,
            I => \N__31737\
        );

    \I__5550\ : CascadeMux
    port map (
            O => \N__31743\,
            I => \N__31734\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__31740\,
            I => \N__31729\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__31737\,
            I => \N__31726\
        );

    \I__5547\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31723\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__31733\,
            I => \N__31719\
        );

    \I__5545\ : InMux
    port map (
            O => \N__31732\,
            I => \N__31714\
        );

    \I__5544\ : Span4Mux_h
    port map (
            O => \N__31729\,
            I => \N__31707\
        );

    \I__5543\ : Span4Mux_h
    port map (
            O => \N__31726\,
            I => \N__31707\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__31723\,
            I => \N__31707\
        );

    \I__5541\ : InMux
    port map (
            O => \N__31722\,
            I => \N__31704\
        );

    \I__5540\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31701\
        );

    \I__5539\ : InMux
    port map (
            O => \N__31718\,
            I => \N__31697\
        );

    \I__5538\ : InMux
    port map (
            O => \N__31717\,
            I => \N__31694\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__31714\,
            I => \N__31691\
        );

    \I__5536\ : Span4Mux_v
    port map (
            O => \N__31707\,
            I => \N__31688\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__31704\,
            I => \N__31685\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__31701\,
            I => \N__31682\
        );

    \I__5533\ : InMux
    port map (
            O => \N__31700\,
            I => \N__31679\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__31697\,
            I => un7_spon_12
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__31694\,
            I => un7_spon_12
        );

    \I__5530\ : Odrv12
    port map (
            O => \N__31691\,
            I => un7_spon_12
        );

    \I__5529\ : Odrv4
    port map (
            O => \N__31688\,
            I => un7_spon_12
        );

    \I__5528\ : Odrv4
    port map (
            O => \N__31685\,
            I => un7_spon_12
        );

    \I__5527\ : Odrv12
    port map (
            O => \N__31682\,
            I => un7_spon_12
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__31679\,
            I => un7_spon_12
        );

    \I__5525\ : CascadeMux
    port map (
            O => \N__31664\,
            I => \N__31661\
        );

    \I__5524\ : InMux
    port map (
            O => \N__31661\,
            I => \N__31655\
        );

    \I__5523\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31652\
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__31659\,
            I => \N__31649\
        );

    \I__5521\ : CascadeMux
    port map (
            O => \N__31658\,
            I => \N__31646\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__31655\,
            I => \N__31640\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__31652\,
            I => \N__31637\
        );

    \I__5518\ : InMux
    port map (
            O => \N__31649\,
            I => \N__31634\
        );

    \I__5517\ : InMux
    port map (
            O => \N__31646\,
            I => \N__31631\
        );

    \I__5516\ : InMux
    port map (
            O => \N__31645\,
            I => \N__31627\
        );

    \I__5515\ : InMux
    port map (
            O => \N__31644\,
            I => \N__31624\
        );

    \I__5514\ : InMux
    port map (
            O => \N__31643\,
            I => \N__31621\
        );

    \I__5513\ : Span4Mux_h
    port map (
            O => \N__31640\,
            I => \N__31614\
        );

    \I__5512\ : Span4Mux_h
    port map (
            O => \N__31637\,
            I => \N__31614\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__31634\,
            I => \N__31614\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__31631\,
            I => \N__31611\
        );

    \I__5509\ : InMux
    port map (
            O => \N__31630\,
            I => \N__31607\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__31627\,
            I => \N__31602\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__31624\,
            I => \N__31602\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__31621\,
            I => \N__31599\
        );

    \I__5505\ : Span4Mux_v
    port map (
            O => \N__31614\,
            I => \N__31594\
        );

    \I__5504\ : Span4Mux_v
    port map (
            O => \N__31611\,
            I => \N__31594\
        );

    \I__5503\ : InMux
    port map (
            O => \N__31610\,
            I => \N__31591\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__31607\,
            I => un7_spon_13
        );

    \I__5501\ : Odrv12
    port map (
            O => \N__31602\,
            I => un7_spon_13
        );

    \I__5500\ : Odrv4
    port map (
            O => \N__31599\,
            I => un7_spon_13
        );

    \I__5499\ : Odrv4
    port map (
            O => \N__31594\,
            I => un7_spon_13
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__31591\,
            I => un7_spon_13
        );

    \I__5497\ : CascadeMux
    port map (
            O => \N__31580\,
            I => \N__31575\
        );

    \I__5496\ : CascadeMux
    port map (
            O => \N__31579\,
            I => \N__31570\
        );

    \I__5495\ : InMux
    port map (
            O => \N__31578\,
            I => \N__31566\
        );

    \I__5494\ : InMux
    port map (
            O => \N__31575\,
            I => \N__31563\
        );

    \I__5493\ : CascadeMux
    port map (
            O => \N__31574\,
            I => \N__31560\
        );

    \I__5492\ : CascadeMux
    port map (
            O => \N__31573\,
            I => \N__31557\
        );

    \I__5491\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31554\
        );

    \I__5490\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31551\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__31566\,
            I => \N__31547\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__31563\,
            I => \N__31544\
        );

    \I__5487\ : InMux
    port map (
            O => \N__31560\,
            I => \N__31541\
        );

    \I__5486\ : InMux
    port map (
            O => \N__31557\,
            I => \N__31538\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__31554\,
            I => \N__31534\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__31551\,
            I => \N__31531\
        );

    \I__5483\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31528\
        );

    \I__5482\ : Span4Mux_h
    port map (
            O => \N__31547\,
            I => \N__31521\
        );

    \I__5481\ : Span4Mux_h
    port map (
            O => \N__31544\,
            I => \N__31521\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__31541\,
            I => \N__31521\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__31538\,
            I => \N__31518\
        );

    \I__5478\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31514\
        );

    \I__5477\ : Span4Mux_h
    port map (
            O => \N__31534\,
            I => \N__31511\
        );

    \I__5476\ : Span4Mux_h
    port map (
            O => \N__31531\,
            I => \N__31508\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__31528\,
            I => \N__31505\
        );

    \I__5474\ : Span4Mux_v
    port map (
            O => \N__31521\,
            I => \N__31500\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__31518\,
            I => \N__31500\
        );

    \I__5472\ : InMux
    port map (
            O => \N__31517\,
            I => \N__31497\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__31514\,
            I => un7_spon_14
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__31511\,
            I => un7_spon_14
        );

    \I__5469\ : Odrv4
    port map (
            O => \N__31508\,
            I => un7_spon_14
        );

    \I__5468\ : Odrv4
    port map (
            O => \N__31505\,
            I => un7_spon_14
        );

    \I__5467\ : Odrv4
    port map (
            O => \N__31500\,
            I => un7_spon_14
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__31497\,
            I => un7_spon_14
        );

    \I__5465\ : CascadeMux
    port map (
            O => \N__31484\,
            I => \N__31481\
        );

    \I__5464\ : InMux
    port map (
            O => \N__31481\,
            I => \N__31476\
        );

    \I__5463\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31473\
        );

    \I__5462\ : CascadeMux
    port map (
            O => \N__31479\,
            I => \N__31469\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__31476\,
            I => \N__31464\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__31473\,
            I => \N__31461\
        );

    \I__5459\ : InMux
    port map (
            O => \N__31472\,
            I => \N__31458\
        );

    \I__5458\ : InMux
    port map (
            O => \N__31469\,
            I => \N__31455\
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__31468\,
            I => \N__31451\
        );

    \I__5456\ : CascadeMux
    port map (
            O => \N__31467\,
            I => \N__31447\
        );

    \I__5455\ : Span4Mux_h
    port map (
            O => \N__31464\,
            I => \N__31440\
        );

    \I__5454\ : Span4Mux_h
    port map (
            O => \N__31461\,
            I => \N__31440\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__31458\,
            I => \N__31440\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__31455\,
            I => \N__31437\
        );

    \I__5451\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31434\
        );

    \I__5450\ : InMux
    port map (
            O => \N__31451\,
            I => \N__31431\
        );

    \I__5449\ : InMux
    port map (
            O => \N__31450\,
            I => \N__31427\
        );

    \I__5448\ : InMux
    port map (
            O => \N__31447\,
            I => \N__31424\
        );

    \I__5447\ : Span4Mux_v
    port map (
            O => \N__31440\,
            I => \N__31421\
        );

    \I__5446\ : Span4Mux_v
    port map (
            O => \N__31437\,
            I => \N__31418\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__31434\,
            I => \N__31413\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__31431\,
            I => \N__31413\
        );

    \I__5443\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31410\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__31427\,
            I => un7_spon_15
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__31424\,
            I => un7_spon_15
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__31421\,
            I => un7_spon_15
        );

    \I__5439\ : Odrv4
    port map (
            O => \N__31418\,
            I => un7_spon_15
        );

    \I__5438\ : Odrv12
    port map (
            O => \N__31413\,
            I => un7_spon_15
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__31410\,
            I => un7_spon_15
        );

    \I__5436\ : CascadeMux
    port map (
            O => \N__31397\,
            I => \N__31394\
        );

    \I__5435\ : InMux
    port map (
            O => \N__31394\,
            I => \N__31390\
        );

    \I__5434\ : CascadeMux
    port map (
            O => \N__31393\,
            I => \N__31384\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__31390\,
            I => \N__31381\
        );

    \I__5432\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31378\
        );

    \I__5431\ : InMux
    port map (
            O => \N__31388\,
            I => \N__31373\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__31387\,
            I => \N__31370\
        );

    \I__5429\ : InMux
    port map (
            O => \N__31384\,
            I => \N__31367\
        );

    \I__5428\ : Span4Mux_v
    port map (
            O => \N__31381\,
            I => \N__31362\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__31378\,
            I => \N__31359\
        );

    \I__5426\ : InMux
    port map (
            O => \N__31377\,
            I => \N__31354\
        );

    \I__5425\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31354\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__31373\,
            I => \N__31351\
        );

    \I__5423\ : InMux
    port map (
            O => \N__31370\,
            I => \N__31348\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__31367\,
            I => \N__31345\
        );

    \I__5421\ : InMux
    port map (
            O => \N__31366\,
            I => \N__31342\
        );

    \I__5420\ : InMux
    port map (
            O => \N__31365\,
            I => \N__31339\
        );

    \I__5419\ : Span4Mux_h
    port map (
            O => \N__31362\,
            I => \N__31327\
        );

    \I__5418\ : Span4Mux_h
    port map (
            O => \N__31359\,
            I => \N__31327\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__31354\,
            I => \N__31327\
        );

    \I__5416\ : Span4Mux_v
    port map (
            O => \N__31351\,
            I => \N__31327\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__31348\,
            I => \N__31324\
        );

    \I__5414\ : Span4Mux_v
    port map (
            O => \N__31345\,
            I => \N__31319\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__31342\,
            I => \N__31319\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__31339\,
            I => \N__31316\
        );

    \I__5411\ : InMux
    port map (
            O => \N__31338\,
            I => \N__31313\
        );

    \I__5410\ : InMux
    port map (
            O => \N__31337\,
            I => \N__31310\
        );

    \I__5409\ : InMux
    port map (
            O => \N__31336\,
            I => \N__31307\
        );

    \I__5408\ : Span4Mux_v
    port map (
            O => \N__31327\,
            I => \N__31302\
        );

    \I__5407\ : Span4Mux_h
    port map (
            O => \N__31324\,
            I => \N__31302\
        );

    \I__5406\ : Span4Mux_v
    port map (
            O => \N__31319\,
            I => \N__31297\
        );

    \I__5405\ : Span4Mux_v
    port map (
            O => \N__31316\,
            I => \N__31297\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__31313\,
            I => un7_spon_16
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__31310\,
            I => un7_spon_16
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__31307\,
            I => un7_spon_16
        );

    \I__5401\ : Odrv4
    port map (
            O => \N__31302\,
            I => un7_spon_16
        );

    \I__5400\ : Odrv4
    port map (
            O => \N__31297\,
            I => un7_spon_16
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__31286\,
            I => \N__31280\
        );

    \I__5398\ : InMux
    port map (
            O => \N__31285\,
            I => \N__31277\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__31284\,
            I => \N__31273\
        );

    \I__5396\ : InMux
    port map (
            O => \N__31283\,
            I => \N__31270\
        );

    \I__5395\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31263\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__31277\,
            I => \N__31258\
        );

    \I__5393\ : InMux
    port map (
            O => \N__31276\,
            I => \N__31255\
        );

    \I__5392\ : InMux
    port map (
            O => \N__31273\,
            I => \N__31252\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__31270\,
            I => \N__31249\
        );

    \I__5390\ : InMux
    port map (
            O => \N__31269\,
            I => \N__31246\
        );

    \I__5389\ : CascadeMux
    port map (
            O => \N__31268\,
            I => \N__31243\
        );

    \I__5388\ : CascadeMux
    port map (
            O => \N__31267\,
            I => \N__31240\
        );

    \I__5387\ : InMux
    port map (
            O => \N__31266\,
            I => \N__31236\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__31263\,
            I => \N__31233\
        );

    \I__5385\ : InMux
    port map (
            O => \N__31262\,
            I => \N__31230\
        );

    \I__5384\ : InMux
    port map (
            O => \N__31261\,
            I => \N__31227\
        );

    \I__5383\ : Span4Mux_v
    port map (
            O => \N__31258\,
            I => \N__31222\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__31255\,
            I => \N__31222\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__31252\,
            I => \N__31219\
        );

    \I__5380\ : Span4Mux_v
    port map (
            O => \N__31249\,
            I => \N__31214\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__31246\,
            I => \N__31214\
        );

    \I__5378\ : InMux
    port map (
            O => \N__31243\,
            I => \N__31211\
        );

    \I__5377\ : InMux
    port map (
            O => \N__31240\,
            I => \N__31206\
        );

    \I__5376\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31206\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__31236\,
            I => \N__31203\
        );

    \I__5374\ : Span4Mux_v
    port map (
            O => \N__31233\,
            I => \N__31200\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__31230\,
            I => \N__31189\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__31227\,
            I => \N__31189\
        );

    \I__5371\ : Span4Mux_v
    port map (
            O => \N__31222\,
            I => \N__31189\
        );

    \I__5370\ : Span4Mux_h
    port map (
            O => \N__31219\,
            I => \N__31189\
        );

    \I__5369\ : Span4Mux_v
    port map (
            O => \N__31214\,
            I => \N__31189\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__31211\,
            I => un7_spon_17
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__31206\,
            I => un7_spon_17
        );

    \I__5366\ : Odrv12
    port map (
            O => \N__31203\,
            I => un7_spon_17
        );

    \I__5365\ : Odrv4
    port map (
            O => \N__31200\,
            I => un7_spon_17
        );

    \I__5364\ : Odrv4
    port map (
            O => \N__31189\,
            I => un7_spon_17
        );

    \I__5363\ : CascadeMux
    port map (
            O => \N__31178\,
            I => \N__31173\
        );

    \I__5362\ : CascadeMux
    port map (
            O => \N__31177\,
            I => \N__31170\
        );

    \I__5361\ : CascadeMux
    port map (
            O => \N__31176\,
            I => \N__31167\
        );

    \I__5360\ : InMux
    port map (
            O => \N__31173\,
            I => \N__31164\
        );

    \I__5359\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31157\
        );

    \I__5358\ : InMux
    port map (
            O => \N__31167\,
            I => \N__31154\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__31164\,
            I => \N__31151\
        );

    \I__5356\ : InMux
    port map (
            O => \N__31163\,
            I => \N__31145\
        );

    \I__5355\ : InMux
    port map (
            O => \N__31162\,
            I => \N__31142\
        );

    \I__5354\ : InMux
    port map (
            O => \N__31161\,
            I => \N__31137\
        );

    \I__5353\ : InMux
    port map (
            O => \N__31160\,
            I => \N__31137\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__31157\,
            I => \N__31134\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__31154\,
            I => \N__31131\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__31151\,
            I => \N__31128\
        );

    \I__5349\ : InMux
    port map (
            O => \N__31150\,
            I => \N__31125\
        );

    \I__5348\ : InMux
    port map (
            O => \N__31149\,
            I => \N__31120\
        );

    \I__5347\ : InMux
    port map (
            O => \N__31148\,
            I => \N__31117\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__31145\,
            I => \N__31114\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__31142\,
            I => \N__31111\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__31137\,
            I => \N__31108\
        );

    \I__5343\ : Span4Mux_h
    port map (
            O => \N__31134\,
            I => \N__31105\
        );

    \I__5342\ : Span4Mux_v
    port map (
            O => \N__31131\,
            I => \N__31098\
        );

    \I__5341\ : Span4Mux_h
    port map (
            O => \N__31128\,
            I => \N__31098\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__31125\,
            I => \N__31098\
        );

    \I__5339\ : InMux
    port map (
            O => \N__31124\,
            I => \N__31095\
        );

    \I__5338\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31092\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__31120\,
            I => \N__31089\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__31117\,
            I => \N__31076\
        );

    \I__5335\ : Span4Mux_h
    port map (
            O => \N__31114\,
            I => \N__31076\
        );

    \I__5334\ : Span4Mux_h
    port map (
            O => \N__31111\,
            I => \N__31076\
        );

    \I__5333\ : Span4Mux_v
    port map (
            O => \N__31108\,
            I => \N__31076\
        );

    \I__5332\ : Span4Mux_v
    port map (
            O => \N__31105\,
            I => \N__31076\
        );

    \I__5331\ : Span4Mux_v
    port map (
            O => \N__31098\,
            I => \N__31076\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__31095\,
            I => un7_spon_18
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__31092\,
            I => un7_spon_18
        );

    \I__5328\ : Odrv12
    port map (
            O => \N__31089\,
            I => un7_spon_18
        );

    \I__5327\ : Odrv4
    port map (
            O => \N__31076\,
            I => un7_spon_18
        );

    \I__5326\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31064\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__31064\,
            I => \sEEPonPoffZ0Z_4\
        );

    \I__5324\ : CascadeMux
    port map (
            O => \N__31061\,
            I => \N__31056\
        );

    \I__5323\ : CascadeMux
    port map (
            O => \N__31060\,
            I => \N__31053\
        );

    \I__5322\ : InMux
    port map (
            O => \N__31059\,
            I => \N__31049\
        );

    \I__5321\ : InMux
    port map (
            O => \N__31056\,
            I => \N__31045\
        );

    \I__5320\ : InMux
    port map (
            O => \N__31053\,
            I => \N__31042\
        );

    \I__5319\ : CascadeMux
    port map (
            O => \N__31052\,
            I => \N__31039\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__31049\,
            I => \N__31035\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__31048\,
            I => \N__31030\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__31045\,
            I => \N__31026\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__31042\,
            I => \N__31023\
        );

    \I__5314\ : InMux
    port map (
            O => \N__31039\,
            I => \N__31020\
        );

    \I__5313\ : CascadeMux
    port map (
            O => \N__31038\,
            I => \N__31017\
        );

    \I__5312\ : Span4Mux_v
    port map (
            O => \N__31035\,
            I => \N__31013\
        );

    \I__5311\ : InMux
    port map (
            O => \N__31034\,
            I => \N__31008\
        );

    \I__5310\ : InMux
    port map (
            O => \N__31033\,
            I => \N__31008\
        );

    \I__5309\ : InMux
    port map (
            O => \N__31030\,
            I => \N__31005\
        );

    \I__5308\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31002\
        );

    \I__5307\ : Span4Mux_h
    port map (
            O => \N__31026\,
            I => \N__30996\
        );

    \I__5306\ : Span4Mux_v
    port map (
            O => \N__31023\,
            I => \N__30991\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__31020\,
            I => \N__30991\
        );

    \I__5304\ : InMux
    port map (
            O => \N__31017\,
            I => \N__30988\
        );

    \I__5303\ : CascadeMux
    port map (
            O => \N__31016\,
            I => \N__30985\
        );

    \I__5302\ : Span4Mux_v
    port map (
            O => \N__31013\,
            I => \N__30975\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__31008\,
            I => \N__30975\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__31005\,
            I => \N__30975\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__31002\,
            I => \N__30975\
        );

    \I__5298\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30972\
        );

    \I__5297\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30969\
        );

    \I__5296\ : InMux
    port map (
            O => \N__30999\,
            I => \N__30966\
        );

    \I__5295\ : Span4Mux_v
    port map (
            O => \N__30996\,
            I => \N__30959\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__30991\,
            I => \N__30959\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__30988\,
            I => \N__30959\
        );

    \I__5292\ : InMux
    port map (
            O => \N__30985\,
            I => \N__30956\
        );

    \I__5291\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30952\
        );

    \I__5290\ : Span4Mux_v
    port map (
            O => \N__30975\,
            I => \N__30949\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__30972\,
            I => \N__30946\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__30969\,
            I => \N__30939\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__30966\,
            I => \N__30939\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__30959\,
            I => \N__30939\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__30956\,
            I => \N__30936\
        );

    \I__5284\ : InMux
    port map (
            O => \N__30955\,
            I => \N__30933\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__30952\,
            I => un7_spon_4
        );

    \I__5282\ : Odrv4
    port map (
            O => \N__30949\,
            I => un7_spon_4
        );

    \I__5281\ : Odrv12
    port map (
            O => \N__30946\,
            I => un7_spon_4
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__30939\,
            I => un7_spon_4
        );

    \I__5279\ : Odrv12
    port map (
            O => \N__30936\,
            I => un7_spon_4
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__30933\,
            I => un7_spon_4
        );

    \I__5277\ : InMux
    port map (
            O => \N__30920\,
            I => \N__30917\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__30917\,
            I => \sEEPonPoff_i_4\
        );

    \I__5275\ : InMux
    port map (
            O => \N__30914\,
            I => \N__30911\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__30911\,
            I => \sEEPonPoffZ0Z_5\
        );

    \I__5273\ : CascadeMux
    port map (
            O => \N__30908\,
            I => \N__30904\
        );

    \I__5272\ : CascadeMux
    port map (
            O => \N__30907\,
            I => \N__30901\
        );

    \I__5271\ : InMux
    port map (
            O => \N__30904\,
            I => \N__30895\
        );

    \I__5270\ : InMux
    port map (
            O => \N__30901\,
            I => \N__30892\
        );

    \I__5269\ : CascadeMux
    port map (
            O => \N__30900\,
            I => \N__30889\
        );

    \I__5268\ : CascadeMux
    port map (
            O => \N__30899\,
            I => \N__30885\
        );

    \I__5267\ : InMux
    port map (
            O => \N__30898\,
            I => \N__30882\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__30895\,
            I => \N__30876\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__30892\,
            I => \N__30873\
        );

    \I__5264\ : InMux
    port map (
            O => \N__30889\,
            I => \N__30870\
        );

    \I__5263\ : InMux
    port map (
            O => \N__30888\,
            I => \N__30867\
        );

    \I__5262\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30864\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__30882\,
            I => \N__30860\
        );

    \I__5260\ : InMux
    port map (
            O => \N__30881\,
            I => \N__30857\
        );

    \I__5259\ : InMux
    port map (
            O => \N__30880\,
            I => \N__30852\
        );

    \I__5258\ : InMux
    port map (
            O => \N__30879\,
            I => \N__30852\
        );

    \I__5257\ : Span4Mux_h
    port map (
            O => \N__30876\,
            I => \N__30845\
        );

    \I__5256\ : Span4Mux_h
    port map (
            O => \N__30873\,
            I => \N__30845\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__30870\,
            I => \N__30845\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__30867\,
            I => \N__30842\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__30864\,
            I => \N__30839\
        );

    \I__5252\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30835\
        );

    \I__5251\ : Span4Mux_h
    port map (
            O => \N__30860\,
            I => \N__30832\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__30857\,
            I => \N__30829\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__30852\,
            I => \N__30824\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__30845\,
            I => \N__30824\
        );

    \I__5247\ : Span4Mux_h
    port map (
            O => \N__30842\,
            I => \N__30819\
        );

    \I__5246\ : Span4Mux_v
    port map (
            O => \N__30839\,
            I => \N__30819\
        );

    \I__5245\ : InMux
    port map (
            O => \N__30838\,
            I => \N__30816\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__30835\,
            I => un7_spon_5
        );

    \I__5243\ : Odrv4
    port map (
            O => \N__30832\,
            I => un7_spon_5
        );

    \I__5242\ : Odrv4
    port map (
            O => \N__30829\,
            I => un7_spon_5
        );

    \I__5241\ : Odrv4
    port map (
            O => \N__30824\,
            I => un7_spon_5
        );

    \I__5240\ : Odrv4
    port map (
            O => \N__30819\,
            I => un7_spon_5
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__30816\,
            I => un7_spon_5
        );

    \I__5238\ : InMux
    port map (
            O => \N__30803\,
            I => \N__30800\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__30800\,
            I => \sEEPonPoff_i_5\
        );

    \I__5236\ : InMux
    port map (
            O => \N__30797\,
            I => \N__30794\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__30794\,
            I => \sEEPonPoffZ0Z_6\
        );

    \I__5234\ : CascadeMux
    port map (
            O => \N__30791\,
            I => \N__30787\
        );

    \I__5233\ : CascadeMux
    port map (
            O => \N__30790\,
            I => \N__30782\
        );

    \I__5232\ : InMux
    port map (
            O => \N__30787\,
            I => \N__30778\
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__30786\,
            I => \N__30775\
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__30785\,
            I => \N__30770\
        );

    \I__5229\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30766\
        );

    \I__5228\ : InMux
    port map (
            O => \N__30781\,
            I => \N__30763\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__30778\,
            I => \N__30759\
        );

    \I__5226\ : InMux
    port map (
            O => \N__30775\,
            I => \N__30756\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__30774\,
            I => \N__30753\
        );

    \I__5224\ : InMux
    port map (
            O => \N__30773\,
            I => \N__30747\
        );

    \I__5223\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30747\
        );

    \I__5222\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30744\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__30766\,
            I => \N__30739\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__30763\,
            I => \N__30739\
        );

    \I__5219\ : InMux
    port map (
            O => \N__30762\,
            I => \N__30736\
        );

    \I__5218\ : Span4Mux_h
    port map (
            O => \N__30759\,
            I => \N__30731\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__30756\,
            I => \N__30731\
        );

    \I__5216\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30728\
        );

    \I__5215\ : InMux
    port map (
            O => \N__30752\,
            I => \N__30724\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__30747\,
            I => \N__30719\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__30744\,
            I => \N__30719\
        );

    \I__5212\ : Span12Mux_v
    port map (
            O => \N__30739\,
            I => \N__30714\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__30736\,
            I => \N__30714\
        );

    \I__5210\ : Span4Mux_v
    port map (
            O => \N__30731\,
            I => \N__30711\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__30728\,
            I => \N__30708\
        );

    \I__5208\ : InMux
    port map (
            O => \N__30727\,
            I => \N__30705\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__30724\,
            I => un7_spon_6
        );

    \I__5206\ : Odrv4
    port map (
            O => \N__30719\,
            I => un7_spon_6
        );

    \I__5205\ : Odrv12
    port map (
            O => \N__30714\,
            I => un7_spon_6
        );

    \I__5204\ : Odrv4
    port map (
            O => \N__30711\,
            I => un7_spon_6
        );

    \I__5203\ : Odrv12
    port map (
            O => \N__30708\,
            I => un7_spon_6
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__30705\,
            I => un7_spon_6
        );

    \I__5201\ : InMux
    port map (
            O => \N__30692\,
            I => \N__30689\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__30689\,
            I => \sEEPonPoff_i_6\
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__30686\,
            I => \N__30683\
        );

    \I__5198\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30679\
        );

    \I__5197\ : CascadeMux
    port map (
            O => \N__30682\,
            I => \N__30676\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__30679\,
            I => \N__30671\
        );

    \I__5195\ : InMux
    port map (
            O => \N__30676\,
            I => \N__30668\
        );

    \I__5194\ : InMux
    port map (
            O => \N__30675\,
            I => \N__30664\
        );

    \I__5193\ : InMux
    port map (
            O => \N__30674\,
            I => \N__30661\
        );

    \I__5192\ : Span4Mux_h
    port map (
            O => \N__30671\,
            I => \N__30656\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__30668\,
            I => \N__30656\
        );

    \I__5190\ : InMux
    port map (
            O => \N__30667\,
            I => \N__30653\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__30664\,
            I => \N__30644\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__30661\,
            I => \N__30644\
        );

    \I__5187\ : Span4Mux_h
    port map (
            O => \N__30656\,
            I => \N__30641\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__30653\,
            I => \N__30638\
        );

    \I__5185\ : InMux
    port map (
            O => \N__30652\,
            I => \N__30635\
        );

    \I__5184\ : InMux
    port map (
            O => \N__30651\,
            I => \N__30631\
        );

    \I__5183\ : InMux
    port map (
            O => \N__30650\,
            I => \N__30628\
        );

    \I__5182\ : InMux
    port map (
            O => \N__30649\,
            I => \N__30624\
        );

    \I__5181\ : Span4Mux_h
    port map (
            O => \N__30644\,
            I => \N__30621\
        );

    \I__5180\ : Span4Mux_v
    port map (
            O => \N__30641\,
            I => \N__30616\
        );

    \I__5179\ : Span4Mux_h
    port map (
            O => \N__30638\,
            I => \N__30616\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__30635\,
            I => \N__30613\
        );

    \I__5177\ : InMux
    port map (
            O => \N__30634\,
            I => \N__30610\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__30631\,
            I => \N__30605\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__30628\,
            I => \N__30605\
        );

    \I__5174\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30602\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__30624\,
            I => un7_spon_7
        );

    \I__5172\ : Odrv4
    port map (
            O => \N__30621\,
            I => un7_spon_7
        );

    \I__5171\ : Odrv4
    port map (
            O => \N__30616\,
            I => un7_spon_7
        );

    \I__5170\ : Odrv12
    port map (
            O => \N__30613\,
            I => un7_spon_7
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__30610\,
            I => un7_spon_7
        );

    \I__5168\ : Odrv12
    port map (
            O => \N__30605\,
            I => un7_spon_7
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__30602\,
            I => un7_spon_7
        );

    \I__5166\ : InMux
    port map (
            O => \N__30587\,
            I => \N__30584\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__30584\,
            I => \sEEPonPoffZ0Z_7\
        );

    \I__5164\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30578\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__30578\,
            I => \sEEPonPoff_i_7\
        );

    \I__5162\ : CascadeMux
    port map (
            O => \N__30575\,
            I => \N__30572\
        );

    \I__5161\ : InMux
    port map (
            O => \N__30572\,
            I => \N__30567\
        );

    \I__5160\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30564\
        );

    \I__5159\ : CascadeMux
    port map (
            O => \N__30570\,
            I => \N__30559\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__30567\,
            I => \N__30556\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__30564\,
            I => \N__30552\
        );

    \I__5156\ : InMux
    port map (
            O => \N__30563\,
            I => \N__30548\
        );

    \I__5155\ : CascadeMux
    port map (
            O => \N__30562\,
            I => \N__30545\
        );

    \I__5154\ : InMux
    port map (
            O => \N__30559\,
            I => \N__30542\
        );

    \I__5153\ : Span4Mux_v
    port map (
            O => \N__30556\,
            I => \N__30538\
        );

    \I__5152\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30535\
        );

    \I__5151\ : Span4Mux_v
    port map (
            O => \N__30552\,
            I => \N__30530\
        );

    \I__5150\ : InMux
    port map (
            O => \N__30551\,
            I => \N__30527\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__30548\,
            I => \N__30524\
        );

    \I__5148\ : InMux
    port map (
            O => \N__30545\,
            I => \N__30521\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__30542\,
            I => \N__30518\
        );

    \I__5146\ : InMux
    port map (
            O => \N__30541\,
            I => \N__30514\
        );

    \I__5145\ : Span4Mux_v
    port map (
            O => \N__30538\,
            I => \N__30509\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__30535\,
            I => \N__30509\
        );

    \I__5143\ : InMux
    port map (
            O => \N__30534\,
            I => \N__30504\
        );

    \I__5142\ : InMux
    port map (
            O => \N__30533\,
            I => \N__30504\
        );

    \I__5141\ : Span4Mux_v
    port map (
            O => \N__30530\,
            I => \N__30499\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__30527\,
            I => \N__30499\
        );

    \I__5139\ : Span4Mux_h
    port map (
            O => \N__30524\,
            I => \N__30496\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__30521\,
            I => \N__30493\
        );

    \I__5137\ : Span4Mux_h
    port map (
            O => \N__30518\,
            I => \N__30490\
        );

    \I__5136\ : InMux
    port map (
            O => \N__30517\,
            I => \N__30487\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__30514\,
            I => un7_spon_8
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__30509\,
            I => un7_spon_8
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__30504\,
            I => un7_spon_8
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__30499\,
            I => un7_spon_8
        );

    \I__5131\ : Odrv4
    port map (
            O => \N__30496\,
            I => un7_spon_8
        );

    \I__5130\ : Odrv12
    port map (
            O => \N__30493\,
            I => un7_spon_8
        );

    \I__5129\ : Odrv4
    port map (
            O => \N__30490\,
            I => un7_spon_8
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__30487\,
            I => un7_spon_8
        );

    \I__5127\ : CascadeMux
    port map (
            O => \N__30470\,
            I => \N__30467\
        );

    \I__5126\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30462\
        );

    \I__5125\ : InMux
    port map (
            O => \N__30466\,
            I => \N__30459\
        );

    \I__5124\ : CascadeMux
    port map (
            O => \N__30465\,
            I => \N__30453\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__30462\,
            I => \N__30450\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__30459\,
            I => \N__30447\
        );

    \I__5121\ : InMux
    port map (
            O => \N__30458\,
            I => \N__30442\
        );

    \I__5120\ : InMux
    port map (
            O => \N__30457\,
            I => \N__30439\
        );

    \I__5119\ : CascadeMux
    port map (
            O => \N__30456\,
            I => \N__30436\
        );

    \I__5118\ : InMux
    port map (
            O => \N__30453\,
            I => \N__30433\
        );

    \I__5117\ : Span4Mux_v
    port map (
            O => \N__30450\,
            I => \N__30430\
        );

    \I__5116\ : Span4Mux_v
    port map (
            O => \N__30447\,
            I => \N__30427\
        );

    \I__5115\ : CascadeMux
    port map (
            O => \N__30446\,
            I => \N__30423\
        );

    \I__5114\ : InMux
    port map (
            O => \N__30445\,
            I => \N__30419\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__30442\,
            I => \N__30414\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__30439\,
            I => \N__30414\
        );

    \I__5111\ : InMux
    port map (
            O => \N__30436\,
            I => \N__30411\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__30433\,
            I => \N__30408\
        );

    \I__5109\ : Span4Mux_v
    port map (
            O => \N__30430\,
            I => \N__30402\
        );

    \I__5108\ : Span4Mux_v
    port map (
            O => \N__30427\,
            I => \N__30402\
        );

    \I__5107\ : InMux
    port map (
            O => \N__30426\,
            I => \N__30399\
        );

    \I__5106\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30394\
        );

    \I__5105\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30394\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__30419\,
            I => \N__30391\
        );

    \I__5103\ : Span4Mux_h
    port map (
            O => \N__30414\,
            I => \N__30388\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__30411\,
            I => \N__30385\
        );

    \I__5101\ : Span4Mux_h
    port map (
            O => \N__30408\,
            I => \N__30382\
        );

    \I__5100\ : InMux
    port map (
            O => \N__30407\,
            I => \N__30379\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__30402\,
            I => un7_spon_9
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__30399\,
            I => un7_spon_9
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__30394\,
            I => un7_spon_9
        );

    \I__5096\ : Odrv4
    port map (
            O => \N__30391\,
            I => un7_spon_9
        );

    \I__5095\ : Odrv4
    port map (
            O => \N__30388\,
            I => un7_spon_9
        );

    \I__5094\ : Odrv12
    port map (
            O => \N__30385\,
            I => un7_spon_9
        );

    \I__5093\ : Odrv4
    port map (
            O => \N__30382\,
            I => un7_spon_9
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__30379\,
            I => un7_spon_9
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__30362\,
            I => \N__30357\
        );

    \I__5090\ : CascadeMux
    port map (
            O => \N__30361\,
            I => \N__30354\
        );

    \I__5089\ : InMux
    port map (
            O => \N__30360\,
            I => \N__30350\
        );

    \I__5088\ : InMux
    port map (
            O => \N__30357\,
            I => \N__30347\
        );

    \I__5087\ : InMux
    port map (
            O => \N__30354\,
            I => \N__30342\
        );

    \I__5086\ : CascadeMux
    port map (
            O => \N__30353\,
            I => \N__30338\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__30350\,
            I => \N__30334\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__30347\,
            I => \N__30331\
        );

    \I__5083\ : InMux
    port map (
            O => \N__30346\,
            I => \N__30328\
        );

    \I__5082\ : InMux
    port map (
            O => \N__30345\,
            I => \N__30325\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__30342\,
            I => \N__30322\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__30341\,
            I => \N__30319\
        );

    \I__5079\ : InMux
    port map (
            O => \N__30338\,
            I => \N__30316\
        );

    \I__5078\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30311\
        );

    \I__5077\ : Span4Mux_v
    port map (
            O => \N__30334\,
            I => \N__30308\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__30331\,
            I => \N__30303\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__30328\,
            I => \N__30303\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__30325\,
            I => \N__30300\
        );

    \I__5073\ : Span4Mux_v
    port map (
            O => \N__30322\,
            I => \N__30297\
        );

    \I__5072\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30294\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__30316\,
            I => \N__30291\
        );

    \I__5070\ : InMux
    port map (
            O => \N__30315\,
            I => \N__30287\
        );

    \I__5069\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30284\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__30311\,
            I => \N__30281\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__30308\,
            I => \N__30272\
        );

    \I__5066\ : Span4Mux_v
    port map (
            O => \N__30303\,
            I => \N__30272\
        );

    \I__5065\ : Span4Mux_h
    port map (
            O => \N__30300\,
            I => \N__30272\
        );

    \I__5064\ : Span4Mux_h
    port map (
            O => \N__30297\,
            I => \N__30272\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__30294\,
            I => \N__30269\
        );

    \I__5062\ : Span4Mux_h
    port map (
            O => \N__30291\,
            I => \N__30266\
        );

    \I__5061\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30263\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__30287\,
            I => un7_spon_10
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__30284\,
            I => un7_spon_10
        );

    \I__5058\ : Odrv4
    port map (
            O => \N__30281\,
            I => un7_spon_10
        );

    \I__5057\ : Odrv4
    port map (
            O => \N__30272\,
            I => un7_spon_10
        );

    \I__5056\ : Odrv12
    port map (
            O => \N__30269\,
            I => un7_spon_10
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__30266\,
            I => un7_spon_10
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__30263\,
            I => un7_spon_10
        );

    \I__5053\ : InMux
    port map (
            O => \N__30248\,
            I => \N__30245\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__30245\,
            I => \sEEPonPoffZ0Z_0\
        );

    \I__5051\ : CascadeMux
    port map (
            O => \N__30242\,
            I => \N__30238\
        );

    \I__5050\ : InMux
    port map (
            O => \N__30241\,
            I => \N__30234\
        );

    \I__5049\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30230\
        );

    \I__5048\ : CascadeMux
    port map (
            O => \N__30237\,
            I => \N__30226\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__30234\,
            I => \N__30223\
        );

    \I__5046\ : InMux
    port map (
            O => \N__30233\,
            I => \N__30220\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__30230\,
            I => \N__30217\
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__30229\,
            I => \N__30213\
        );

    \I__5043\ : InMux
    port map (
            O => \N__30226\,
            I => \N__30210\
        );

    \I__5042\ : Span4Mux_v
    port map (
            O => \N__30223\,
            I => \N__30207\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__30220\,
            I => \N__30201\
        );

    \I__5040\ : Span4Mux_v
    port map (
            O => \N__30217\,
            I => \N__30198\
        );

    \I__5039\ : InMux
    port map (
            O => \N__30216\,
            I => \N__30195\
        );

    \I__5038\ : InMux
    port map (
            O => \N__30213\,
            I => \N__30192\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__30210\,
            I => \N__30189\
        );

    \I__5036\ : Span4Mux_v
    port map (
            O => \N__30207\,
            I => \N__30185\
        );

    \I__5035\ : InMux
    port map (
            O => \N__30206\,
            I => \N__30182\
        );

    \I__5034\ : InMux
    port map (
            O => \N__30205\,
            I => \N__30177\
        );

    \I__5033\ : InMux
    port map (
            O => \N__30204\,
            I => \N__30177\
        );

    \I__5032\ : Span4Mux_h
    port map (
            O => \N__30201\,
            I => \N__30174\
        );

    \I__5031\ : Span4Mux_v
    port map (
            O => \N__30198\,
            I => \N__30169\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__30195\,
            I => \N__30169\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__30192\,
            I => \N__30166\
        );

    \I__5028\ : Span4Mux_h
    port map (
            O => \N__30189\,
            I => \N__30163\
        );

    \I__5027\ : InMux
    port map (
            O => \N__30188\,
            I => \N__30160\
        );

    \I__5026\ : Odrv4
    port map (
            O => \N__30185\,
            I => un7_spon_0
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__30182\,
            I => un7_spon_0
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__30177\,
            I => un7_spon_0
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__30174\,
            I => un7_spon_0
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__30169\,
            I => un7_spon_0
        );

    \I__5021\ : Odrv12
    port map (
            O => \N__30166\,
            I => un7_spon_0
        );

    \I__5020\ : Odrv4
    port map (
            O => \N__30163\,
            I => un7_spon_0
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__30160\,
            I => un7_spon_0
        );

    \I__5018\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30140\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__30140\,
            I => \sEEPonPoff_i_0\
        );

    \I__5016\ : CascadeMux
    port map (
            O => \N__30137\,
            I => \N__30134\
        );

    \I__5015\ : InMux
    port map (
            O => \N__30134\,
            I => \N__30131\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__30131\,
            I => \N__30127\
        );

    \I__5013\ : CascadeMux
    port map (
            O => \N__30130\,
            I => \N__30124\
        );

    \I__5012\ : Span4Mux_v
    port map (
            O => \N__30127\,
            I => \N__30121\
        );

    \I__5011\ : InMux
    port map (
            O => \N__30124\,
            I => \N__30118\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__30121\,
            I => \N__30112\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__30118\,
            I => \N__30112\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__30117\,
            I => \N__30106\
        );

    \I__5007\ : Span4Mux_v
    port map (
            O => \N__30112\,
            I => \N__30103\
        );

    \I__5006\ : InMux
    port map (
            O => \N__30111\,
            I => \N__30100\
        );

    \I__5005\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30097\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__30109\,
            I => \N__30093\
        );

    \I__5003\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30090\
        );

    \I__5002\ : Span4Mux_h
    port map (
            O => \N__30103\,
            I => \N__30082\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__30100\,
            I => \N__30082\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__30097\,
            I => \N__30082\
        );

    \I__4999\ : InMux
    port map (
            O => \N__30096\,
            I => \N__30077\
        );

    \I__4998\ : InMux
    port map (
            O => \N__30093\,
            I => \N__30074\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__30090\,
            I => \N__30071\
        );

    \I__4996\ : InMux
    port map (
            O => \N__30089\,
            I => \N__30067\
        );

    \I__4995\ : Span4Mux_v
    port map (
            O => \N__30082\,
            I => \N__30064\
        );

    \I__4994\ : InMux
    port map (
            O => \N__30081\,
            I => \N__30059\
        );

    \I__4993\ : InMux
    port map (
            O => \N__30080\,
            I => \N__30059\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__30077\,
            I => \N__30056\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__30074\,
            I => \N__30053\
        );

    \I__4990\ : Span4Mux_h
    port map (
            O => \N__30071\,
            I => \N__30050\
        );

    \I__4989\ : InMux
    port map (
            O => \N__30070\,
            I => \N__30047\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__30067\,
            I => un7_spon_1
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__30064\,
            I => un7_spon_1
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__30059\,
            I => un7_spon_1
        );

    \I__4985\ : Odrv12
    port map (
            O => \N__30056\,
            I => un7_spon_1
        );

    \I__4984\ : Odrv12
    port map (
            O => \N__30053\,
            I => un7_spon_1
        );

    \I__4983\ : Odrv4
    port map (
            O => \N__30050\,
            I => un7_spon_1
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__30047\,
            I => un7_spon_1
        );

    \I__4981\ : InMux
    port map (
            O => \N__30032\,
            I => \N__30029\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__30029\,
            I => \sEEPonPoffZ0Z_1\
        );

    \I__4979\ : InMux
    port map (
            O => \N__30026\,
            I => \N__30023\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__30023\,
            I => \sEEPonPoff_i_1\
        );

    \I__4977\ : InMux
    port map (
            O => \N__30020\,
            I => \N__30017\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__30017\,
            I => \sEEPonPoffZ0Z_2\
        );

    \I__4975\ : CascadeMux
    port map (
            O => \N__30014\,
            I => \N__30010\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__30013\,
            I => \N__30007\
        );

    \I__4973\ : InMux
    port map (
            O => \N__30010\,
            I => \N__30002\
        );

    \I__4972\ : InMux
    port map (
            O => \N__30007\,
            I => \N__29999\
        );

    \I__4971\ : CascadeMux
    port map (
            O => \N__30006\,
            I => \N__29993\
        );

    \I__4970\ : InMux
    port map (
            O => \N__30005\,
            I => \N__29990\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__30002\,
            I => \N__29987\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__29999\,
            I => \N__29984\
        );

    \I__4967\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29980\
        );

    \I__4966\ : CascadeMux
    port map (
            O => \N__29997\,
            I => \N__29977\
        );

    \I__4965\ : CascadeMux
    port map (
            O => \N__29996\,
            I => \N__29974\
        );

    \I__4964\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29971\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__29990\,
            I => \N__29966\
        );

    \I__4962\ : Span4Mux_h
    port map (
            O => \N__29987\,
            I => \N__29961\
        );

    \I__4961\ : Span4Mux_h
    port map (
            O => \N__29984\,
            I => \N__29961\
        );

    \I__4960\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29958\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__29980\,
            I => \N__29955\
        );

    \I__4958\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29952\
        );

    \I__4957\ : InMux
    port map (
            O => \N__29974\,
            I => \N__29949\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__29971\,
            I => \N__29946\
        );

    \I__4955\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29942\
        );

    \I__4954\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29939\
        );

    \I__4953\ : Span4Mux_v
    port map (
            O => \N__29966\,
            I => \N__29936\
        );

    \I__4952\ : Span4Mux_v
    port map (
            O => \N__29961\,
            I => \N__29931\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__29958\,
            I => \N__29931\
        );

    \I__4950\ : Span4Mux_h
    port map (
            O => \N__29955\,
            I => \N__29928\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__29952\,
            I => \N__29925\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__29949\,
            I => \N__29922\
        );

    \I__4947\ : Span4Mux_h
    port map (
            O => \N__29946\,
            I => \N__29919\
        );

    \I__4946\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29916\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__29942\,
            I => un7_spon_2
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__29939\,
            I => un7_spon_2
        );

    \I__4943\ : Odrv4
    port map (
            O => \N__29936\,
            I => un7_spon_2
        );

    \I__4942\ : Odrv4
    port map (
            O => \N__29931\,
            I => un7_spon_2
        );

    \I__4941\ : Odrv4
    port map (
            O => \N__29928\,
            I => un7_spon_2
        );

    \I__4940\ : Odrv12
    port map (
            O => \N__29925\,
            I => un7_spon_2
        );

    \I__4939\ : Odrv12
    port map (
            O => \N__29922\,
            I => un7_spon_2
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__29919\,
            I => un7_spon_2
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__29916\,
            I => un7_spon_2
        );

    \I__4936\ : InMux
    port map (
            O => \N__29897\,
            I => \N__29894\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__29894\,
            I => \sEEPonPoff_i_2\
        );

    \I__4934\ : InMux
    port map (
            O => \N__29891\,
            I => \N__29888\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__29888\,
            I => \sEEPonPoffZ0Z_3\
        );

    \I__4932\ : CascadeMux
    port map (
            O => \N__29885\,
            I => \N__29881\
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__29884\,
            I => \N__29878\
        );

    \I__4930\ : InMux
    port map (
            O => \N__29881\,
            I => \N__29874\
        );

    \I__4929\ : InMux
    port map (
            O => \N__29878\,
            I => \N__29868\
        );

    \I__4928\ : CascadeMux
    port map (
            O => \N__29877\,
            I => \N__29864\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__29874\,
            I => \N__29861\
        );

    \I__4926\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29858\
        );

    \I__4925\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29855\
        );

    \I__4924\ : InMux
    port map (
            O => \N__29871\,
            I => \N__29852\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__29868\,
            I => \N__29848\
        );

    \I__4922\ : InMux
    port map (
            O => \N__29867\,
            I => \N__29845\
        );

    \I__4921\ : InMux
    port map (
            O => \N__29864\,
            I => \N__29842\
        );

    \I__4920\ : Span4Mux_v
    port map (
            O => \N__29861\,
            I => \N__29833\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__29858\,
            I => \N__29833\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__29855\,
            I => \N__29833\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__29852\,
            I => \N__29830\
        );

    \I__4916\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29827\
        );

    \I__4915\ : Span4Mux_h
    port map (
            O => \N__29848\,
            I => \N__29822\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__29845\,
            I => \N__29822\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__29842\,
            I => \N__29819\
        );

    \I__4912\ : InMux
    port map (
            O => \N__29841\,
            I => \N__29815\
        );

    \I__4911\ : InMux
    port map (
            O => \N__29840\,
            I => \N__29812\
        );

    \I__4910\ : Span4Mux_v
    port map (
            O => \N__29833\,
            I => \N__29807\
        );

    \I__4909\ : Span4Mux_h
    port map (
            O => \N__29830\,
            I => \N__29807\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__29827\,
            I => \N__29802\
        );

    \I__4907\ : Span4Mux_v
    port map (
            O => \N__29822\,
            I => \N__29802\
        );

    \I__4906\ : Span4Mux_h
    port map (
            O => \N__29819\,
            I => \N__29799\
        );

    \I__4905\ : InMux
    port map (
            O => \N__29818\,
            I => \N__29796\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__29815\,
            I => un7_spon_3
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__29812\,
            I => un7_spon_3
        );

    \I__4902\ : Odrv4
    port map (
            O => \N__29807\,
            I => un7_spon_3
        );

    \I__4901\ : Odrv4
    port map (
            O => \N__29802\,
            I => un7_spon_3
        );

    \I__4900\ : Odrv4
    port map (
            O => \N__29799\,
            I => un7_spon_3
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__29796\,
            I => un7_spon_3
        );

    \I__4898\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29780\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__29780\,
            I => \sEEPonPoff_i_3\
        );

    \I__4896\ : InMux
    port map (
            O => \N__29777\,
            I => \N__29774\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__29774\,
            I => \N__29771\
        );

    \I__4894\ : Odrv4
    port map (
            O => \N__29771\,
            I => \sDAC_mem_27Z0Z_2\
        );

    \I__4893\ : InMux
    port map (
            O => \N__29768\,
            I => \N__29765\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__29765\,
            I => \N__29762\
        );

    \I__4891\ : Span4Mux_h
    port map (
            O => \N__29762\,
            I => \N__29759\
        );

    \I__4890\ : Odrv4
    port map (
            O => \N__29759\,
            I => \sDAC_mem_27Z0Z_4\
        );

    \I__4889\ : InMux
    port map (
            O => \N__29756\,
            I => \N__29753\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__29753\,
            I => \N__29750\
        );

    \I__4887\ : Odrv4
    port map (
            O => \N__29750\,
            I => \sDAC_mem_27Z0Z_5\
        );

    \I__4886\ : InMux
    port map (
            O => \N__29747\,
            I => \N__29744\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__29744\,
            I => \N__29741\
        );

    \I__4884\ : Span4Mux_v
    port map (
            O => \N__29741\,
            I => \N__29738\
        );

    \I__4883\ : Odrv4
    port map (
            O => \N__29738\,
            I => \sDAC_mem_27Z0Z_6\
        );

    \I__4882\ : InMux
    port map (
            O => \N__29735\,
            I => \N__29732\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__29732\,
            I => \N__29729\
        );

    \I__4880\ : Odrv4
    port map (
            O => \N__29729\,
            I => \sDAC_mem_27Z0Z_7\
        );

    \I__4879\ : CEMux
    port map (
            O => \N__29726\,
            I => \N__29723\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__29723\,
            I => \N__29720\
        );

    \I__4877\ : Span12Mux_h
    port map (
            O => \N__29720\,
            I => \N__29717\
        );

    \I__4876\ : Odrv12
    port map (
            O => \N__29717\,
            I => \sDAC_mem_27_1_sqmuxa\
        );

    \I__4875\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29711\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__29711\,
            I => \sDAC_mem_28Z0Z_6\
        );

    \I__4873\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29705\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__29705\,
            I => \N__29702\
        );

    \I__4871\ : Odrv12
    port map (
            O => \N__29702\,
            I => \sDAC_mem_31Z0Z_0\
        );

    \I__4870\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29696\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__29696\,
            I => \N__29693\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__29693\,
            I => \N__29690\
        );

    \I__4867\ : Span4Mux_h
    port map (
            O => \N__29690\,
            I => \N__29687\
        );

    \I__4866\ : Odrv4
    port map (
            O => \N__29687\,
            I => \sDAC_mem_30Z0Z_0\
        );

    \I__4865\ : InMux
    port map (
            O => \N__29684\,
            I => \N__29681\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__29681\,
            I => \N__29678\
        );

    \I__4863\ : Odrv12
    port map (
            O => \N__29678\,
            I => \sDAC_mem_31Z0Z_3\
        );

    \I__4862\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29672\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__29672\,
            I => \N__29669\
        );

    \I__4860\ : Span12Mux_h
    port map (
            O => \N__29669\,
            I => \N__29666\
        );

    \I__4859\ : Odrv12
    port map (
            O => \N__29666\,
            I => \sDAC_mem_30Z0Z_3\
        );

    \I__4858\ : InMux
    port map (
            O => \N__29663\,
            I => \N__29660\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__29660\,
            I => \N__29657\
        );

    \I__4856\ : Span4Mux_h
    port map (
            O => \N__29657\,
            I => \N__29654\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__29654\,
            I => \sDAC_mem_31Z0Z_6\
        );

    \I__4854\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29648\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__29648\,
            I => \N__29645\
        );

    \I__4852\ : Span4Mux_h
    port map (
            O => \N__29645\,
            I => \N__29642\
        );

    \I__4851\ : Span4Mux_h
    port map (
            O => \N__29642\,
            I => \N__29639\
        );

    \I__4850\ : Odrv4
    port map (
            O => \N__29639\,
            I => \sDAC_mem_30Z0Z_6\
        );

    \I__4849\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29633\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__29633\,
            I => \N__29630\
        );

    \I__4847\ : Span4Mux_v
    port map (
            O => \N__29630\,
            I => \N__29627\
        );

    \I__4846\ : Odrv4
    port map (
            O => \N__29627\,
            I => \sDAC_data_RNO_24Z0Z_9\
        );

    \I__4845\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29621\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__29621\,
            I => \N__29618\
        );

    \I__4843\ : Span4Mux_h
    port map (
            O => \N__29618\,
            I => \N__29615\
        );

    \I__4842\ : Span4Mux_h
    port map (
            O => \N__29615\,
            I => \N__29612\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__29612\,
            I => \sDAC_mem_16Z0Z_0\
        );

    \I__4840\ : InMux
    port map (
            O => \N__29609\,
            I => \N__29606\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__29606\,
            I => \N__29603\
        );

    \I__4838\ : Span4Mux_h
    port map (
            O => \N__29603\,
            I => \N__29600\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__29600\,
            I => \N__29597\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__29597\,
            I => \sDAC_mem_16Z0Z_1\
        );

    \I__4835\ : InMux
    port map (
            O => \N__29594\,
            I => \N__29591\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__29591\,
            I => \N__29588\
        );

    \I__4833\ : Span4Mux_v
    port map (
            O => \N__29588\,
            I => \N__29585\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__29585\,
            I => \sDAC_data_RNO_28Z0Z_4\
        );

    \I__4831\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29579\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__29579\,
            I => \N__29576\
        );

    \I__4829\ : Span12Mux_h
    port map (
            O => \N__29576\,
            I => \N__29573\
        );

    \I__4828\ : Odrv12
    port map (
            O => \N__29573\,
            I => \sDAC_mem_16Z0Z_2\
        );

    \I__4827\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29567\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__29567\,
            I => \N__29564\
        );

    \I__4825\ : Odrv4
    port map (
            O => \N__29564\,
            I => \sDAC_mem_27Z0Z_1\
        );

    \I__4824\ : InMux
    port map (
            O => \N__29561\,
            I => \N__29558\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__29558\,
            I => \N__29551\
        );

    \I__4822\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29548\
        );

    \I__4821\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29545\
        );

    \I__4820\ : InMux
    port map (
            O => \N__29555\,
            I => \N__29540\
        );

    \I__4819\ : InMux
    port map (
            O => \N__29554\,
            I => \N__29540\
        );

    \I__4818\ : Span12Mux_v
    port map (
            O => \N__29551\,
            I => \N__29535\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__29548\,
            I => \N__29535\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__29545\,
            I => \N_106\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__29540\,
            I => \N_106\
        );

    \I__4814\ : Odrv12
    port map (
            O => \N__29535\,
            I => \N_106\
        );

    \I__4813\ : InMux
    port map (
            O => \N__29528\,
            I => \bfn_14_13_0_\
        );

    \I__4812\ : InMux
    port map (
            O => \N__29525\,
            I => \N__29522\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__29522\,
            I => \N__29519\
        );

    \I__4810\ : Span4Mux_h
    port map (
            O => \N__29519\,
            I => \N__29516\
        );

    \I__4809\ : Odrv4
    port map (
            O => \N__29516\,
            I => \sDAC_mem_24Z0Z_7\
        );

    \I__4808\ : InMux
    port map (
            O => \N__29513\,
            I => \N__29510\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__29510\,
            I => \N__29507\
        );

    \I__4806\ : Span4Mux_h
    port map (
            O => \N__29507\,
            I => \N__29504\
        );

    \I__4805\ : Span4Mux_h
    port map (
            O => \N__29504\,
            I => \N__29501\
        );

    \I__4804\ : Odrv4
    port map (
            O => \N__29501\,
            I => \sDAC_mem_26Z0Z_7\
        );

    \I__4803\ : InMux
    port map (
            O => \N__29498\,
            I => \N__29495\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__29495\,
            I => \N__29492\
        );

    \I__4801\ : Span4Mux_v
    port map (
            O => \N__29492\,
            I => \N__29489\
        );

    \I__4800\ : Span4Mux_h
    port map (
            O => \N__29489\,
            I => \N__29486\
        );

    \I__4799\ : Span4Mux_v
    port map (
            O => \N__29486\,
            I => \N__29483\
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__29483\,
            I => \sDAC_dataZ0Z_10\
        );

    \I__4797\ : InMux
    port map (
            O => \N__29480\,
            I => \N__29477\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__29477\,
            I => \N__29474\
        );

    \I__4795\ : Span4Mux_h
    port map (
            O => \N__29474\,
            I => \N__29471\
        );

    \I__4794\ : Odrv4
    port map (
            O => \N__29471\,
            I => \sDAC_mem_24Z0Z_2\
        );

    \I__4793\ : InMux
    port map (
            O => \N__29468\,
            I => \N__29465\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__29465\,
            I => \sDAC_data_RNO_30Z0Z_5\
        );

    \I__4791\ : InMux
    port map (
            O => \N__29462\,
            I => \N__29459\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__29459\,
            I => \N__29456\
        );

    \I__4789\ : Span4Mux_v
    port map (
            O => \N__29456\,
            I => \N__29453\
        );

    \I__4788\ : Odrv4
    port map (
            O => \N__29453\,
            I => \sDAC_mem_24Z0Z_5\
        );

    \I__4787\ : InMux
    port map (
            O => \N__29450\,
            I => \N__29447\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__29447\,
            I => \N__29444\
        );

    \I__4785\ : Span4Mux_h
    port map (
            O => \N__29444\,
            I => \N__29441\
        );

    \I__4784\ : Odrv4
    port map (
            O => \N__29441\,
            I => \sDAC_data_RNO_30Z0Z_8\
        );

    \I__4783\ : InMux
    port map (
            O => \N__29438\,
            I => \N__29435\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__29435\,
            I => \N__29432\
        );

    \I__4781\ : Span4Mux_h
    port map (
            O => \N__29432\,
            I => \N__29429\
        );

    \I__4780\ : Span4Mux_h
    port map (
            O => \N__29429\,
            I => \N__29426\
        );

    \I__4779\ : Odrv4
    port map (
            O => \N__29426\,
            I => \sDAC_mem_29Z0Z_6\
        );

    \I__4778\ : InMux
    port map (
            O => \N__29423\,
            I => \N__29420\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__29420\,
            I => \N__29417\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__29417\,
            I => \N__29414\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__29414\,
            I => \sDAC_data_RNO_23Z0Z_9\
        );

    \I__4774\ : InMux
    port map (
            O => \N__29411\,
            I => \N__29408\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__29408\,
            I => \N__29404\
        );

    \I__4772\ : CascadeMux
    port map (
            O => \N__29407\,
            I => \N__29401\
        );

    \I__4771\ : Span4Mux_h
    port map (
            O => \N__29404\,
            I => \N__29398\
        );

    \I__4770\ : InMux
    port map (
            O => \N__29401\,
            I => \N__29395\
        );

    \I__4769\ : Odrv4
    port map (
            O => \N__29398\,
            I => \sEEACQZ0Z_15\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__29395\,
            I => \sEEACQZ0Z_15\
        );

    \I__4767\ : CascadeMux
    port map (
            O => \N__29390\,
            I => \N__29387\
        );

    \I__4766\ : InMux
    port map (
            O => \N__29387\,
            I => \N__29384\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__29384\,
            I => \N__29381\
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__29381\,
            I => \sEEACQ_i_15\
        );

    \I__4763\ : InMux
    port map (
            O => \N__29378\,
            I => \N__29374\
        );

    \I__4762\ : CascadeMux
    port map (
            O => \N__29377\,
            I => \N__29371\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__29374\,
            I => \N__29368\
        );

    \I__4760\ : InMux
    port map (
            O => \N__29371\,
            I => \N__29365\
        );

    \I__4759\ : Span4Mux_h
    port map (
            O => \N__29368\,
            I => \N__29362\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__29365\,
            I => \N__29357\
        );

    \I__4757\ : Span4Mux_v
    port map (
            O => \N__29362\,
            I => \N__29357\
        );

    \I__4756\ : Odrv4
    port map (
            O => \N__29357\,
            I => \sEEACQZ0Z_7\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__29354\,
            I => \N__29351\
        );

    \I__4754\ : InMux
    port map (
            O => \N__29351\,
            I => \N__29348\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__29348\,
            I => \sEEACQ_i_7\
        );

    \I__4752\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29342\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__29342\,
            I => \N__29338\
        );

    \I__4750\ : CascadeMux
    port map (
            O => \N__29341\,
            I => \N__29335\
        );

    \I__4749\ : Span12Mux_v
    port map (
            O => \N__29338\,
            I => \N__29332\
        );

    \I__4748\ : InMux
    port map (
            O => \N__29335\,
            I => \N__29329\
        );

    \I__4747\ : Odrv12
    port map (
            O => \N__29332\,
            I => \sEEACQZ0Z_8\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__29329\,
            I => \sEEACQZ0Z_8\
        );

    \I__4745\ : CascadeMux
    port map (
            O => \N__29324\,
            I => \N__29321\
        );

    \I__4744\ : InMux
    port map (
            O => \N__29321\,
            I => \N__29318\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__29318\,
            I => \sEEACQ_i_8\
        );

    \I__4742\ : InMux
    port map (
            O => \N__29315\,
            I => \N__29312\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__29312\,
            I => \N__29309\
        );

    \I__4740\ : Span4Mux_h
    port map (
            O => \N__29309\,
            I => \N__29305\
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__29308\,
            I => \N__29302\
        );

    \I__4738\ : Span4Mux_v
    port map (
            O => \N__29305\,
            I => \N__29299\
        );

    \I__4737\ : InMux
    port map (
            O => \N__29302\,
            I => \N__29296\
        );

    \I__4736\ : Odrv4
    port map (
            O => \N__29299\,
            I => \sEEACQZ0Z_9\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__29296\,
            I => \sEEACQZ0Z_9\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__29291\,
            I => \N__29288\
        );

    \I__4733\ : InMux
    port map (
            O => \N__29288\,
            I => \N__29285\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__29285\,
            I => \sEEACQ_i_9\
        );

    \I__4731\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29279\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29275\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__29278\,
            I => \N__29272\
        );

    \I__4728\ : Span4Mux_h
    port map (
            O => \N__29275\,
            I => \N__29269\
        );

    \I__4727\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29266\
        );

    \I__4726\ : Span4Mux_v
    port map (
            O => \N__29269\,
            I => \N__29261\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__29266\,
            I => \N__29261\
        );

    \I__4724\ : Odrv4
    port map (
            O => \N__29261\,
            I => \sEEACQZ0Z_10\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__29258\,
            I => \N__29255\
        );

    \I__4722\ : InMux
    port map (
            O => \N__29255\,
            I => \N__29252\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__29252\,
            I => \sEEACQ_i_10\
        );

    \I__4720\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29245\
        );

    \I__4719\ : CascadeMux
    port map (
            O => \N__29248\,
            I => \N__29242\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__29245\,
            I => \N__29239\
        );

    \I__4717\ : InMux
    port map (
            O => \N__29242\,
            I => \N__29236\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__29239\,
            I => \N__29233\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__29236\,
            I => \N__29230\
        );

    \I__4714\ : Odrv4
    port map (
            O => \N__29233\,
            I => \sEEACQZ0Z_11\
        );

    \I__4713\ : Odrv4
    port map (
            O => \N__29230\,
            I => \sEEACQZ0Z_11\
        );

    \I__4712\ : CascadeMux
    port map (
            O => \N__29225\,
            I => \N__29222\
        );

    \I__4711\ : InMux
    port map (
            O => \N__29222\,
            I => \N__29219\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__29219\,
            I => \sEEACQ_i_11\
        );

    \I__4709\ : InMux
    port map (
            O => \N__29216\,
            I => \N__29213\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__29213\,
            I => \N__29209\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__29212\,
            I => \N__29206\
        );

    \I__4706\ : Span4Mux_h
    port map (
            O => \N__29209\,
            I => \N__29203\
        );

    \I__4705\ : InMux
    port map (
            O => \N__29206\,
            I => \N__29200\
        );

    \I__4704\ : Odrv4
    port map (
            O => \N__29203\,
            I => \sEEACQZ0Z_12\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__29200\,
            I => \sEEACQZ0Z_12\
        );

    \I__4702\ : CascadeMux
    port map (
            O => \N__29195\,
            I => \N__29192\
        );

    \I__4701\ : InMux
    port map (
            O => \N__29192\,
            I => \N__29189\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__29189\,
            I => \sEEACQ_i_12\
        );

    \I__4699\ : InMux
    port map (
            O => \N__29186\,
            I => \N__29183\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__29183\,
            I => \N__29179\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__29182\,
            I => \N__29176\
        );

    \I__4696\ : Span4Mux_h
    port map (
            O => \N__29179\,
            I => \N__29173\
        );

    \I__4695\ : InMux
    port map (
            O => \N__29176\,
            I => \N__29170\
        );

    \I__4694\ : Odrv4
    port map (
            O => \N__29173\,
            I => \sEEACQZ0Z_13\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__29170\,
            I => \sEEACQZ0Z_13\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__29165\,
            I => \N__29162\
        );

    \I__4691\ : InMux
    port map (
            O => \N__29162\,
            I => \N__29159\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__29159\,
            I => \sEEACQ_i_13\
        );

    \I__4689\ : InMux
    port map (
            O => \N__29156\,
            I => \N__29152\
        );

    \I__4688\ : CascadeMux
    port map (
            O => \N__29155\,
            I => \N__29149\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__29152\,
            I => \N__29146\
        );

    \I__4686\ : InMux
    port map (
            O => \N__29149\,
            I => \N__29143\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__29146\,
            I => \N__29140\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__29143\,
            I => \N__29137\
        );

    \I__4683\ : Odrv4
    port map (
            O => \N__29140\,
            I => \sEEACQZ0Z_14\
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__29137\,
            I => \sEEACQZ0Z_14\
        );

    \I__4681\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29129\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__29129\,
            I => \sEEACQ_i_14\
        );

    \I__4679\ : InMux
    port map (
            O => \N__29126\,
            I => \N__29123\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__29123\,
            I => \sDAC_mem_12Z0Z_3\
        );

    \I__4677\ : InMux
    port map (
            O => \N__29120\,
            I => \N__29116\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__29119\,
            I => \N__29113\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__29116\,
            I => \N__29110\
        );

    \I__4674\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29107\
        );

    \I__4673\ : Span4Mux_h
    port map (
            O => \N__29110\,
            I => \N__29104\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__29107\,
            I => \N__29101\
        );

    \I__4671\ : Odrv4
    port map (
            O => \N__29104\,
            I => \sEEACQZ0Z_0\
        );

    \I__4670\ : Odrv4
    port map (
            O => \N__29101\,
            I => \sEEACQZ0Z_0\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__29096\,
            I => \N__29093\
        );

    \I__4668\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29090\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__29090\,
            I => \sEEACQ_i_0\
        );

    \I__4666\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29083\
        );

    \I__4665\ : CascadeMux
    port map (
            O => \N__29086\,
            I => \N__29080\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__29083\,
            I => \N__29077\
        );

    \I__4663\ : InMux
    port map (
            O => \N__29080\,
            I => \N__29074\
        );

    \I__4662\ : Span4Mux_h
    port map (
            O => \N__29077\,
            I => \N__29071\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__29074\,
            I => \N__29068\
        );

    \I__4660\ : Odrv4
    port map (
            O => \N__29071\,
            I => \sEEACQZ0Z_1\
        );

    \I__4659\ : Odrv4
    port map (
            O => \N__29068\,
            I => \sEEACQZ0Z_1\
        );

    \I__4658\ : CascadeMux
    port map (
            O => \N__29063\,
            I => \N__29060\
        );

    \I__4657\ : InMux
    port map (
            O => \N__29060\,
            I => \N__29057\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__29057\,
            I => \sEEACQ_i_1\
        );

    \I__4655\ : InMux
    port map (
            O => \N__29054\,
            I => \N__29051\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__29051\,
            I => \N__29047\
        );

    \I__4653\ : CascadeMux
    port map (
            O => \N__29050\,
            I => \N__29044\
        );

    \I__4652\ : Span4Mux_h
    port map (
            O => \N__29047\,
            I => \N__29041\
        );

    \I__4651\ : InMux
    port map (
            O => \N__29044\,
            I => \N__29038\
        );

    \I__4650\ : Odrv4
    port map (
            O => \N__29041\,
            I => \sEEACQZ0Z_2\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__29038\,
            I => \sEEACQZ0Z_2\
        );

    \I__4648\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29030\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__29030\,
            I => \sEEACQ_i_2\
        );

    \I__4646\ : InMux
    port map (
            O => \N__29027\,
            I => \N__29024\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__29024\,
            I => \N__29020\
        );

    \I__4644\ : CascadeMux
    port map (
            O => \N__29023\,
            I => \N__29017\
        );

    \I__4643\ : Span4Mux_h
    port map (
            O => \N__29020\,
            I => \N__29014\
        );

    \I__4642\ : InMux
    port map (
            O => \N__29017\,
            I => \N__29011\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__29014\,
            I => \sEEACQZ0Z_3\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__29011\,
            I => \sEEACQZ0Z_3\
        );

    \I__4639\ : CascadeMux
    port map (
            O => \N__29006\,
            I => \N__29003\
        );

    \I__4638\ : InMux
    port map (
            O => \N__29003\,
            I => \N__29000\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__29000\,
            I => \sEEACQ_i_3\
        );

    \I__4636\ : InMux
    port map (
            O => \N__28997\,
            I => \N__28993\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__28996\,
            I => \N__28990\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__28993\,
            I => \N__28987\
        );

    \I__4633\ : InMux
    port map (
            O => \N__28990\,
            I => \N__28984\
        );

    \I__4632\ : Span4Mux_h
    port map (
            O => \N__28987\,
            I => \N__28981\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__28984\,
            I => \N__28978\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__28981\,
            I => \sEEACQZ0Z_4\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__28978\,
            I => \sEEACQZ0Z_4\
        );

    \I__4628\ : CascadeMux
    port map (
            O => \N__28973\,
            I => \N__28970\
        );

    \I__4627\ : InMux
    port map (
            O => \N__28970\,
            I => \N__28967\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__28967\,
            I => \sEEACQ_i_4\
        );

    \I__4625\ : InMux
    port map (
            O => \N__28964\,
            I => \N__28961\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__28961\,
            I => \N__28957\
        );

    \I__4623\ : CascadeMux
    port map (
            O => \N__28960\,
            I => \N__28954\
        );

    \I__4622\ : Span4Mux_h
    port map (
            O => \N__28957\,
            I => \N__28951\
        );

    \I__4621\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28948\
        );

    \I__4620\ : Odrv4
    port map (
            O => \N__28951\,
            I => \sEEACQZ0Z_5\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__28948\,
            I => \sEEACQZ0Z_5\
        );

    \I__4618\ : CascadeMux
    port map (
            O => \N__28943\,
            I => \N__28940\
        );

    \I__4617\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28937\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__28937\,
            I => \sEEACQ_i_5\
        );

    \I__4615\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28931\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__28931\,
            I => \N__28927\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__28930\,
            I => \N__28924\
        );

    \I__4612\ : Span12Mux_v
    port map (
            O => \N__28927\,
            I => \N__28921\
        );

    \I__4611\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28918\
        );

    \I__4610\ : Odrv12
    port map (
            O => \N__28921\,
            I => \sEEACQZ0Z_6\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__28918\,
            I => \sEEACQZ0Z_6\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__28913\,
            I => \N__28910\
        );

    \I__4607\ : InMux
    port map (
            O => \N__28910\,
            I => \N__28907\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__28907\,
            I => \sEEACQ_i_6\
        );

    \I__4605\ : InMux
    port map (
            O => \N__28904\,
            I => \N__28901\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__28901\,
            I => \sDAC_data_2_14_ns_1_4\
        );

    \I__4603\ : InMux
    port map (
            O => \N__28898\,
            I => \N__28895\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__28895\,
            I => \sDAC_data_2_32_ns_1_4\
        );

    \I__4601\ : InMux
    port map (
            O => \N__28892\,
            I => \N__28889\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__28889\,
            I => \N__28886\
        );

    \I__4599\ : Odrv12
    port map (
            O => \N__28886\,
            I => \sDAC_mem_15Z0Z_2\
        );

    \I__4598\ : InMux
    port map (
            O => \N__28883\,
            I => \N__28880\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__28880\,
            I => \N__28877\
        );

    \I__4596\ : Span4Mux_h
    port map (
            O => \N__28877\,
            I => \N__28874\
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__28874\,
            I => \sDAC_mem_14Z0Z_2\
        );

    \I__4594\ : CascadeMux
    port map (
            O => \N__28871\,
            I => \sDAC_data_RNO_18Z0Z_5_cascade_\
        );

    \I__4593\ : InMux
    port map (
            O => \N__28868\,
            I => \N__28865\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__28865\,
            I => \sDAC_data_RNO_19Z0Z_5\
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__28862\,
            I => \sDAC_data_RNO_18Z0Z_6_cascade_\
        );

    \I__4590\ : InMux
    port map (
            O => \N__28859\,
            I => \N__28856\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__28856\,
            I => \N__28853\
        );

    \I__4588\ : Span4Mux_h
    port map (
            O => \N__28853\,
            I => \N__28850\
        );

    \I__4587\ : Odrv4
    port map (
            O => \N__28850\,
            I => \sDAC_data_2_24_ns_1_6\
        );

    \I__4586\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28844\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__28844\,
            I => \N__28841\
        );

    \I__4584\ : Odrv12
    port map (
            O => \N__28841\,
            I => \sDAC_mem_15Z0Z_3\
        );

    \I__4583\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28835\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__28835\,
            I => \N__28832\
        );

    \I__4581\ : Span4Mux_h
    port map (
            O => \N__28832\,
            I => \N__28829\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__28829\,
            I => \sDAC_mem_14Z0Z_3\
        );

    \I__4579\ : InMux
    port map (
            O => \N__28826\,
            I => \N__28823\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__28823\,
            I => \sDAC_data_RNO_19Z0Z_6\
        );

    \I__4577\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28817\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__28817\,
            I => \sDAC_mem_12Z0Z_2\
        );

    \I__4575\ : InMux
    port map (
            O => \N__28814\,
            I => \N__28811\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__28811\,
            I => \sDAC_data_RNO_28Z0Z_8\
        );

    \I__4573\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28805\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__28805\,
            I => \sDAC_mem_16Z0Z_5\
        );

    \I__4571\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28799\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__28799\,
            I => \sDAC_mem_16Z0Z_6\
        );

    \I__4569\ : CascadeMux
    port map (
            O => \N__28796\,
            I => \sDAC_data_RNO_10Z0Z_4_cascade_\
        );

    \I__4568\ : InMux
    port map (
            O => \N__28793\,
            I => \N__28790\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__28790\,
            I => \N__28787\
        );

    \I__4566\ : Span4Mux_h
    port map (
            O => \N__28787\,
            I => \N__28784\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__28784\,
            I => \sDAC_data_RNO_11Z0Z_4\
        );

    \I__4564\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28778\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__28778\,
            I => \N__28775\
        );

    \I__4562\ : Span4Mux_h
    port map (
            O => \N__28775\,
            I => \N__28772\
        );

    \I__4561\ : Odrv4
    port map (
            O => \N__28772\,
            I => \sDAC_data_RNO_5Z0Z_4\
        );

    \I__4560\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28766\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__28766\,
            I => \sDAC_data_RNO_2Z0Z_4\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__28763\,
            I => \sDAC_data_RNO_1Z0Z_4_cascade_\
        );

    \I__4557\ : InMux
    port map (
            O => \N__28760\,
            I => \N__28757\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__28757\,
            I => \sDAC_data_2_41_ns_1_4\
        );

    \I__4555\ : CascadeMux
    port map (
            O => \N__28754\,
            I => \sDAC_data_2_4_cascade_\
        );

    \I__4554\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28748\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__28748\,
            I => \sDAC_data_RNO_15Z0Z_4\
        );

    \I__4552\ : InMux
    port map (
            O => \N__28745\,
            I => \N__28742\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__28742\,
            I => \N__28739\
        );

    \I__4550\ : Span4Mux_h
    port map (
            O => \N__28739\,
            I => \N__28736\
        );

    \I__4549\ : Odrv4
    port map (
            O => \N__28736\,
            I => \sDAC_mem_38Z0Z_3\
        );

    \I__4548\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28730\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__28730\,
            I => \N__28727\
        );

    \I__4546\ : Span4Mux_h
    port map (
            O => \N__28727\,
            I => \N__28724\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__28724\,
            I => \sDAC_mem_39Z0Z_3\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__28721\,
            I => \sDAC_data_2_13_bm_1_6_cascade_\
        );

    \I__4543\ : InMux
    port map (
            O => \N__28718\,
            I => \N__28715\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__28715\,
            I => \sDAC_data_RNO_5Z0Z_6\
        );

    \I__4541\ : InMux
    port map (
            O => \N__28712\,
            I => \N__28709\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__28709\,
            I => \sDAC_mem_6Z0Z_3\
        );

    \I__4539\ : InMux
    port map (
            O => \N__28706\,
            I => \N__28703\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__28703\,
            I => \N__28700\
        );

    \I__4537\ : Odrv12
    port map (
            O => \N__28700\,
            I => \sDAC_mem_38Z0Z_4\
        );

    \I__4536\ : InMux
    port map (
            O => \N__28697\,
            I => \N__28694\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__28694\,
            I => \N__28691\
        );

    \I__4534\ : Span4Mux_v
    port map (
            O => \N__28691\,
            I => \N__28688\
        );

    \I__4533\ : Sp12to4
    port map (
            O => \N__28688\,
            I => \N__28685\
        );

    \I__4532\ : Odrv12
    port map (
            O => \N__28685\,
            I => \sDAC_mem_39Z0Z_4\
        );

    \I__4531\ : CascadeMux
    port map (
            O => \N__28682\,
            I => \sDAC_data_2_13_bm_1_7_cascade_\
        );

    \I__4530\ : InMux
    port map (
            O => \N__28679\,
            I => \N__28676\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__28676\,
            I => \N__28673\
        );

    \I__4528\ : Odrv4
    port map (
            O => \N__28673\,
            I => \sDAC_data_RNO_28Z0Z_6\
        );

    \I__4527\ : InMux
    port map (
            O => \N__28670\,
            I => \N__28667\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__28667\,
            I => \sDAC_mem_16Z0Z_3\
        );

    \I__4525\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28661\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__28661\,
            I => \sDAC_mem_16Z0Z_4\
        );

    \I__4523\ : CascadeMux
    port map (
            O => \N__28658\,
            I => \sDAC_data_RNO_18Z0Z_8_cascade_\
        );

    \I__4522\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28652\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__28652\,
            I => \sDAC_data_2_24_ns_1_8\
        );

    \I__4520\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28646\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__28646\,
            I => \N__28643\
        );

    \I__4518\ : Span4Mux_h
    port map (
            O => \N__28643\,
            I => \N__28640\
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__28640\,
            I => \sDAC_mem_15Z0Z_5\
        );

    \I__4516\ : InMux
    port map (
            O => \N__28637\,
            I => \N__28634\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__28634\,
            I => \N__28631\
        );

    \I__4514\ : Span4Mux_h
    port map (
            O => \N__28631\,
            I => \N__28628\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__28628\,
            I => \sDAC_mem_14Z0Z_5\
        );

    \I__4512\ : InMux
    port map (
            O => \N__28625\,
            I => \N__28622\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__28622\,
            I => \sDAC_data_RNO_19Z0Z_8\
        );

    \I__4510\ : InMux
    port map (
            O => \N__28619\,
            I => \N__28616\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__28616\,
            I => \sDAC_mem_12Z0Z_4\
        );

    \I__4508\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28610\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__28610\,
            I => \sDAC_mem_12Z0Z_5\
        );

    \I__4506\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28604\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__28604\,
            I => \N__28601\
        );

    \I__4504\ : Odrv12
    port map (
            O => \N__28601\,
            I => \sDAC_mem_38Z0Z_2\
        );

    \I__4503\ : InMux
    port map (
            O => \N__28598\,
            I => \N__28595\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__28595\,
            I => \N__28592\
        );

    \I__4501\ : Span4Mux_h
    port map (
            O => \N__28592\,
            I => \N__28589\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__28589\,
            I => \sDAC_mem_39Z0Z_2\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__28586\,
            I => \sDAC_data_2_13_bm_1_5_cascade_\
        );

    \I__4498\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28580\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__28580\,
            I => \sDAC_mem_6Z0Z_2\
        );

    \I__4496\ : InMux
    port map (
            O => \N__28577\,
            I => \N__28574\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__28574\,
            I => \sDAC_mem_18Z0Z_3\
        );

    \I__4494\ : InMux
    port map (
            O => \N__28571\,
            I => \N__28568\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__28568\,
            I => \sDAC_mem_18Z0Z_4\
        );

    \I__4492\ : InMux
    port map (
            O => \N__28565\,
            I => \N__28562\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__28562\,
            I => \N__28559\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__28559\,
            I => \sDAC_data_RNO_29Z0Z_8\
        );

    \I__4489\ : InMux
    port map (
            O => \N__28556\,
            I => \N__28553\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__28553\,
            I => \sDAC_mem_18Z0Z_5\
        );

    \I__4487\ : InMux
    port map (
            O => \N__28550\,
            I => \N__28547\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__28547\,
            I => \sDAC_mem_18Z0Z_6\
        );

    \I__4485\ : CEMux
    port map (
            O => \N__28544\,
            I => \N__28541\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__28541\,
            I => \N__28537\
        );

    \I__4483\ : CEMux
    port map (
            O => \N__28540\,
            I => \N__28534\
        );

    \I__4482\ : Span4Mux_h
    port map (
            O => \N__28537\,
            I => \N__28531\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__28534\,
            I => \N__28528\
        );

    \I__4480\ : Span4Mux_v
    port map (
            O => \N__28531\,
            I => \N__28523\
        );

    \I__4479\ : Span4Mux_v
    port map (
            O => \N__28528\,
            I => \N__28523\
        );

    \I__4478\ : Span4Mux_h
    port map (
            O => \N__28523\,
            I => \N__28520\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__28520\,
            I => \sDAC_mem_18_1_sqmuxa\
        );

    \I__4476\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28514\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__28514\,
            I => \N__28511\
        );

    \I__4474\ : Span12Mux_v
    port map (
            O => \N__28511\,
            I => \N__28508\
        );

    \I__4473\ : Odrv12
    port map (
            O => \N__28508\,
            I => \sDAC_mem_15Z0Z_4\
        );

    \I__4472\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28502\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__28502\,
            I => \N__28499\
        );

    \I__4470\ : Span4Mux_h
    port map (
            O => \N__28499\,
            I => \N__28496\
        );

    \I__4469\ : Odrv4
    port map (
            O => \N__28496\,
            I => \sDAC_mem_14Z0Z_4\
        );

    \I__4468\ : CascadeMux
    port map (
            O => \N__28493\,
            I => \sDAC_data_RNO_18Z0Z_7_cascade_\
        );

    \I__4467\ : InMux
    port map (
            O => \N__28490\,
            I => \N__28487\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__28487\,
            I => \sDAC_data_RNO_19Z0Z_7\
        );

    \I__4465\ : CEMux
    port map (
            O => \N__28484\,
            I => \N__28481\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__28481\,
            I => \sDAC_mem_36_1_sqmuxa\
        );

    \I__4463\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28475\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__28475\,
            I => \sDAC_data_RNO_29Z0Z_6\
        );

    \I__4461\ : InMux
    port map (
            O => \N__28472\,
            I => \sRAM_pointer_read_cry_9\
        );

    \I__4460\ : InMux
    port map (
            O => \N__28469\,
            I => \sRAM_pointer_read_cry_10\
        );

    \I__4459\ : InMux
    port map (
            O => \N__28466\,
            I => \sRAM_pointer_read_cry_11\
        );

    \I__4458\ : InMux
    port map (
            O => \N__28463\,
            I => \sRAM_pointer_read_cry_12\
        );

    \I__4457\ : InMux
    port map (
            O => \N__28460\,
            I => \sRAM_pointer_read_cry_13\
        );

    \I__4456\ : InMux
    port map (
            O => \N__28457\,
            I => \sRAM_pointer_read_cry_14\
        );

    \I__4455\ : InMux
    port map (
            O => \N__28454\,
            I => \bfn_13_20_0_\
        );

    \I__4454\ : InMux
    port map (
            O => \N__28451\,
            I => \sRAM_pointer_read_cry_16\
        );

    \I__4453\ : InMux
    port map (
            O => \N__28448\,
            I => \sRAM_pointer_read_cry_17\
        );

    \I__4452\ : CEMux
    port map (
            O => \N__28445\,
            I => \N__28436\
        );

    \I__4451\ : CEMux
    port map (
            O => \N__28444\,
            I => \N__28436\
        );

    \I__4450\ : CEMux
    port map (
            O => \N__28443\,
            I => \N__28436\
        );

    \I__4449\ : GlobalMux
    port map (
            O => \N__28436\,
            I => \N__28433\
        );

    \I__4448\ : gio2CtrlBuf
    port map (
            O => \N__28433\,
            I => \N_28_g\
        );

    \I__4447\ : InMux
    port map (
            O => \N__28430\,
            I => \sRAM_pointer_read_cry_0\
        );

    \I__4446\ : InMux
    port map (
            O => \N__28427\,
            I => \sRAM_pointer_read_cry_1\
        );

    \I__4445\ : InMux
    port map (
            O => \N__28424\,
            I => \sRAM_pointer_read_cry_2\
        );

    \I__4444\ : InMux
    port map (
            O => \N__28421\,
            I => \sRAM_pointer_read_cry_3\
        );

    \I__4443\ : InMux
    port map (
            O => \N__28418\,
            I => \sRAM_pointer_read_cry_4\
        );

    \I__4442\ : InMux
    port map (
            O => \N__28415\,
            I => \sRAM_pointer_read_cry_5\
        );

    \I__4441\ : InMux
    port map (
            O => \N__28412\,
            I => \sRAM_pointer_read_cry_6\
        );

    \I__4440\ : InMux
    port map (
            O => \N__28409\,
            I => \bfn_13_19_0_\
        );

    \I__4439\ : InMux
    port map (
            O => \N__28406\,
            I => \sRAM_pointer_read_cry_8\
        );

    \I__4438\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28400\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__28400\,
            I => un1_sacqtime_cry_20_sf
        );

    \I__4436\ : InMux
    port map (
            O => \N__28397\,
            I => \N__28394\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__28394\,
            I => un1_sacqtime_cry_21_sf
        );

    \I__4434\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28388\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__28388\,
            I => un1_sacqtime_cry_22_sf
        );

    \I__4432\ : InMux
    port map (
            O => \N__28385\,
            I => \N__28382\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__28382\,
            I => un1_sacqtime_cry_23_sf
        );

    \I__4430\ : InMux
    port map (
            O => \N__28379\,
            I => \bfn_13_17_0_\
        );

    \I__4429\ : CascadeMux
    port map (
            O => \N__28376\,
            I => \N__28373\
        );

    \I__4428\ : InMux
    port map (
            O => \N__28373\,
            I => \N__28367\
        );

    \I__4427\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28367\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__28367\,
            I => \sADC_clk_prevZ0\
        );

    \I__4425\ : CascadeMux
    port map (
            O => \N__28364\,
            I => \N_71_cascade_\
        );

    \I__4424\ : InMux
    port map (
            O => \N__28361\,
            I => \bfn_13_18_0_\
        );

    \I__4423\ : InMux
    port map (
            O => \N__28358\,
            I => \N__28354\
        );

    \I__4422\ : CascadeMux
    port map (
            O => \N__28357\,
            I => \N__28351\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__28354\,
            I => \N__28348\
        );

    \I__4420\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28345\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__28348\,
            I => \N__28342\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__28345\,
            I => \sCounter_i_11\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__28342\,
            I => \sCounter_i_11\
        );

    \I__4416\ : InMux
    port map (
            O => \N__28337\,
            I => \N__28333\
        );

    \I__4415\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28330\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__28333\,
            I => \N__28327\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__28330\,
            I => \N__28322\
        );

    \I__4412\ : Span4Mux_v
    port map (
            O => \N__28327\,
            I => \N__28322\
        );

    \I__4411\ : Odrv4
    port map (
            O => \N__28322\,
            I => \sCounter_i_12\
        );

    \I__4410\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28315\
        );

    \I__4409\ : CascadeMux
    port map (
            O => \N__28318\,
            I => \N__28312\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__28315\,
            I => \N__28309\
        );

    \I__4407\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28306\
        );

    \I__4406\ : Span4Mux_v
    port map (
            O => \N__28309\,
            I => \N__28303\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__28306\,
            I => \sCounter_i_13\
        );

    \I__4404\ : Odrv4
    port map (
            O => \N__28303\,
            I => \sCounter_i_13\
        );

    \I__4403\ : InMux
    port map (
            O => \N__28298\,
            I => \N__28294\
        );

    \I__4402\ : CascadeMux
    port map (
            O => \N__28297\,
            I => \N__28291\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__28294\,
            I => \N__28288\
        );

    \I__4400\ : InMux
    port map (
            O => \N__28291\,
            I => \N__28285\
        );

    \I__4399\ : Span4Mux_v
    port map (
            O => \N__28288\,
            I => \N__28282\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__28285\,
            I => \sCounter_i_14\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__28282\,
            I => \sCounter_i_14\
        );

    \I__4396\ : InMux
    port map (
            O => \N__28277\,
            I => \N__28274\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__28274\,
            I => \N__28270\
        );

    \I__4394\ : InMux
    port map (
            O => \N__28273\,
            I => \N__28267\
        );

    \I__4393\ : Span4Mux_v
    port map (
            O => \N__28270\,
            I => \N__28264\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__28267\,
            I => \sCounter_i_15\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__28264\,
            I => \sCounter_i_15\
        );

    \I__4390\ : InMux
    port map (
            O => \N__28259\,
            I => \N__28256\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__28256\,
            I => un1_sacqtime_cry_16_sf
        );

    \I__4388\ : InMux
    port map (
            O => \N__28253\,
            I => \N__28250\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__28250\,
            I => un1_sacqtime_cry_17_sf
        );

    \I__4386\ : InMux
    port map (
            O => \N__28247\,
            I => \N__28244\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__28244\,
            I => un1_sacqtime_cry_18_sf
        );

    \I__4384\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28238\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__28238\,
            I => un1_sacqtime_cry_19_sf
        );

    \I__4382\ : InMux
    port map (
            O => \N__28235\,
            I => \N__28231\
        );

    \I__4381\ : CascadeMux
    port map (
            O => \N__28234\,
            I => \N__28228\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__28231\,
            I => \N__28225\
        );

    \I__4379\ : InMux
    port map (
            O => \N__28228\,
            I => \N__28222\
        );

    \I__4378\ : Span4Mux_v
    port map (
            O => \N__28225\,
            I => \N__28219\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__28222\,
            I => \sCounter_i_3\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__28219\,
            I => \sCounter_i_3\
        );

    \I__4375\ : InMux
    port map (
            O => \N__28214\,
            I => \N__28210\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__28213\,
            I => \N__28207\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__28210\,
            I => \N__28204\
        );

    \I__4372\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28201\
        );

    \I__4371\ : Span4Mux_v
    port map (
            O => \N__28204\,
            I => \N__28198\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__28201\,
            I => \sCounter_i_4\
        );

    \I__4369\ : Odrv4
    port map (
            O => \N__28198\,
            I => \sCounter_i_4\
        );

    \I__4368\ : InMux
    port map (
            O => \N__28193\,
            I => \N__28190\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__28190\,
            I => \N__28186\
        );

    \I__4366\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28183\
        );

    \I__4365\ : Span4Mux_v
    port map (
            O => \N__28186\,
            I => \N__28180\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__28183\,
            I => \sCounter_i_5\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__28180\,
            I => \sCounter_i_5\
        );

    \I__4362\ : InMux
    port map (
            O => \N__28175\,
            I => \N__28171\
        );

    \I__4361\ : CascadeMux
    port map (
            O => \N__28174\,
            I => \N__28168\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__28171\,
            I => \N__28165\
        );

    \I__4359\ : InMux
    port map (
            O => \N__28168\,
            I => \N__28162\
        );

    \I__4358\ : Span4Mux_v
    port map (
            O => \N__28165\,
            I => \N__28159\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__28162\,
            I => \sCounter_i_6\
        );

    \I__4356\ : Odrv4
    port map (
            O => \N__28159\,
            I => \sCounter_i_6\
        );

    \I__4355\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28151\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__28151\,
            I => \N__28147\
        );

    \I__4353\ : InMux
    port map (
            O => \N__28150\,
            I => \N__28144\
        );

    \I__4352\ : Span4Mux_v
    port map (
            O => \N__28147\,
            I => \N__28141\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__28144\,
            I => \sCounter_i_7\
        );

    \I__4350\ : Odrv4
    port map (
            O => \N__28141\,
            I => \sCounter_i_7\
        );

    \I__4349\ : InMux
    port map (
            O => \N__28136\,
            I => \N__28132\
        );

    \I__4348\ : CascadeMux
    port map (
            O => \N__28135\,
            I => \N__28129\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__28132\,
            I => \N__28126\
        );

    \I__4346\ : InMux
    port map (
            O => \N__28129\,
            I => \N__28123\
        );

    \I__4345\ : Span4Mux_v
    port map (
            O => \N__28126\,
            I => \N__28120\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__28123\,
            I => \sCounter_i_8\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__28120\,
            I => \sCounter_i_8\
        );

    \I__4342\ : InMux
    port map (
            O => \N__28115\,
            I => \N__28112\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__28112\,
            I => \N__28108\
        );

    \I__4340\ : InMux
    port map (
            O => \N__28111\,
            I => \N__28105\
        );

    \I__4339\ : Span4Mux_v
    port map (
            O => \N__28108\,
            I => \N__28102\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__28105\,
            I => \sCounter_i_9\
        );

    \I__4337\ : Odrv4
    port map (
            O => \N__28102\,
            I => \sCounter_i_9\
        );

    \I__4336\ : InMux
    port map (
            O => \N__28097\,
            I => \N__28093\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__28096\,
            I => \N__28090\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__28093\,
            I => \N__28087\
        );

    \I__4333\ : InMux
    port map (
            O => \N__28090\,
            I => \N__28084\
        );

    \I__4332\ : Span4Mux_v
    port map (
            O => \N__28087\,
            I => \N__28081\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__28084\,
            I => \sCounter_i_10\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__28081\,
            I => \sCounter_i_10\
        );

    \I__4329\ : InMux
    port map (
            O => \N__28076\,
            I => \N__28073\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__28073\,
            I => \sDAC_data_RNO_31Z0Z_5\
        );

    \I__4327\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28067\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__28067\,
            I => \sDAC_mem_26Z0Z_2\
        );

    \I__4325\ : InMux
    port map (
            O => \N__28064\,
            I => \N__28061\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__28061\,
            I => \N__28058\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__28058\,
            I => \sDAC_data_RNO_31Z0Z_8\
        );

    \I__4322\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28052\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__28052\,
            I => \sDAC_mem_26Z0Z_5\
        );

    \I__4320\ : CEMux
    port map (
            O => \N__28049\,
            I => \N__28046\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__28046\,
            I => \N__28042\
        );

    \I__4318\ : CEMux
    port map (
            O => \N__28045\,
            I => \N__28039\
        );

    \I__4317\ : Span4Mux_h
    port map (
            O => \N__28042\,
            I => \N__28034\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__28039\,
            I => \N__28034\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__28034\,
            I => \N__28031\
        );

    \I__4314\ : Span4Mux_h
    port map (
            O => \N__28031\,
            I => \N__28028\
        );

    \I__4313\ : Odrv4
    port map (
            O => \N__28028\,
            I => \sDAC_mem_26_1_sqmuxa\
        );

    \I__4312\ : InMux
    port map (
            O => \N__28025\,
            I => \N__28022\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__28022\,
            I => \N__28019\
        );

    \I__4310\ : Span4Mux_h
    port map (
            O => \N__28019\,
            I => \N__28016\
        );

    \I__4309\ : Span4Mux_v
    port map (
            O => \N__28016\,
            I => \N__28013\
        );

    \I__4308\ : Span4Mux_v
    port map (
            O => \N__28013\,
            I => \N__28010\
        );

    \I__4307\ : Odrv4
    port map (
            O => \N__28010\,
            I => \spi_master_inst.sclk_gen_u0.delay_clk_iZ0\
        );

    \I__4306\ : InMux
    port map (
            O => \N__28007\,
            I => \N__28004\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__28004\,
            I => \N__28001\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__28001\,
            I => \N__27997\
        );

    \I__4303\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27994\
        );

    \I__4302\ : Span4Mux_h
    port map (
            O => \N__27997\,
            I => \N__27990\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__27994\,
            I => \N__27986\
        );

    \I__4300\ : InMux
    port map (
            O => \N__27993\,
            I => \N__27983\
        );

    \I__4299\ : Span4Mux_v
    port map (
            O => \N__27990\,
            I => \N__27980\
        );

    \I__4298\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27977\
        );

    \I__4297\ : Odrv4
    port map (
            O => \N__27986\,
            I => \spi_master_inst.sclk_gen_u0.div_clk_iZ0\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__27983\,
            I => \spi_master_inst.sclk_gen_u0.div_clk_iZ0\
        );

    \I__4295\ : Odrv4
    port map (
            O => \N__27980\,
            I => \spi_master_inst.sclk_gen_u0.div_clk_iZ0\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__27977\,
            I => \spi_master_inst.sclk_gen_u0.div_clk_iZ0\
        );

    \I__4293\ : CEMux
    port map (
            O => \N__27968\,
            I => \N__27965\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__27965\,
            I => \N__27962\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__27962\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i\
        );

    \I__4290\ : InMux
    port map (
            O => \N__27959\,
            I => \N__27953\
        );

    \I__4289\ : InMux
    port map (
            O => \N__27958\,
            I => \N__27953\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__27953\,
            I => \N__27950\
        );

    \I__4287\ : Span4Mux_h
    port map (
            O => \N__27950\,
            I => \N__27947\
        );

    \I__4286\ : Span4Mux_h
    port map (
            O => \N__27947\,
            I => \N__27944\
        );

    \I__4285\ : Span4Mux_h
    port map (
            O => \N__27944\,
            I => \N__27940\
        );

    \I__4284\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27937\
        );

    \I__4283\ : Span4Mux_v
    port map (
            O => \N__27940\,
            I => \N__27934\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__27937\,
            I => \spi_master_inst.sclk_gen_u0.falling_count_start_iZ0\
        );

    \I__4281\ : Odrv4
    port map (
            O => \N__27934\,
            I => \spi_master_inst.sclk_gen_u0.falling_count_start_iZ0\
        );

    \I__4280\ : InMux
    port map (
            O => \N__27929\,
            I => \N__27911\
        );

    \I__4279\ : InMux
    port map (
            O => \N__27928\,
            I => \N__27911\
        );

    \I__4278\ : InMux
    port map (
            O => \N__27927\,
            I => \N__27911\
        );

    \I__4277\ : InMux
    port map (
            O => \N__27926\,
            I => \N__27911\
        );

    \I__4276\ : InMux
    port map (
            O => \N__27925\,
            I => \N__27911\
        );

    \I__4275\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27904\
        );

    \I__4274\ : InMux
    port map (
            O => \N__27923\,
            I => \N__27904\
        );

    \I__4273\ : InMux
    port map (
            O => \N__27922\,
            I => \N__27904\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__27911\,
            I => \N__27899\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__27904\,
            I => \N__27899\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__27899\,
            I => \spi_master_inst.sclk_gen_u0.falling_count_start_i_i\
        );

    \I__4269\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27893\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__27893\,
            I => \N__27889\
        );

    \I__4267\ : InMux
    port map (
            O => \N__27892\,
            I => \N__27886\
        );

    \I__4266\ : Span4Mux_v
    port map (
            O => \N__27889\,
            I => \N__27883\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__27886\,
            I => \sCounter_i_0\
        );

    \I__4264\ : Odrv4
    port map (
            O => \N__27883\,
            I => \sCounter_i_0\
        );

    \I__4263\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27874\
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__27877\,
            I => \N__27871\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__27874\,
            I => \N__27868\
        );

    \I__4260\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27865\
        );

    \I__4259\ : Span4Mux_v
    port map (
            O => \N__27868\,
            I => \N__27862\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__27865\,
            I => \sCounter_i_1\
        );

    \I__4257\ : Odrv4
    port map (
            O => \N__27862\,
            I => \sCounter_i_1\
        );

    \I__4256\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27853\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__27856\,
            I => \N__27850\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__27853\,
            I => \N__27847\
        );

    \I__4253\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27844\
        );

    \I__4252\ : Span4Mux_v
    port map (
            O => \N__27847\,
            I => \N__27841\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__27844\,
            I => \sCounter_i_2\
        );

    \I__4250\ : Odrv4
    port map (
            O => \N__27841\,
            I => \sCounter_i_2\
        );

    \I__4249\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27833\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__27833\,
            I => \N__27830\
        );

    \I__4247\ : Span4Mux_h
    port map (
            O => \N__27830\,
            I => \N__27827\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__27827\,
            I => \sDAC_mem_26Z0Z_1\
        );

    \I__4245\ : CascadeMux
    port map (
            O => \N__27824\,
            I => \sDAC_data_RNO_30Z0Z_4_cascade_\
        );

    \I__4244\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27818\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__27818\,
            I => \sDAC_data_RNO_31Z0Z_4\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__27815\,
            I => \sDAC_data_2_39_ns_1_4_cascade_\
        );

    \I__4241\ : InMux
    port map (
            O => \N__27812\,
            I => \N__27809\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__27809\,
            I => \N__27806\
        );

    \I__4239\ : Span4Mux_h
    port map (
            O => \N__27806\,
            I => \N__27803\
        );

    \I__4238\ : Odrv4
    port map (
            O => \N__27803\,
            I => \sDAC_mem_28Z0Z_1\
        );

    \I__4237\ : InMux
    port map (
            O => \N__27800\,
            I => \N__27797\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__27797\,
            I => \N__27794\
        );

    \I__4235\ : Span12Mux_h
    port map (
            O => \N__27794\,
            I => \N__27791\
        );

    \I__4234\ : Odrv12
    port map (
            O => \N__27791\,
            I => \sDAC_mem_29Z0Z_1\
        );

    \I__4233\ : InMux
    port map (
            O => \N__27788\,
            I => \N__27785\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__27785\,
            I => \sDAC_data_RNO_23Z0Z_4\
        );

    \I__4231\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27779\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__27779\,
            I => \N__27776\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__27776\,
            I => \N__27773\
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__27773\,
            I => \sDAC_mem_31Z0Z_1\
        );

    \I__4227\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27767\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__27767\,
            I => \N__27764\
        );

    \I__4225\ : Span12Mux_h
    port map (
            O => \N__27764\,
            I => \N__27761\
        );

    \I__4224\ : Odrv12
    port map (
            O => \N__27761\,
            I => \sDAC_mem_30Z0Z_1\
        );

    \I__4223\ : InMux
    port map (
            O => \N__27758\,
            I => \N__27755\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__27755\,
            I => \sDAC_data_RNO_24Z0Z_4\
        );

    \I__4221\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27749\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__27749\,
            I => \sDAC_mem_24Z0Z_1\
        );

    \I__4219\ : CEMux
    port map (
            O => \N__27746\,
            I => \N__27742\
        );

    \I__4218\ : CEMux
    port map (
            O => \N__27745\,
            I => \N__27738\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__27742\,
            I => \N__27735\
        );

    \I__4216\ : CEMux
    port map (
            O => \N__27741\,
            I => \N__27732\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__27738\,
            I => \N__27729\
        );

    \I__4214\ : Span4Mux_v
    port map (
            O => \N__27735\,
            I => \N__27726\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__27732\,
            I => \N__27723\
        );

    \I__4212\ : Span4Mux_v
    port map (
            O => \N__27729\,
            I => \N__27720\
        );

    \I__4211\ : Span4Mux_h
    port map (
            O => \N__27726\,
            I => \N__27715\
        );

    \I__4210\ : Span4Mux_v
    port map (
            O => \N__27723\,
            I => \N__27715\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__27720\,
            I => \sDAC_mem_24_1_sqmuxa\
        );

    \I__4208\ : Odrv4
    port map (
            O => \N__27715\,
            I => \sDAC_mem_24_1_sqmuxa\
        );

    \I__4207\ : InMux
    port map (
            O => \N__27710\,
            I => \N__27707\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__27707\,
            I => \N__27704\
        );

    \I__4205\ : Span4Mux_h
    port map (
            O => \N__27704\,
            I => \N__27701\
        );

    \I__4204\ : Span4Mux_h
    port map (
            O => \N__27701\,
            I => \N__27698\
        );

    \I__4203\ : Odrv4
    port map (
            O => \N__27698\,
            I => \sDAC_mem_26Z0Z_6\
        );

    \I__4202\ : InMux
    port map (
            O => \N__27695\,
            I => \N__27692\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__27692\,
            I => \sDAC_data_RNO_31Z0Z_9\
        );

    \I__4200\ : CascadeMux
    port map (
            O => \N__27689\,
            I => \sDAC_data_RNO_30Z0Z_7_cascade_\
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__27686\,
            I => \sDAC_data_2_39_ns_1_7_cascade_\
        );

    \I__4198\ : InMux
    port map (
            O => \N__27683\,
            I => \N__27680\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__27680\,
            I => \N__27677\
        );

    \I__4196\ : Span4Mux_h
    port map (
            O => \N__27677\,
            I => \N__27674\
        );

    \I__4195\ : Odrv4
    port map (
            O => \N__27674\,
            I => \sDAC_mem_26Z0Z_4\
        );

    \I__4194\ : InMux
    port map (
            O => \N__27671\,
            I => \N__27668\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__27668\,
            I => \sDAC_data_RNO_31Z0Z_7\
        );

    \I__4192\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27662\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__27662\,
            I => \N__27659\
        );

    \I__4190\ : Span4Mux_v
    port map (
            O => \N__27659\,
            I => \N__27656\
        );

    \I__4189\ : Span4Mux_h
    port map (
            O => \N__27656\,
            I => \N__27653\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__27653\,
            I => \sDAC_mem_29Z0Z_4\
        );

    \I__4187\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27647\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__27647\,
            I => \N__27644\
        );

    \I__4185\ : Span4Mux_h
    port map (
            O => \N__27644\,
            I => \N__27641\
        );

    \I__4184\ : Span4Mux_v
    port map (
            O => \N__27641\,
            I => \N__27638\
        );

    \I__4183\ : Odrv4
    port map (
            O => \N__27638\,
            I => \sDAC_mem_28Z0Z_4\
        );

    \I__4182\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27632\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__27632\,
            I => \sDAC_data_RNO_23Z0Z_7\
        );

    \I__4180\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27626\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__27626\,
            I => \N__27623\
        );

    \I__4178\ : Span4Mux_h
    port map (
            O => \N__27623\,
            I => \N__27620\
        );

    \I__4177\ : Odrv4
    port map (
            O => \N__27620\,
            I => \sDAC_mem_30Z0Z_4\
        );

    \I__4176\ : InMux
    port map (
            O => \N__27617\,
            I => \N__27614\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__27614\,
            I => \N__27611\
        );

    \I__4174\ : Span4Mux_v
    port map (
            O => \N__27611\,
            I => \N__27608\
        );

    \I__4173\ : Span4Mux_h
    port map (
            O => \N__27608\,
            I => \N__27605\
        );

    \I__4172\ : Odrv4
    port map (
            O => \N__27605\,
            I => \sDAC_mem_31Z0Z_4\
        );

    \I__4171\ : InMux
    port map (
            O => \N__27602\,
            I => \N__27599\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__27599\,
            I => \sDAC_data_RNO_24Z0Z_7\
        );

    \I__4169\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27593\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__27593\,
            I => \sDAC_mem_24Z0Z_4\
        );

    \I__4167\ : InMux
    port map (
            O => \N__27590\,
            I => \N__27587\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__27587\,
            I => \sDAC_data_2_39_ns_1_8\
        );

    \I__4165\ : InMux
    port map (
            O => \N__27584\,
            I => \N__27581\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__27581\,
            I => \sDAC_mem_12Z0Z_0\
        );

    \I__4163\ : InMux
    port map (
            O => \N__27578\,
            I => \N__27575\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__27575\,
            I => \sDAC_mem_12Z0Z_1\
        );

    \I__4161\ : InMux
    port map (
            O => \N__27572\,
            I => \N__27569\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__27569\,
            I => \N__27566\
        );

    \I__4159\ : Span4Mux_h
    port map (
            O => \N__27566\,
            I => \N__27563\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__27563\,
            I => \sDAC_mem_31Z0Z_5\
        );

    \I__4157\ : InMux
    port map (
            O => \N__27560\,
            I => \N__27557\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__27557\,
            I => \N__27554\
        );

    \I__4155\ : Span4Mux_h
    port map (
            O => \N__27554\,
            I => \N__27551\
        );

    \I__4154\ : Span4Mux_v
    port map (
            O => \N__27551\,
            I => \N__27548\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__27548\,
            I => \sDAC_mem_30Z0Z_5\
        );

    \I__4152\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27542\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__27542\,
            I => \N__27539\
        );

    \I__4150\ : Span4Mux_v
    port map (
            O => \N__27539\,
            I => \N__27536\
        );

    \I__4149\ : Span4Mux_h
    port map (
            O => \N__27536\,
            I => \N__27533\
        );

    \I__4148\ : Odrv4
    port map (
            O => \N__27533\,
            I => \sDAC_mem_29Z0Z_5\
        );

    \I__4147\ : InMux
    port map (
            O => \N__27530\,
            I => \N__27527\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__27527\,
            I => \sDAC_data_RNO_24Z0Z_8\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__27524\,
            I => \sDAC_data_RNO_23Z0Z_8_cascade_\
        );

    \I__4144\ : InMux
    port map (
            O => \N__27521\,
            I => \N__27518\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__27518\,
            I => \N__27515\
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__27515\,
            I => \sDAC_data_RNO_11Z0Z_8\
        );

    \I__4141\ : InMux
    port map (
            O => \N__27512\,
            I => \N__27509\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__27509\,
            I => \sDAC_mem_28Z0Z_5\
        );

    \I__4139\ : InMux
    port map (
            O => \N__27506\,
            I => \N__27503\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__27503\,
            I => \N__27500\
        );

    \I__4137\ : Span4Mux_v
    port map (
            O => \N__27500\,
            I => \N__27497\
        );

    \I__4136\ : Span4Mux_h
    port map (
            O => \N__27497\,
            I => \N__27494\
        );

    \I__4135\ : Odrv4
    port map (
            O => \N__27494\,
            I => \sDAC_mem_24Z0Z_6\
        );

    \I__4134\ : CascadeMux
    port map (
            O => \N__27491\,
            I => \sDAC_data_RNO_30Z0Z_9_cascade_\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__27488\,
            I => \sDAC_data_2_39_ns_1_9_cascade_\
        );

    \I__4132\ : InMux
    port map (
            O => \N__27485\,
            I => \N__27482\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__27482\,
            I => \N__27479\
        );

    \I__4130\ : Odrv12
    port map (
            O => \N__27479\,
            I => \sDAC_mem_40Z0Z_1\
        );

    \I__4129\ : InMux
    port map (
            O => \N__27476\,
            I => \N__27473\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__27473\,
            I => \N__27470\
        );

    \I__4127\ : Span4Mux_v
    port map (
            O => \N__27470\,
            I => \N__27467\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__27467\,
            I => \sDAC_mem_8Z0Z_1\
        );

    \I__4125\ : CascadeMux
    port map (
            O => \N__27464\,
            I => \sDAC_data_2_20_am_1_4_cascade_\
        );

    \I__4124\ : CascadeMux
    port map (
            O => \N__27461\,
            I => \sDAC_data_RNO_7Z0Z_4_cascade_\
        );

    \I__4123\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27455\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__27455\,
            I => \sDAC_data_RNO_8Z0Z_4\
        );

    \I__4121\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27449\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__27449\,
            I => \N__27446\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__27446\,
            I => \sDAC_mem_15Z0Z_0\
        );

    \I__4118\ : InMux
    port map (
            O => \N__27443\,
            I => \N__27440\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__27440\,
            I => \N__27437\
        );

    \I__4116\ : Span4Mux_v
    port map (
            O => \N__27437\,
            I => \N__27434\
        );

    \I__4115\ : Odrv4
    port map (
            O => \N__27434\,
            I => \sDAC_mem_14Z0Z_0\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__27431\,
            I => \sDAC_data_RNO_18Z0Z_3_cascade_\
        );

    \I__4113\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27425\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__27425\,
            I => \sDAC_data_RNO_19Z0Z_3\
        );

    \I__4111\ : CascadeMux
    port map (
            O => \N__27422\,
            I => \sDAC_data_RNO_18Z0Z_4_cascade_\
        );

    \I__4110\ : InMux
    port map (
            O => \N__27419\,
            I => \N__27416\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__27416\,
            I => \sDAC_data_2_24_ns_1_4\
        );

    \I__4108\ : InMux
    port map (
            O => \N__27413\,
            I => \N__27410\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__27410\,
            I => \N__27407\
        );

    \I__4106\ : Odrv4
    port map (
            O => \N__27407\,
            I => \sDAC_mem_15Z0Z_1\
        );

    \I__4105\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27401\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__27401\,
            I => \N__27398\
        );

    \I__4103\ : Span4Mux_v
    port map (
            O => \N__27398\,
            I => \N__27395\
        );

    \I__4102\ : Odrv4
    port map (
            O => \N__27395\,
            I => \sDAC_mem_14Z0Z_1\
        );

    \I__4101\ : InMux
    port map (
            O => \N__27392\,
            I => \N__27389\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__27389\,
            I => \sDAC_data_RNO_19Z0Z_4\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__27386\,
            I => \sDAC_data_2_8_cascade_\
        );

    \I__4098\ : CascadeMux
    port map (
            O => \N__27383\,
            I => \sDAC_data_2_32_ns_1_8_cascade_\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__27380\,
            I => \sDAC_data_RNO_10Z0Z_8_cascade_\
        );

    \I__4096\ : InMux
    port map (
            O => \N__27377\,
            I => \N__27374\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__27374\,
            I => \sDAC_data_2_41_ns_1_8\
        );

    \I__4094\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27368\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__27368\,
            I => \sDAC_mem_34Z0Z_1\
        );

    \I__4092\ : InMux
    port map (
            O => \N__27365\,
            I => \N__27362\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__27362\,
            I => \N__27359\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__27359\,
            I => \sDAC_mem_2Z0Z_1\
        );

    \I__4089\ : InMux
    port map (
            O => \N__27356\,
            I => \N__27353\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__27353\,
            I => \sDAC_mem_3Z0Z_1\
        );

    \I__4087\ : InMux
    port map (
            O => \N__27350\,
            I => \N__27347\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__27347\,
            I => \N__27344\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__27344\,
            I => \N__27341\
        );

    \I__4084\ : Span4Mux_h
    port map (
            O => \N__27341\,
            I => \N__27338\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__27338\,
            I => \sDAC_mem_35Z0Z_1\
        );

    \I__4082\ : CascadeMux
    port map (
            O => \N__27335\,
            I => \sDAC_data_2_6_bm_1_4_cascade_\
        );

    \I__4081\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27329\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__27329\,
            I => \N__27326\
        );

    \I__4079\ : Span4Mux_v
    port map (
            O => \N__27326\,
            I => \N__27323\
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__27323\,
            I => \sDAC_mem_42Z0Z_1\
        );

    \I__4077\ : InMux
    port map (
            O => \N__27320\,
            I => \N__27317\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__27317\,
            I => \N__27314\
        );

    \I__4075\ : Span4Mux_v
    port map (
            O => \N__27314\,
            I => \N__27311\
        );

    \I__4074\ : Odrv4
    port map (
            O => \N__27311\,
            I => \sDAC_mem_10Z0Z_1\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__27308\,
            I => \sDAC_data_RNO_17Z0Z_4_cascade_\
        );

    \I__4072\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27302\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__27302\,
            I => \N__27299\
        );

    \I__4070\ : Span4Mux_h
    port map (
            O => \N__27299\,
            I => \N__27296\
        );

    \I__4069\ : Span4Mux_h
    port map (
            O => \N__27296\,
            I => \N__27293\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__27293\,
            I => \sDAC_mem_11Z0Z_1\
        );

    \I__4067\ : InMux
    port map (
            O => \N__27290\,
            I => \N__27287\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__27287\,
            I => \N__27284\
        );

    \I__4065\ : Span4Mux_v
    port map (
            O => \N__27284\,
            I => \N__27281\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__27281\,
            I => \sDAC_mem_42Z0Z_5\
        );

    \I__4063\ : InMux
    port map (
            O => \N__27278\,
            I => \N__27275\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__27275\,
            I => \N__27272\
        );

    \I__4061\ : Span4Mux_v
    port map (
            O => \N__27272\,
            I => \N__27269\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__27269\,
            I => \sDAC_mem_10Z0Z_5\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__27266\,
            I => \sDAC_data_RNO_17Z0Z_8_cascade_\
        );

    \I__4058\ : InMux
    port map (
            O => \N__27263\,
            I => \N__27260\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__27260\,
            I => \N__27257\
        );

    \I__4056\ : Odrv12
    port map (
            O => \N__27257\,
            I => \sDAC_mem_11Z0Z_5\
        );

    \I__4055\ : InMux
    port map (
            O => \N__27254\,
            I => \N__27251\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__27251\,
            I => \N__27248\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__27248\,
            I => \sDAC_mem_40Z0Z_5\
        );

    \I__4052\ : InMux
    port map (
            O => \N__27245\,
            I => \N__27242\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__27242\,
            I => \N__27239\
        );

    \I__4050\ : Odrv4
    port map (
            O => \N__27239\,
            I => \sDAC_mem_8Z0Z_5\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__27236\,
            I => \sDAC_data_2_20_am_1_8_cascade_\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__27233\,
            I => \sDAC_data_RNO_7Z0Z_8_cascade_\
        );

    \I__4047\ : InMux
    port map (
            O => \N__27230\,
            I => \N__27227\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__27227\,
            I => \sDAC_data_RNO_8Z0Z_8\
        );

    \I__4045\ : InMux
    port map (
            O => \N__27224\,
            I => \N__27221\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__27221\,
            I => \sDAC_data_RNO_15Z0Z_8\
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__27218\,
            I => \sDAC_data_2_14_ns_1_8_cascade_\
        );

    \I__4042\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__27212\,
            I => \sDAC_data_RNO_2Z0Z_8\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__27209\,
            I => \sDAC_data_RNO_1Z0Z_8_cascade_\
        );

    \I__4039\ : CascadeMux
    port map (
            O => \N__27206\,
            I => \sDAC_data_2_32_ns_1_6_cascade_\
        );

    \I__4038\ : InMux
    port map (
            O => \N__27203\,
            I => \N__27200\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__27200\,
            I => \sDAC_data_RNO_15Z0Z_6\
        );

    \I__4036\ : CascadeMux
    port map (
            O => \N__27197\,
            I => \sDAC_data_2_14_ns_1_6_cascade_\
        );

    \I__4035\ : InMux
    port map (
            O => \N__27194\,
            I => \N__27191\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__27191\,
            I => \sDAC_data_RNO_10Z0Z_6\
        );

    \I__4033\ : InMux
    port map (
            O => \N__27188\,
            I => \N__27185\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__27185\,
            I => \sDAC_data_RNO_2Z0Z_6\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__27182\,
            I => \sDAC_data_2_41_ns_1_6_cascade_\
        );

    \I__4030\ : InMux
    port map (
            O => \N__27179\,
            I => \N__27176\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__27176\,
            I => \sDAC_data_RNO_1Z0Z_6\
        );

    \I__4028\ : CascadeMux
    port map (
            O => \N__27173\,
            I => \sDAC_data_2_6_cascade_\
        );

    \I__4027\ : InMux
    port map (
            O => \N__27170\,
            I => \N__27167\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__27167\,
            I => \N__27164\
        );

    \I__4025\ : Odrv12
    port map (
            O => \N__27164\,
            I => \sDAC_dataZ0Z_6\
        );

    \I__4024\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27158\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__27158\,
            I => \N__27155\
        );

    \I__4022\ : Span4Mux_h
    port map (
            O => \N__27155\,
            I => \N__27152\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__27152\,
            I => \sDAC_mem_34Z0Z_5\
        );

    \I__4020\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27146\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__27146\,
            I => \sDAC_mem_2Z0Z_5\
        );

    \I__4018\ : InMux
    port map (
            O => \N__27143\,
            I => \N__27140\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__27140\,
            I => \N__27137\
        );

    \I__4016\ : Odrv12
    port map (
            O => \N__27137\,
            I => \sDAC_mem_35Z0Z_5\
        );

    \I__4015\ : CascadeMux
    port map (
            O => \N__27134\,
            I => \sDAC_data_2_6_bm_1_8_cascade_\
        );

    \I__4014\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27128\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__27128\,
            I => \sDAC_mem_3Z0Z_5\
        );

    \I__4012\ : CEMux
    port map (
            O => \N__27125\,
            I => \N__27122\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__27122\,
            I => \N__27119\
        );

    \I__4010\ : Odrv12
    port map (
            O => \N__27119\,
            I => \sDAC_mem_40_1_sqmuxa\
        );

    \I__4009\ : CEMux
    port map (
            O => \N__27116\,
            I => \N__27113\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__27113\,
            I => \sDAC_mem_8_1_sqmuxa\
        );

    \I__4007\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27107\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__27107\,
            I => \N__27103\
        );

    \I__4005\ : InMux
    port map (
            O => \N__27106\,
            I => \N__27100\
        );

    \I__4004\ : Span4Mux_h
    port map (
            O => \N__27103\,
            I => \N__27095\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__27100\,
            I => \N__27095\
        );

    \I__4002\ : Span4Mux_h
    port map (
            O => \N__27095\,
            I => \N__27087\
        );

    \I__4001\ : InMux
    port map (
            O => \N__27094\,
            I => \N__27084\
        );

    \I__4000\ : InMux
    port map (
            O => \N__27093\,
            I => \N__27081\
        );

    \I__3999\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27078\
        );

    \I__3998\ : InMux
    port map (
            O => \N__27091\,
            I => \N__27073\
        );

    \I__3997\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27073\
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__27087\,
            I => \N_317\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__27084\,
            I => \N_317\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__27081\,
            I => \N_317\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__27078\,
            I => \N_317\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__27073\,
            I => \N_317\
        );

    \I__3991\ : InMux
    port map (
            O => \N__27062\,
            I => \N__27058\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__27061\,
            I => \N__27054\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__27058\,
            I => \N__27051\
        );

    \I__3988\ : InMux
    port map (
            O => \N__27057\,
            I => \N__27046\
        );

    \I__3987\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27046\
        );

    \I__3986\ : Span4Mux_v
    port map (
            O => \N__27051\,
            I => \N__27043\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__27046\,
            I => \N__27040\
        );

    \I__3984\ : Span4Mux_v
    port map (
            O => \N__27043\,
            I => \N__27037\
        );

    \I__3983\ : Span4Mux_h
    port map (
            O => \N__27040\,
            I => \N__27034\
        );

    \I__3982\ : Span4Mux_v
    port map (
            O => \N__27037\,
            I => \N__27031\
        );

    \I__3981\ : Span4Mux_v
    port map (
            O => \N__27034\,
            I => \N__27028\
        );

    \I__3980\ : Odrv4
    port map (
            O => \N__27031\,
            I => \sAddress_RNI6VH7_4Z0Z_1\
        );

    \I__3979\ : Odrv4
    port map (
            O => \N__27028\,
            I => \sAddress_RNI6VH7_4Z0Z_1\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__27023\,
            I => \N__27016\
        );

    \I__3977\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27006\
        );

    \I__3976\ : InMux
    port map (
            O => \N__27021\,
            I => \N__27006\
        );

    \I__3975\ : InMux
    port map (
            O => \N__27020\,
            I => \N__27006\
        );

    \I__3974\ : InMux
    port map (
            O => \N__27019\,
            I => \N__27006\
        );

    \I__3973\ : InMux
    port map (
            O => \N__27016\,
            I => \N__27003\
        );

    \I__3972\ : InMux
    port map (
            O => \N__27015\,
            I => \N__27000\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__27006\,
            I => \N__26997\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__27003\,
            I => \N__26992\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__27000\,
            I => \N__26992\
        );

    \I__3968\ : Span12Mux_v
    port map (
            O => \N__26997\,
            I => \N__26989\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__26992\,
            I => \sAddress_RNI70I7Z0Z_1\
        );

    \I__3966\ : Odrv12
    port map (
            O => \N__26989\,
            I => \sAddress_RNI70I7Z0Z_1\
        );

    \I__3965\ : InMux
    port map (
            O => \N__26984\,
            I => \N__26981\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__26981\,
            I => \N__26978\
        );

    \I__3963\ : Span4Mux_h
    port map (
            O => \N__26978\,
            I => \N__26974\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__26977\,
            I => \N__26971\
        );

    \I__3961\ : Span4Mux_v
    port map (
            O => \N__26974\,
            I => \N__26968\
        );

    \I__3960\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26965\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__26968\,
            I => \sAddress_RNIAM2A_0Z0Z_1\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__26965\,
            I => \sAddress_RNIAM2A_0Z0Z_1\
        );

    \I__3957\ : InMux
    port map (
            O => \N__26960\,
            I => \N__26957\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__26957\,
            I => \N__26954\
        );

    \I__3955\ : Span4Mux_v
    port map (
            O => \N__26954\,
            I => \N__26951\
        );

    \I__3954\ : Span4Mux_h
    port map (
            O => \N__26951\,
            I => \N__26946\
        );

    \I__3953\ : InMux
    port map (
            O => \N__26950\,
            I => \N__26943\
        );

    \I__3952\ : InMux
    port map (
            O => \N__26949\,
            I => \N__26940\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__26946\,
            I => \sTrigCounterZ0Z_1\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__26943\,
            I => \sTrigCounterZ0Z_1\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__26940\,
            I => \sTrigCounterZ0Z_1\
        );

    \I__3948\ : IoInMux
    port map (
            O => \N__26933\,
            I => \N__26930\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__26930\,
            I => \N__26927\
        );

    \I__3946\ : Span4Mux_s2_h
    port map (
            O => \N__26927\,
            I => \N__26924\
        );

    \I__3945\ : Span4Mux_h
    port map (
            O => \N__26924\,
            I => \N__26921\
        );

    \I__3944\ : Sp12to4
    port map (
            O => \N__26921\,
            I => \N__26918\
        );

    \I__3943\ : Span12Mux_v
    port map (
            O => \N__26918\,
            I => \N__26915\
        );

    \I__3942\ : Odrv12
    port map (
            O => \N__26915\,
            I => \RAM_DATA_1Z0Z_14\
        );

    \I__3941\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26909\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__26909\,
            I => \N__26906\
        );

    \I__3939\ : Span4Mux_v
    port map (
            O => \N__26906\,
            I => \N__26903\
        );

    \I__3938\ : Sp12to4
    port map (
            O => \N__26903\,
            I => \N__26900\
        );

    \I__3937\ : Span12Mux_h
    port map (
            O => \N__26900\,
            I => \N__26897\
        );

    \I__3936\ : Odrv12
    port map (
            O => \N__26897\,
            I => \ADC2_c\
        );

    \I__3935\ : IoInMux
    port map (
            O => \N__26894\,
            I => \N__26891\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__26891\,
            I => \N__26888\
        );

    \I__3933\ : Span12Mux_s8_v
    port map (
            O => \N__26888\,
            I => \N__26885\
        );

    \I__3932\ : Span12Mux_h
    port map (
            O => \N__26885\,
            I => \N__26882\
        );

    \I__3931\ : Odrv12
    port map (
            O => \N__26882\,
            I => \RAM_DATA_1Z0Z_2\
        );

    \I__3930\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26876\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__26876\,
            I => \N__26873\
        );

    \I__3928\ : Span4Mux_v
    port map (
            O => \N__26873\,
            I => \N__26870\
        );

    \I__3927\ : Sp12to4
    port map (
            O => \N__26870\,
            I => \N__26867\
        );

    \I__3926\ : Span12Mux_h
    port map (
            O => \N__26867\,
            I => \N__26864\
        );

    \I__3925\ : Odrv12
    port map (
            O => \N__26864\,
            I => \ADC6_c\
        );

    \I__3924\ : IoInMux
    port map (
            O => \N__26861\,
            I => \N__26858\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__26858\,
            I => \N__26855\
        );

    \I__3922\ : Span4Mux_s2_v
    port map (
            O => \N__26855\,
            I => \N__26852\
        );

    \I__3921\ : Span4Mux_h
    port map (
            O => \N__26852\,
            I => \N__26849\
        );

    \I__3920\ : Span4Mux_v
    port map (
            O => \N__26849\,
            I => \N__26846\
        );

    \I__3919\ : Sp12to4
    port map (
            O => \N__26846\,
            I => \N__26843\
        );

    \I__3918\ : Odrv12
    port map (
            O => \N__26843\,
            I => \RAM_DATA_1Z0Z_6\
        );

    \I__3917\ : InMux
    port map (
            O => \N__26840\,
            I => \N__26837\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__26837\,
            I => \N__26834\
        );

    \I__3915\ : Span4Mux_v
    port map (
            O => \N__26834\,
            I => \N__26831\
        );

    \I__3914\ : Span4Mux_h
    port map (
            O => \N__26831\,
            I => \N__26828\
        );

    \I__3913\ : Span4Mux_h
    port map (
            O => \N__26828\,
            I => \N__26825\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__26825\,
            I => \ADC0_c\
        );

    \I__3911\ : IoInMux
    port map (
            O => \N__26822\,
            I => \N__26819\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__26819\,
            I => \N__26816\
        );

    \I__3909\ : Span4Mux_s2_v
    port map (
            O => \N__26816\,
            I => \N__26813\
        );

    \I__3908\ : Span4Mux_v
    port map (
            O => \N__26813\,
            I => \N__26810\
        );

    \I__3907\ : Sp12to4
    port map (
            O => \N__26810\,
            I => \N__26807\
        );

    \I__3906\ : Odrv12
    port map (
            O => \N__26807\,
            I => \RAM_DATA_1Z0Z_0\
        );

    \I__3905\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26801\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__26801\,
            I => \N__26798\
        );

    \I__3903\ : Odrv4
    port map (
            O => \N__26798\,
            I => \sDAC_mem_40Z0Z_3\
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__26795\,
            I => \N__26792\
        );

    \I__3901\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26789\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__26789\,
            I => \N__26786\
        );

    \I__3899\ : Span12Mux_v
    port map (
            O => \N__26786\,
            I => \N__26783\
        );

    \I__3898\ : Odrv12
    port map (
            O => \N__26783\,
            I => \sEEPoffZ0Z_15\
        );

    \I__3897\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26777\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__3895\ : Span4Mux_v
    port map (
            O => \N__26774\,
            I => \N__26771\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__26771\,
            I => \sEEPoffZ0Z_8\
        );

    \I__3893\ : CascadeMux
    port map (
            O => \N__26768\,
            I => \N__26765\
        );

    \I__3892\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26762\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__26762\,
            I => \N__26759\
        );

    \I__3890\ : Odrv12
    port map (
            O => \N__26759\,
            I => \sEEPoffZ0Z_9\
        );

    \I__3889\ : CEMux
    port map (
            O => \N__26756\,
            I => \N__26752\
        );

    \I__3888\ : CEMux
    port map (
            O => \N__26755\,
            I => \N__26749\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__26752\,
            I => \sAddress_RNIA6242_2Z0Z_0\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__26749\,
            I => \sAddress_RNIA6242_2Z0Z_0\
        );

    \I__3885\ : IoInMux
    port map (
            O => \N__26744\,
            I => \N__26741\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__26741\,
            I => \N__26738\
        );

    \I__3883\ : IoSpan4Mux
    port map (
            O => \N__26738\,
            I => \N__26735\
        );

    \I__3882\ : Span4Mux_s3_h
    port map (
            O => \N__26735\,
            I => \N__26732\
        );

    \I__3881\ : Span4Mux_h
    port map (
            O => \N__26732\,
            I => \N__26729\
        );

    \I__3880\ : Span4Mux_h
    port map (
            O => \N__26729\,
            I => \N__26726\
        );

    \I__3879\ : Span4Mux_h
    port map (
            O => \N__26726\,
            I => \N__26723\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__26723\,
            I => \un4_sacqtime_cry_23_c_RNI2CQMZ0\
        );

    \I__3877\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26717\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__26717\,
            I => \N__26714\
        );

    \I__3875\ : Span4Mux_v
    port map (
            O => \N__26714\,
            I => \N__26711\
        );

    \I__3874\ : Sp12to4
    port map (
            O => \N__26711\,
            I => \N__26708\
        );

    \I__3873\ : Span12Mux_h
    port map (
            O => \N__26708\,
            I => \N__26705\
        );

    \I__3872\ : Odrv12
    port map (
            O => \N__26705\,
            I => \ADC5_c\
        );

    \I__3871\ : IoInMux
    port map (
            O => \N__26702\,
            I => \N__26699\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__26699\,
            I => \N__26696\
        );

    \I__3869\ : IoSpan4Mux
    port map (
            O => \N__26696\,
            I => \N__26693\
        );

    \I__3868\ : IoSpan4Mux
    port map (
            O => \N__26693\,
            I => \N__26690\
        );

    \I__3867\ : Span4Mux_s2_v
    port map (
            O => \N__26690\,
            I => \N__26687\
        );

    \I__3866\ : Sp12to4
    port map (
            O => \N__26687\,
            I => \N__26684\
        );

    \I__3865\ : Span12Mux_s8_v
    port map (
            O => \N__26684\,
            I => \N__26681\
        );

    \I__3864\ : Odrv12
    port map (
            O => \N__26681\,
            I => \RAM_DATA_1Z0Z_5\
        );

    \I__3863\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26675\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__26675\,
            I => \N__26672\
        );

    \I__3861\ : Span4Mux_v
    port map (
            O => \N__26672\,
            I => \N__26669\
        );

    \I__3860\ : Sp12to4
    port map (
            O => \N__26669\,
            I => \N__26666\
        );

    \I__3859\ : Span12Mux_h
    port map (
            O => \N__26666\,
            I => \N__26663\
        );

    \I__3858\ : Odrv12
    port map (
            O => \N__26663\,
            I => \ADC1_c\
        );

    \I__3857\ : IoInMux
    port map (
            O => \N__26660\,
            I => \N__26657\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__26657\,
            I => \N__26654\
        );

    \I__3855\ : Span12Mux_s11_v
    port map (
            O => \N__26654\,
            I => \N__26651\
        );

    \I__3854\ : Span12Mux_h
    port map (
            O => \N__26651\,
            I => \N__26648\
        );

    \I__3853\ : Odrv12
    port map (
            O => \N__26648\,
            I => \RAM_DATA_1Z0Z_1\
        );

    \I__3852\ : InMux
    port map (
            O => \N__26645\,
            I => \N__26642\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__26642\,
            I => \N__26639\
        );

    \I__3850\ : Span4Mux_v
    port map (
            O => \N__26639\,
            I => \N__26636\
        );

    \I__3849\ : Sp12to4
    port map (
            O => \N__26636\,
            I => \N__26633\
        );

    \I__3848\ : Span12Mux_h
    port map (
            O => \N__26633\,
            I => \N__26630\
        );

    \I__3847\ : Odrv12
    port map (
            O => \N__26630\,
            I => \ADC9_c\
        );

    \I__3846\ : IoInMux
    port map (
            O => \N__26627\,
            I => \N__26624\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__26624\,
            I => \N__26621\
        );

    \I__3844\ : Span12Mux_s4_h
    port map (
            O => \N__26621\,
            I => \N__26618\
        );

    \I__3843\ : Span12Mux_v
    port map (
            O => \N__26618\,
            I => \N__26615\
        );

    \I__3842\ : Span12Mux_h
    port map (
            O => \N__26615\,
            I => \N__26612\
        );

    \I__3841\ : Odrv12
    port map (
            O => \N__26612\,
            I => \RAM_DATA_1Z0Z_10\
        );

    \I__3840\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26606\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__26606\,
            I => \N__26603\
        );

    \I__3838\ : Span12Mux_v
    port map (
            O => \N__26603\,
            I => \N__26600\
        );

    \I__3837\ : Span12Mux_h
    port map (
            O => \N__26600\,
            I => \N__26597\
        );

    \I__3836\ : Odrv12
    port map (
            O => \N__26597\,
            I => top_tour1_c
        );

    \I__3835\ : IoInMux
    port map (
            O => \N__26594\,
            I => \N__26591\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26588\
        );

    \I__3833\ : IoSpan4Mux
    port map (
            O => \N__26588\,
            I => \N__26585\
        );

    \I__3832\ : Span4Mux_s2_h
    port map (
            O => \N__26585\,
            I => \N__26582\
        );

    \I__3831\ : Sp12to4
    port map (
            O => \N__26582\,
            I => \N__26579\
        );

    \I__3830\ : Span12Mux_h
    port map (
            O => \N__26579\,
            I => \N__26576\
        );

    \I__3829\ : Odrv12
    port map (
            O => \N__26576\,
            I => \RAM_DATA_1Z0Z_11\
        );

    \I__3828\ : InMux
    port map (
            O => \N__26573\,
            I => \N__26570\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__26570\,
            I => \N__26567\
        );

    \I__3826\ : Span4Mux_v
    port map (
            O => \N__26567\,
            I => \N__26564\
        );

    \I__3825\ : Span4Mux_h
    port map (
            O => \N__26564\,
            I => \N__26559\
        );

    \I__3824\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26556\
        );

    \I__3823\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26553\
        );

    \I__3822\ : Odrv4
    port map (
            O => \N__26559\,
            I => \sTrigCounterZ0Z_0\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__26556\,
            I => \sTrigCounterZ0Z_0\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__26553\,
            I => \sTrigCounterZ0Z_0\
        );

    \I__3819\ : IoInMux
    port map (
            O => \N__26546\,
            I => \N__26543\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__26543\,
            I => \N__26540\
        );

    \I__3817\ : IoSpan4Mux
    port map (
            O => \N__26540\,
            I => \N__26537\
        );

    \I__3816\ : Span4Mux_s2_h
    port map (
            O => \N__26537\,
            I => \N__26534\
        );

    \I__3815\ : Sp12to4
    port map (
            O => \N__26534\,
            I => \N__26531\
        );

    \I__3814\ : Span12Mux_h
    port map (
            O => \N__26531\,
            I => \N__26528\
        );

    \I__3813\ : Odrv12
    port map (
            O => \N__26528\,
            I => \RAM_DATA_1Z0Z_13\
        );

    \I__3812\ : CEMux
    port map (
            O => \N__26525\,
            I => \N__26522\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__26522\,
            I => \N__26519\
        );

    \I__3810\ : Odrv12
    port map (
            O => \N__26519\,
            I => \sAddress_RNIA6242_0Z0Z_0\
        );

    \I__3809\ : InMux
    port map (
            O => \N__26516\,
            I => \N__26513\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__26513\,
            I => \N__26510\
        );

    \I__3807\ : Span4Mux_v
    port map (
            O => \N__26510\,
            I => \N__26507\
        );

    \I__3806\ : Odrv4
    port map (
            O => \N__26507\,
            I => \sEEPoffZ0Z_11\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__26504\,
            I => \N__26501\
        );

    \I__3804\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26498\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__26498\,
            I => \N__26495\
        );

    \I__3802\ : Odrv12
    port map (
            O => \N__26495\,
            I => \sEEPoffZ0Z_12\
        );

    \I__3801\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26489\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__26489\,
            I => \N__26486\
        );

    \I__3799\ : Span4Mux_v
    port map (
            O => \N__26486\,
            I => \N__26483\
        );

    \I__3798\ : Odrv4
    port map (
            O => \N__26483\,
            I => \sEEPoffZ0Z_13\
        );

    \I__3797\ : InMux
    port map (
            O => \N__26480\,
            I => \N__26477\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__26477\,
            I => \N__26474\
        );

    \I__3795\ : Odrv12
    port map (
            O => \N__26474\,
            I => \sEEPoffZ0Z_14\
        );

    \I__3794\ : CEMux
    port map (
            O => \N__26471\,
            I => \N__26468\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__26468\,
            I => \N__26465\
        );

    \I__3792\ : Span4Mux_v
    port map (
            O => \N__26465\,
            I => \N__26462\
        );

    \I__3791\ : Span4Mux_h
    port map (
            O => \N__26462\,
            I => \N__26459\
        );

    \I__3790\ : Odrv4
    port map (
            O => \N__26459\,
            I => \sAddress_RNIA6242_1Z0Z_0\
        );

    \I__3789\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26453\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__26453\,
            I => \sCounter_i_19\
        );

    \I__3787\ : InMux
    port map (
            O => \N__26450\,
            I => \N__26447\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__26447\,
            I => \sCounter_i_20\
        );

    \I__3785\ : InMux
    port map (
            O => \N__26444\,
            I => \N__26441\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__26441\,
            I => \sCounter_i_21\
        );

    \I__3783\ : InMux
    port map (
            O => \N__26438\,
            I => \N__26435\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__26435\,
            I => \sCounter_i_22\
        );

    \I__3781\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26429\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__26429\,
            I => \sCounter_i_23\
        );

    \I__3779\ : InMux
    port map (
            O => \N__26426\,
            I => \bfn_12_13_0_\
        );

    \I__3778\ : IoInMux
    port map (
            O => \N__26423\,
            I => \N__26420\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__3776\ : IoSpan4Mux
    port map (
            O => \N__26417\,
            I => \N__26414\
        );

    \I__3775\ : Span4Mux_s1_h
    port map (
            O => \N__26414\,
            I => \N__26411\
        );

    \I__3774\ : Span4Mux_h
    port map (
            O => \N__26411\,
            I => \N__26408\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__26408\,
            I => \N__26405\
        );

    \I__3772\ : Span4Mux_h
    port map (
            O => \N__26405\,
            I => \N__26402\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__26402\,
            I => \N_1683_i\
        );

    \I__3770\ : InMux
    port map (
            O => \N__26399\,
            I => \N__26396\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__26396\,
            I => \N__26393\
        );

    \I__3768\ : Span4Mux_v
    port map (
            O => \N__26393\,
            I => \N__26390\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__26390\,
            I => \N__26386\
        );

    \I__3766\ : CascadeMux
    port map (
            O => \N__26389\,
            I => \N__26383\
        );

    \I__3765\ : Span4Mux_h
    port map (
            O => \N__26386\,
            I => \N__26380\
        );

    \I__3764\ : InMux
    port map (
            O => \N__26383\,
            I => \N__26377\
        );

    \I__3763\ : Odrv4
    port map (
            O => \N__26380\,
            I => \sbuttonModeStatusZ0\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__26377\,
            I => \sbuttonModeStatusZ0\
        );

    \I__3761\ : InMux
    port map (
            O => \N__26372\,
            I => \N__26369\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__3759\ : Odrv4
    port map (
            O => \N__26366\,
            I => \sbuttonModeStatus_0_sqmuxa_0\
        );

    \I__3758\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26360\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__26360\,
            I => \sbuttonModeStatus_0_sqmuxa_18\
        );

    \I__3756\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26354\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__26354\,
            I => \sCounter_i_16\
        );

    \I__3754\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26348\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__26348\,
            I => \sCounter_i_17\
        );

    \I__3752\ : InMux
    port map (
            O => \N__26345\,
            I => \N__26342\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__26342\,
            I => \sCounter_i_18\
        );

    \I__3750\ : InMux
    port map (
            O => \N__26339\,
            I => \N__26336\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__26336\,
            I => \N__26333\
        );

    \I__3748\ : Span4Mux_v
    port map (
            O => \N__26333\,
            I => \N__26330\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__26330\,
            I => \sEEPoffZ0Z_2\
        );

    \I__3746\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26324\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__26324\,
            I => \N__26321\
        );

    \I__3744\ : Span4Mux_v
    port map (
            O => \N__26321\,
            I => \N__26318\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__26318\,
            I => \sEEPoffZ0Z_3\
        );

    \I__3742\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__26312\,
            I => \N__26309\
        );

    \I__3740\ : Span4Mux_v
    port map (
            O => \N__26309\,
            I => \N__26306\
        );

    \I__3739\ : Odrv4
    port map (
            O => \N__26306\,
            I => \sEEPoffZ0Z_4\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__26303\,
            I => \N__26300\
        );

    \I__3737\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26297\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__26297\,
            I => \N__26294\
        );

    \I__3735\ : Span4Mux_v
    port map (
            O => \N__26294\,
            I => \N__26291\
        );

    \I__3734\ : Odrv4
    port map (
            O => \N__26291\,
            I => \sEEPoffZ0Z_5\
        );

    \I__3733\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26285\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__26285\,
            I => \N__26282\
        );

    \I__3731\ : Span4Mux_v
    port map (
            O => \N__26282\,
            I => \N__26279\
        );

    \I__3730\ : Odrv4
    port map (
            O => \N__26279\,
            I => \sEEPoffZ0Z_6\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__26276\,
            I => \N__26273\
        );

    \I__3728\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26270\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__26270\,
            I => \N__26267\
        );

    \I__3726\ : Span4Mux_v
    port map (
            O => \N__26267\,
            I => \N__26264\
        );

    \I__3725\ : Odrv4
    port map (
            O => \N__26264\,
            I => \sEEPoffZ0Z_7\
        );

    \I__3724\ : InMux
    port map (
            O => \N__26261\,
            I => \N__26258\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__26258\,
            I => \N__26255\
        );

    \I__3722\ : Span4Mux_v
    port map (
            O => \N__26255\,
            I => \N__26252\
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__26252\,
            I => \sEEPoffZ0Z_10\
        );

    \I__3720\ : InMux
    port map (
            O => \N__26249\,
            I => \N__26246\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__26246\,
            I => \N__26243\
        );

    \I__3718\ : Odrv12
    port map (
            O => \N__26243\,
            I => \sDAC_mem_39Z0Z_1\
        );

    \I__3717\ : CEMux
    port map (
            O => \N__26240\,
            I => \N__26237\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__26237\,
            I => \N__26234\
        );

    \I__3715\ : Span4Mux_v
    port map (
            O => \N__26234\,
            I => \N__26231\
        );

    \I__3714\ : Span4Mux_h
    port map (
            O => \N__26231\,
            I => \N__26228\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__26228\,
            I => \sDAC_mem_39_1_sqmuxa\
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__26225\,
            I => \N__26222\
        );

    \I__3711\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26219\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__26219\,
            I => \N__26216\
        );

    \I__3709\ : Span4Mux_v
    port map (
            O => \N__26216\,
            I => \N__26213\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__26213\,
            I => \sEEPoffZ0Z_0\
        );

    \I__3707\ : InMux
    port map (
            O => \N__26210\,
            I => \N__26207\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__26207\,
            I => \N__26204\
        );

    \I__3705\ : Span4Mux_v
    port map (
            O => \N__26204\,
            I => \N__26201\
        );

    \I__3704\ : Odrv4
    port map (
            O => \N__26201\,
            I => \sEEPoffZ0Z_1\
        );

    \I__3703\ : InMux
    port map (
            O => \N__26198\,
            I => \N__26188\
        );

    \I__3702\ : InMux
    port map (
            O => \N__26197\,
            I => \N__26188\
        );

    \I__3701\ : InMux
    port map (
            O => \N__26196\,
            I => \N__26185\
        );

    \I__3700\ : InMux
    port map (
            O => \N__26195\,
            I => \N__26179\
        );

    \I__3699\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26179\
        );

    \I__3698\ : CascadeMux
    port map (
            O => \N__26193\,
            I => \N__26175\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__26188\,
            I => \N__26171\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__26185\,
            I => \N__26168\
        );

    \I__3695\ : CascadeMux
    port map (
            O => \N__26184\,
            I => \N__26159\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__26179\,
            I => \N__26156\
        );

    \I__3693\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26153\
        );

    \I__3692\ : InMux
    port map (
            O => \N__26175\,
            I => \N__26148\
        );

    \I__3691\ : InMux
    port map (
            O => \N__26174\,
            I => \N__26148\
        );

    \I__3690\ : Span12Mux_s11_h
    port map (
            O => \N__26171\,
            I => \N__26145\
        );

    \I__3689\ : Span4Mux_v
    port map (
            O => \N__26168\,
            I => \N__26142\
        );

    \I__3688\ : InMux
    port map (
            O => \N__26167\,
            I => \N__26137\
        );

    \I__3687\ : InMux
    port map (
            O => \N__26166\,
            I => \N__26137\
        );

    \I__3686\ : InMux
    port map (
            O => \N__26165\,
            I => \N__26134\
        );

    \I__3685\ : InMux
    port map (
            O => \N__26164\,
            I => \N__26131\
        );

    \I__3684\ : InMux
    port map (
            O => \N__26163\,
            I => \N__26124\
        );

    \I__3683\ : InMux
    port map (
            O => \N__26162\,
            I => \N__26124\
        );

    \I__3682\ : InMux
    port map (
            O => \N__26159\,
            I => \N__26124\
        );

    \I__3681\ : Span4Mux_v
    port map (
            O => \N__26156\,
            I => \N__26121\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__26153\,
            I => \N__26118\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__26148\,
            I => \sPointerZ0Z_1\
        );

    \I__3678\ : Odrv12
    port map (
            O => \N__26145\,
            I => \sPointerZ0Z_1\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__26142\,
            I => \sPointerZ0Z_1\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__26137\,
            I => \sPointerZ0Z_1\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__26134\,
            I => \sPointerZ0Z_1\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__26131\,
            I => \sPointerZ0Z_1\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__26124\,
            I => \sPointerZ0Z_1\
        );

    \I__3672\ : Odrv4
    port map (
            O => \N__26121\,
            I => \sPointerZ0Z_1\
        );

    \I__3671\ : Odrv4
    port map (
            O => \N__26118\,
            I => \sPointerZ0Z_1\
        );

    \I__3670\ : InMux
    port map (
            O => \N__26099\,
            I => \N__26095\
        );

    \I__3669\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26092\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__26095\,
            I => \N__26084\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__26092\,
            I => \N__26081\
        );

    \I__3666\ : InMux
    port map (
            O => \N__26091\,
            I => \N__26078\
        );

    \I__3665\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26073\
        );

    \I__3664\ : InMux
    port map (
            O => \N__26089\,
            I => \N__26073\
        );

    \I__3663\ : InMux
    port map (
            O => \N__26088\,
            I => \N__26068\
        );

    \I__3662\ : InMux
    port map (
            O => \N__26087\,
            I => \N__26068\
        );

    \I__3661\ : Span4Mux_h
    port map (
            O => \N__26084\,
            I => \N__26065\
        );

    \I__3660\ : Span4Mux_v
    port map (
            O => \N__26081\,
            I => \N__26062\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__26078\,
            I => \N__26059\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__26073\,
            I => \sPointerZ0Z_0\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__26068\,
            I => \sPointerZ0Z_0\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__26065\,
            I => \sPointerZ0Z_0\
        );

    \I__3655\ : Odrv4
    port map (
            O => \N__26062\,
            I => \sPointerZ0Z_0\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__26059\,
            I => \sPointerZ0Z_0\
        );

    \I__3653\ : InMux
    port map (
            O => \N__26048\,
            I => \N__26045\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__26045\,
            I => \N__26038\
        );

    \I__3651\ : InMux
    port map (
            O => \N__26044\,
            I => \N__26031\
        );

    \I__3650\ : InMux
    port map (
            O => \N__26043\,
            I => \N__26031\
        );

    \I__3649\ : InMux
    port map (
            O => \N__26042\,
            I => \N__26031\
        );

    \I__3648\ : InMux
    port map (
            O => \N__26041\,
            I => \N__26028\
        );

    \I__3647\ : Span4Mux_v
    port map (
            O => \N__26038\,
            I => \N__26024\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__26031\,
            I => \N__26019\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__26028\,
            I => \N__26019\
        );

    \I__3644\ : InMux
    port map (
            O => \N__26027\,
            I => \N__26016\
        );

    \I__3643\ : Span4Mux_h
    port map (
            O => \N__26024\,
            I => \N__26009\
        );

    \I__3642\ : Span4Mux_v
    port map (
            O => \N__26019\,
            I => \N__26009\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__26016\,
            I => \N__26009\
        );

    \I__3640\ : Odrv4
    port map (
            O => \N__26009\,
            I => \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1\
        );

    \I__3639\ : InMux
    port map (
            O => \N__26006\,
            I => \N__26003\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__26003\,
            I => \N__26000\
        );

    \I__3637\ : Span4Mux_h
    port map (
            O => \N__26000\,
            I => \N__25997\
        );

    \I__3636\ : Span4Mux_h
    port map (
            O => \N__25997\,
            I => \N__25994\
        );

    \I__3635\ : Odrv4
    port map (
            O => \N__25994\,
            I => \N_1624\
        );

    \I__3634\ : InMux
    port map (
            O => \N__25991\,
            I => \N__25988\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__25988\,
            I => \N__25985\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__25985\,
            I => \sDAC_mem_34Z0Z_3\
        );

    \I__3631\ : CEMux
    port map (
            O => \N__25982\,
            I => \N__25979\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__25979\,
            I => \N__25976\
        );

    \I__3629\ : Span4Mux_h
    port map (
            O => \N__25976\,
            I => \N__25973\
        );

    \I__3628\ : Odrv4
    port map (
            O => \N__25973\,
            I => \sDAC_mem_34_1_sqmuxa\
        );

    \I__3627\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25967\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__25967\,
            I => \sDAC_mem_7Z0Z_1\
        );

    \I__3625\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25961\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__25961\,
            I => \N__25958\
        );

    \I__3623\ : Span4Mux_v
    port map (
            O => \N__25958\,
            I => \N__25955\
        );

    \I__3622\ : Odrv4
    port map (
            O => \N__25955\,
            I => un1_spointer11_2_0_0_a2_5
        );

    \I__3621\ : InMux
    port map (
            O => \N__25952\,
            I => \N__25949\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__25949\,
            I => \N__25946\
        );

    \I__3619\ : Span4Mux_h
    port map (
            O => \N__25946\,
            I => \N__25942\
        );

    \I__3618\ : InMux
    port map (
            O => \N__25945\,
            I => \N__25939\
        );

    \I__3617\ : Span4Mux_h
    port map (
            O => \N__25942\,
            I => \N__25936\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__25939\,
            I => \N__25933\
        );

    \I__3615\ : Odrv4
    port map (
            O => \N__25936\,
            I => \N_183\
        );

    \I__3614\ : Odrv12
    port map (
            O => \N__25933\,
            I => \N_183\
        );

    \I__3613\ : InMux
    port map (
            O => \N__25928\,
            I => \N__25925\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__25925\,
            I => \sDAC_mem_8Z0Z_3\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__25922\,
            I => \sDAC_data_2_20_am_1_6_cascade_\
        );

    \I__3610\ : InMux
    port map (
            O => \N__25919\,
            I => \N__25916\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__25916\,
            I => \N__25913\
        );

    \I__3608\ : Odrv4
    port map (
            O => \N__25913\,
            I => \sDAC_mem_10Z0Z_3\
        );

    \I__3607\ : InMux
    port map (
            O => \N__25910\,
            I => \N__25907\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__25907\,
            I => \N__25904\
        );

    \I__3605\ : Odrv12
    port map (
            O => \N__25904\,
            I => \sDAC_mem_42Z0Z_3\
        );

    \I__3604\ : CascadeMux
    port map (
            O => \N__25901\,
            I => \sDAC_data_RNO_17Z0Z_6_cascade_\
        );

    \I__3603\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25895\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__25895\,
            I => \N__25892\
        );

    \I__3601\ : Span4Mux_v
    port map (
            O => \N__25892\,
            I => \N__25889\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__25889\,
            I => \sDAC_mem_11Z0Z_3\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__25886\,
            I => \sDAC_data_RNO_8Z0Z_6_cascade_\
        );

    \I__3598\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25880\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__25880\,
            I => \sDAC_data_RNO_7Z0Z_6\
        );

    \I__3596\ : InMux
    port map (
            O => \N__25877\,
            I => \N__25874\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__25874\,
            I => \sDAC_mem_2Z0Z_3\
        );

    \I__3594\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25868\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__25868\,
            I => \N__25865\
        );

    \I__3592\ : Span12Mux_s11_v
    port map (
            O => \N__25865\,
            I => \N__25862\
        );

    \I__3591\ : Odrv12
    port map (
            O => \N__25862\,
            I => \sDAC_mem_35Z0Z_3\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__25859\,
            I => \sDAC_data_2_6_bm_1_6_cascade_\
        );

    \I__3589\ : InMux
    port map (
            O => \N__25856\,
            I => \N__25853\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__25853\,
            I => \sDAC_mem_3Z0Z_3\
        );

    \I__3587\ : InMux
    port map (
            O => \N__25850\,
            I => \N__25847\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__25847\,
            I => \N__25844\
        );

    \I__3585\ : Span4Mux_h
    port map (
            O => \N__25844\,
            I => \N__25841\
        );

    \I__3584\ : Span4Mux_v
    port map (
            O => \N__25841\,
            I => \N__25838\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__25838\,
            I => g0_4_0
        );

    \I__3582\ : InMux
    port map (
            O => \N__25835\,
            I => \bfn_11_20_0_\
        );

    \I__3581\ : InMux
    port map (
            O => \N__25832\,
            I => \N__25829\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__25829\,
            I => \N__25826\
        );

    \I__3579\ : Sp12to4
    port map (
            O => \N__25826\,
            I => \N__25823\
        );

    \I__3578\ : Span12Mux_h
    port map (
            O => \N__25823\,
            I => \N__25820\
        );

    \I__3577\ : Odrv12
    port map (
            O => \N__25820\,
            I => spi_sclk_ft_c
        );

    \I__3576\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25814\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__25814\,
            I => \N__25811\
        );

    \I__3574\ : Span4Mux_v
    port map (
            O => \N__25811\,
            I => \N__25808\
        );

    \I__3573\ : Sp12to4
    port map (
            O => \N__25808\,
            I => \N__25805\
        );

    \I__3572\ : Span12Mux_h
    port map (
            O => \N__25805\,
            I => \N__25802\
        );

    \I__3571\ : Odrv12
    port map (
            O => \N__25802\,
            I => spi_sclk_rpi_c
        );

    \I__3570\ : IoInMux
    port map (
            O => \N__25799\,
            I => \N__25796\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__25796\,
            I => \N__25793\
        );

    \I__3568\ : Odrv12
    port map (
            O => \N__25793\,
            I => spi_sclk
        );

    \I__3567\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25787\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__25787\,
            I => \N__25784\
        );

    \I__3565\ : Span4Mux_h
    port map (
            O => \N__25784\,
            I => \N__25781\
        );

    \I__3564\ : Odrv4
    port map (
            O => \N__25781\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3\
        );

    \I__3563\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25775\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__25775\,
            I => \N__25772\
        );

    \I__3561\ : Span4Mux_h
    port map (
            O => \N__25772\,
            I => \N__25769\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__25769\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_12\
        );

    \I__3559\ : InMux
    port map (
            O => \N__25766\,
            I => \N__25763\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__25763\,
            I => \N__25760\
        );

    \I__3557\ : Span4Mux_h
    port map (
            O => \N__25760\,
            I => \N__25757\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__25757\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12\
        );

    \I__3555\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25751\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__25751\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7\
        );

    \I__3553\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25745\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__25745\,
            I => \N__25742\
        );

    \I__3551\ : Odrv12
    port map (
            O => \N__25742\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9\
        );

    \I__3550\ : InMux
    port map (
            O => \N__25739\,
            I => \N__25736\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__25736\,
            I => \sEEDelayACQZ0Z_14\
        );

    \I__3548\ : InMux
    port map (
            O => \N__25733\,
            I => \N__25730\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__25730\,
            I => \sEEDelayACQ_i_14\
        );

    \I__3546\ : InMux
    port map (
            O => \N__25727\,
            I => \N__25724\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__25724\,
            I => \sEEDelayACQZ0Z_15\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__25721\,
            I => \N__25718\
        );

    \I__3543\ : InMux
    port map (
            O => \N__25718\,
            I => \N__25715\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__25715\,
            I => \sEEDelayACQ_i_15\
        );

    \I__3541\ : InMux
    port map (
            O => \N__25712\,
            I => \N__25709\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__25709\,
            I => \N__25706\
        );

    \I__3539\ : Span4Mux_h
    port map (
            O => \N__25706\,
            I => \N__25703\
        );

    \I__3538\ : Span4Mux_v
    port map (
            O => \N__25703\,
            I => \N__25700\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__25700\,
            I => g1_i_a4_4
        );

    \I__3536\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25694\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__25694\,
            I => \sEEDelayACQZ0Z_6\
        );

    \I__3534\ : InMux
    port map (
            O => \N__25691\,
            I => \N__25688\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__25688\,
            I => \sEEDelayACQ_i_6\
        );

    \I__3532\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25682\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__25682\,
            I => \sEEDelayACQZ0Z_7\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__25679\,
            I => \N__25676\
        );

    \I__3529\ : InMux
    port map (
            O => \N__25676\,
            I => \N__25673\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__25673\,
            I => \sEEDelayACQ_i_7\
        );

    \I__3527\ : InMux
    port map (
            O => \N__25670\,
            I => \N__25667\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__25667\,
            I => \sEEDelayACQZ0Z_8\
        );

    \I__3525\ : InMux
    port map (
            O => \N__25664\,
            I => \N__25661\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__25661\,
            I => \sEEDelayACQ_i_8\
        );

    \I__3523\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25655\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__25655\,
            I => \sEEDelayACQZ0Z_9\
        );

    \I__3521\ : InMux
    port map (
            O => \N__25652\,
            I => \N__25649\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__25649\,
            I => \sEEDelayACQ_i_9\
        );

    \I__3519\ : InMux
    port map (
            O => \N__25646\,
            I => \N__25643\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__25643\,
            I => \sEEDelayACQZ0Z_10\
        );

    \I__3517\ : InMux
    port map (
            O => \N__25640\,
            I => \N__25637\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__25637\,
            I => \sEEDelayACQ_i_10\
        );

    \I__3515\ : InMux
    port map (
            O => \N__25634\,
            I => \N__25631\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__25631\,
            I => \sEEDelayACQZ0Z_11\
        );

    \I__3513\ : InMux
    port map (
            O => \N__25628\,
            I => \N__25625\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__25625\,
            I => \sEEDelayACQ_i_11\
        );

    \I__3511\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25619\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__25619\,
            I => \sEEDelayACQZ0Z_12\
        );

    \I__3509\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25613\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__25613\,
            I => \sEEDelayACQ_i_12\
        );

    \I__3507\ : InMux
    port map (
            O => \N__25610\,
            I => \N__25607\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__25607\,
            I => \sEEDelayACQZ0Z_13\
        );

    \I__3505\ : InMux
    port map (
            O => \N__25604\,
            I => \N__25601\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__25601\,
            I => \sEEDelayACQ_i_13\
        );

    \I__3503\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25595\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__25595\,
            I => \sEEDelayACQZ0Z_0\
        );

    \I__3501\ : InMux
    port map (
            O => \N__25592\,
            I => \N__25589\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__25589\,
            I => \sEEDelayACQ_i_0\
        );

    \I__3499\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25583\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__25583\,
            I => \sEEDelayACQZ0Z_1\
        );

    \I__3497\ : InMux
    port map (
            O => \N__25580\,
            I => \N__25577\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__25577\,
            I => \sEEDelayACQ_i_1\
        );

    \I__3495\ : InMux
    port map (
            O => \N__25574\,
            I => \N__25571\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__25571\,
            I => \sEEDelayACQZ0Z_2\
        );

    \I__3493\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25565\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__25565\,
            I => \sEEDelayACQ_i_2\
        );

    \I__3491\ : InMux
    port map (
            O => \N__25562\,
            I => \N__25559\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__25559\,
            I => \sEEDelayACQZ0Z_3\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__25556\,
            I => \N__25553\
        );

    \I__3488\ : InMux
    port map (
            O => \N__25553\,
            I => \N__25550\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__25550\,
            I => \sEEDelayACQ_i_3\
        );

    \I__3486\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25544\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__25544\,
            I => \sEEDelayACQZ0Z_4\
        );

    \I__3484\ : InMux
    port map (
            O => \N__25541\,
            I => \N__25538\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__25538\,
            I => \sEEDelayACQ_i_4\
        );

    \I__3482\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25532\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__25532\,
            I => \sEEDelayACQZ0Z_5\
        );

    \I__3480\ : InMux
    port map (
            O => \N__25529\,
            I => \N__25526\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__25526\,
            I => \sEEDelayACQ_i_5\
        );

    \I__3478\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25517\
        );

    \I__3477\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25510\
        );

    \I__3476\ : InMux
    port map (
            O => \N__25521\,
            I => \N__25510\
        );

    \I__3475\ : InMux
    port map (
            O => \N__25520\,
            I => \N__25510\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__25517\,
            I => \N__25505\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__25510\,
            I => \N__25505\
        );

    \I__3472\ : Span4Mux_h
    port map (
            O => \N__25505\,
            I => \N__25502\
        );

    \I__3471\ : Span4Mux_v
    port map (
            O => \N__25502\,
            I => \N__25499\
        );

    \I__3470\ : Odrv4
    port map (
            O => \N__25499\,
            I => un1_spointer11_5_0_2
        );

    \I__3469\ : CEMux
    port map (
            O => \N__25496\,
            I => \N__25493\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__25493\,
            I => \sAddress_RNIA6242_3Z0Z_0\
        );

    \I__3467\ : InMux
    port map (
            O => \N__25490\,
            I => \N__25486\
        );

    \I__3466\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25483\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__25486\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__25483\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2\
        );

    \I__3463\ : InMux
    port map (
            O => \N__25478\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1\
        );

    \I__3462\ : InMux
    port map (
            O => \N__25475\,
            I => \N__25471\
        );

    \I__3461\ : InMux
    port map (
            O => \N__25474\,
            I => \N__25468\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__25471\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__25468\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3\
        );

    \I__3458\ : InMux
    port map (
            O => \N__25463\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2\
        );

    \I__3457\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25457\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__25457\,
            I => \N__25454\
        );

    \I__3455\ : Span4Mux_h
    port map (
            O => \N__25454\,
            I => \N__25450\
        );

    \I__3454\ : InMux
    port map (
            O => \N__25453\,
            I => \N__25447\
        );

    \I__3453\ : Span4Mux_h
    port map (
            O => \N__25450\,
            I => \N__25444\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__25447\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4\
        );

    \I__3451\ : Odrv4
    port map (
            O => \N__25444\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4\
        );

    \I__3450\ : InMux
    port map (
            O => \N__25439\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__25436\,
            I => \N__25432\
        );

    \I__3448\ : InMux
    port map (
            O => \N__25435\,
            I => \N__25429\
        );

    \I__3447\ : InMux
    port map (
            O => \N__25432\,
            I => \N__25426\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__25429\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__25426\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5\
        );

    \I__3444\ : InMux
    port map (
            O => \N__25421\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4\
        );

    \I__3443\ : InMux
    port map (
            O => \N__25418\,
            I => \N__25414\
        );

    \I__3442\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25411\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__25414\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__25411\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6\
        );

    \I__3439\ : InMux
    port map (
            O => \N__25406\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5\
        );

    \I__3438\ : InMux
    port map (
            O => \N__25403\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6\
        );

    \I__3437\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25396\
        );

    \I__3436\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25393\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__25396\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__25393\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7\
        );

    \I__3433\ : InMux
    port map (
            O => \N__25388\,
            I => \sCounter_cry_16\
        );

    \I__3432\ : InMux
    port map (
            O => \N__25385\,
            I => \sCounter_cry_17\
        );

    \I__3431\ : InMux
    port map (
            O => \N__25382\,
            I => \sCounter_cry_18\
        );

    \I__3430\ : InMux
    port map (
            O => \N__25379\,
            I => \sCounter_cry_19\
        );

    \I__3429\ : InMux
    port map (
            O => \N__25376\,
            I => \sCounter_cry_20\
        );

    \I__3428\ : InMux
    port map (
            O => \N__25373\,
            I => \sCounter_cry_21\
        );

    \I__3427\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25340\
        );

    \I__3426\ : InMux
    port map (
            O => \N__25369\,
            I => \N__25340\
        );

    \I__3425\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25340\
        );

    \I__3424\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25331\
        );

    \I__3423\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25331\
        );

    \I__3422\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25331\
        );

    \I__3421\ : InMux
    port map (
            O => \N__25364\,
            I => \N__25331\
        );

    \I__3420\ : InMux
    port map (
            O => \N__25363\,
            I => \N__25322\
        );

    \I__3419\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25322\
        );

    \I__3418\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25322\
        );

    \I__3417\ : InMux
    port map (
            O => \N__25360\,
            I => \N__25322\
        );

    \I__3416\ : InMux
    port map (
            O => \N__25359\,
            I => \N__25311\
        );

    \I__3415\ : InMux
    port map (
            O => \N__25358\,
            I => \N__25311\
        );

    \I__3414\ : InMux
    port map (
            O => \N__25357\,
            I => \N__25311\
        );

    \I__3413\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25311\
        );

    \I__3412\ : InMux
    port map (
            O => \N__25355\,
            I => \N__25311\
        );

    \I__3411\ : InMux
    port map (
            O => \N__25354\,
            I => \N__25302\
        );

    \I__3410\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25302\
        );

    \I__3409\ : InMux
    port map (
            O => \N__25352\,
            I => \N__25302\
        );

    \I__3408\ : InMux
    port map (
            O => \N__25351\,
            I => \N__25302\
        );

    \I__3407\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25293\
        );

    \I__3406\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25293\
        );

    \I__3405\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25293\
        );

    \I__3404\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25293\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__25340\,
            I => \N__25288\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__25331\,
            I => \N__25288\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__25322\,
            I => \N__25281\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__25311\,
            I => \N__25281\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__25302\,
            I => \N__25281\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__25293\,
            I => \LED_ACQ_c_i\
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__25288\,
            I => \LED_ACQ_c_i\
        );

    \I__3396\ : Odrv4
    port map (
            O => \N__25281\,
            I => \LED_ACQ_c_i\
        );

    \I__3395\ : InMux
    port map (
            O => \N__25274\,
            I => \sCounter_cry_22\
        );

    \I__3394\ : InMux
    port map (
            O => \N__25271\,
            I => \N__25267\
        );

    \I__3393\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25264\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__25267\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__25264\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0\
        );

    \I__3390\ : InMux
    port map (
            O => \N__25259\,
            I => \bfn_11_13_0_\
        );

    \I__3389\ : InMux
    port map (
            O => \N__25256\,
            I => \N__25252\
        );

    \I__3388\ : InMux
    port map (
            O => \N__25255\,
            I => \N__25249\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__25252\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__25249\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1\
        );

    \I__3385\ : InMux
    port map (
            O => \N__25244\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0\
        );

    \I__3384\ : InMux
    port map (
            O => \N__25241\,
            I => \bfn_11_11_0_\
        );

    \I__3383\ : InMux
    port map (
            O => \N__25238\,
            I => \sCounter_cry_8\
        );

    \I__3382\ : InMux
    port map (
            O => \N__25235\,
            I => \sCounter_cry_9\
        );

    \I__3381\ : InMux
    port map (
            O => \N__25232\,
            I => \sCounter_cry_10\
        );

    \I__3380\ : InMux
    port map (
            O => \N__25229\,
            I => \sCounter_cry_11\
        );

    \I__3379\ : InMux
    port map (
            O => \N__25226\,
            I => \sCounter_cry_12\
        );

    \I__3378\ : InMux
    port map (
            O => \N__25223\,
            I => \sCounter_cry_13\
        );

    \I__3377\ : InMux
    port map (
            O => \N__25220\,
            I => \sCounter_cry_14\
        );

    \I__3376\ : InMux
    port map (
            O => \N__25217\,
            I => \bfn_11_12_0_\
        );

    \I__3375\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25210\
        );

    \I__3374\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25207\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__25210\,
            I => \N__25203\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__25207\,
            I => \N__25200\
        );

    \I__3371\ : InMux
    port map (
            O => \N__25206\,
            I => \N__25197\
        );

    \I__3370\ : Span4Mux_v
    port map (
            O => \N__25203\,
            I => \N__25194\
        );

    \I__3369\ : Odrv4
    port map (
            O => \N__25200\,
            I => \sTrigInternalZ0\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__25197\,
            I => \sTrigInternalZ0\
        );

    \I__3367\ : Odrv4
    port map (
            O => \N__25194\,
            I => \sTrigInternalZ0\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__25187\,
            I => \N__25184\
        );

    \I__3365\ : InMux
    port map (
            O => \N__25184\,
            I => \N__25180\
        );

    \I__3364\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25177\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__25180\,
            I => \N__25174\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__25177\,
            I => \N__25171\
        );

    \I__3361\ : Sp12to4
    port map (
            O => \N__25174\,
            I => \N__25168\
        );

    \I__3360\ : Span4Mux_v
    port map (
            O => \N__25171\,
            I => \N__25165\
        );

    \I__3359\ : Odrv12
    port map (
            O => \N__25168\,
            I => op_gt_op_gt_un13_striginternal_0
        );

    \I__3358\ : Odrv4
    port map (
            O => \N__25165\,
            I => op_gt_op_gt_un13_striginternal_0
        );

    \I__3357\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25153\
        );

    \I__3356\ : InMux
    port map (
            O => \N__25159\,
            I => \N__25153\
        );

    \I__3355\ : InMux
    port map (
            O => \N__25158\,
            I => \N__25149\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__25153\,
            I => \N__25146\
        );

    \I__3353\ : InMux
    port map (
            O => \N__25152\,
            I => \N__25143\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__25149\,
            I => \N__25138\
        );

    \I__3351\ : Span4Mux_v
    port map (
            O => \N__25146\,
            I => \N__25138\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__25143\,
            I => \un4_speriod_cry_23_THRU_CO\
        );

    \I__3349\ : Odrv4
    port map (
            O => \N__25138\,
            I => \un4_speriod_cry_23_THRU_CO\
        );

    \I__3348\ : InMux
    port map (
            O => \N__25133\,
            I => \bfn_11_10_0_\
        );

    \I__3347\ : InMux
    port map (
            O => \N__25130\,
            I => \sCounter_cry_0\
        );

    \I__3346\ : InMux
    port map (
            O => \N__25127\,
            I => \sCounter_cry_1\
        );

    \I__3345\ : InMux
    port map (
            O => \N__25124\,
            I => \sCounter_cry_2\
        );

    \I__3344\ : InMux
    port map (
            O => \N__25121\,
            I => \sCounter_cry_3\
        );

    \I__3343\ : InMux
    port map (
            O => \N__25118\,
            I => \sCounter_cry_4\
        );

    \I__3342\ : InMux
    port map (
            O => \N__25115\,
            I => \sCounter_cry_5\
        );

    \I__3341\ : InMux
    port map (
            O => \N__25112\,
            I => \sCounter_cry_6\
        );

    \I__3340\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25106\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__25106\,
            I => \sEEPeriodZ0Z_19\
        );

    \I__3338\ : InMux
    port map (
            O => \N__25103\,
            I => \N__25100\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__25100\,
            I => \sEEPeriod_i_19\
        );

    \I__3336\ : InMux
    port map (
            O => \N__25097\,
            I => \N__25094\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__25094\,
            I => \sEEPeriodZ0Z_20\
        );

    \I__3334\ : InMux
    port map (
            O => \N__25091\,
            I => \N__25088\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__25088\,
            I => \sEEPeriod_i_20\
        );

    \I__3332\ : InMux
    port map (
            O => \N__25085\,
            I => \N__25082\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__25082\,
            I => \sEEPeriodZ0Z_21\
        );

    \I__3330\ : InMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__25076\,
            I => \sEEPeriod_i_21\
        );

    \I__3328\ : InMux
    port map (
            O => \N__25073\,
            I => \N__25070\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__25070\,
            I => \sEEPeriodZ0Z_22\
        );

    \I__3326\ : InMux
    port map (
            O => \N__25067\,
            I => \N__25064\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__25064\,
            I => \sEEPeriod_i_22\
        );

    \I__3324\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25058\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__25058\,
            I => \sEEPeriodZ0Z_23\
        );

    \I__3322\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__25052\,
            I => \sEEPeriod_i_23\
        );

    \I__3320\ : InMux
    port map (
            O => \N__25049\,
            I => \bfn_11_9_0_\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__25046\,
            I => \N__25043\
        );

    \I__3318\ : InMux
    port map (
            O => \N__25043\,
            I => \N__25040\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__25040\,
            I => \N__25037\
        );

    \I__3316\ : Span4Mux_h
    port map (
            O => \N__25037\,
            I => \N__25034\
        );

    \I__3315\ : Odrv4
    port map (
            O => \N__25034\,
            I => un1_spointer11_2_0_0_a2_6
        );

    \I__3314\ : InMux
    port map (
            O => \N__25031\,
            I => \N__25028\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__25028\,
            I => un1_spointer11_2_0_0_a2_1
        );

    \I__3312\ : InMux
    port map (
            O => \N__25025\,
            I => \N__25022\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__25022\,
            I => \sEEPeriodZ0Z_11\
        );

    \I__3310\ : InMux
    port map (
            O => \N__25019\,
            I => \N__25016\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__25016\,
            I => \sEEPeriod_i_11\
        );

    \I__3308\ : InMux
    port map (
            O => \N__25013\,
            I => \N__25010\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__25010\,
            I => \sEEPeriodZ0Z_12\
        );

    \I__3306\ : InMux
    port map (
            O => \N__25007\,
            I => \N__25004\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__25004\,
            I => \sEEPeriod_i_12\
        );

    \I__3304\ : InMux
    port map (
            O => \N__25001\,
            I => \N__24998\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__24998\,
            I => \sEEPeriodZ0Z_13\
        );

    \I__3302\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24992\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__24992\,
            I => \sEEPeriod_i_13\
        );

    \I__3300\ : InMux
    port map (
            O => \N__24989\,
            I => \N__24986\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__24986\,
            I => \sEEPeriodZ0Z_14\
        );

    \I__3298\ : InMux
    port map (
            O => \N__24983\,
            I => \N__24980\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__24980\,
            I => \sEEPeriod_i_14\
        );

    \I__3296\ : InMux
    port map (
            O => \N__24977\,
            I => \N__24974\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__24974\,
            I => \sEEPeriodZ0Z_15\
        );

    \I__3294\ : InMux
    port map (
            O => \N__24971\,
            I => \N__24968\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__24968\,
            I => \sEEPeriod_i_15\
        );

    \I__3292\ : InMux
    port map (
            O => \N__24965\,
            I => \N__24962\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__24962\,
            I => \sEEPeriodZ0Z_16\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24956\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__24956\,
            I => \sEEPeriod_i_16\
        );

    \I__3288\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24950\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__24950\,
            I => \sEEPeriodZ0Z_17\
        );

    \I__3286\ : InMux
    port map (
            O => \N__24947\,
            I => \N__24944\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__24944\,
            I => \sEEPeriod_i_17\
        );

    \I__3284\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24938\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__24938\,
            I => \sEEPeriodZ0Z_18\
        );

    \I__3282\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24932\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__24932\,
            I => \sEEPeriod_i_18\
        );

    \I__3280\ : InMux
    port map (
            O => \N__24929\,
            I => \N__24926\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__24926\,
            I => \sEEPeriod_i_3\
        );

    \I__3278\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24920\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__24920\,
            I => \sEEPeriodZ0Z_4\
        );

    \I__3276\ : InMux
    port map (
            O => \N__24917\,
            I => \N__24914\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__24914\,
            I => \sEEPeriod_i_4\
        );

    \I__3274\ : InMux
    port map (
            O => \N__24911\,
            I => \N__24908\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__24908\,
            I => \sEEPeriodZ0Z_5\
        );

    \I__3272\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24902\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__24902\,
            I => \sEEPeriod_i_5\
        );

    \I__3270\ : InMux
    port map (
            O => \N__24899\,
            I => \N__24896\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__24896\,
            I => \sEEPeriodZ0Z_6\
        );

    \I__3268\ : InMux
    port map (
            O => \N__24893\,
            I => \N__24890\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__24890\,
            I => \sEEPeriod_i_6\
        );

    \I__3266\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24884\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__24884\,
            I => \sEEPeriodZ0Z_7\
        );

    \I__3264\ : CascadeMux
    port map (
            O => \N__24881\,
            I => \N__24878\
        );

    \I__3263\ : InMux
    port map (
            O => \N__24878\,
            I => \N__24875\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__24875\,
            I => \sEEPeriod_i_7\
        );

    \I__3261\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24869\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__24869\,
            I => \sEEPeriodZ0Z_8\
        );

    \I__3259\ : InMux
    port map (
            O => \N__24866\,
            I => \N__24863\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__24863\,
            I => \sEEPeriod_i_8\
        );

    \I__3257\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24857\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__24857\,
            I => \sEEPeriodZ0Z_9\
        );

    \I__3255\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24851\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__24851\,
            I => \sEEPeriod_i_9\
        );

    \I__3253\ : InMux
    port map (
            O => \N__24848\,
            I => \N__24845\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__24845\,
            I => \sEEPeriodZ0Z_10\
        );

    \I__3251\ : InMux
    port map (
            O => \N__24842\,
            I => \N__24839\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__24839\,
            I => \sEEPeriod_i_10\
        );

    \I__3249\ : CEMux
    port map (
            O => \N__24836\,
            I => \N__24833\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__24833\,
            I => \N__24830\
        );

    \I__3247\ : Span4Mux_v
    port map (
            O => \N__24830\,
            I => \N__24827\
        );

    \I__3246\ : Odrv4
    port map (
            O => \N__24827\,
            I => \sAddress_RNIETI62Z0Z_1\
        );

    \I__3245\ : InMux
    port map (
            O => \N__24824\,
            I => \N__24821\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__24821\,
            I => \sEEPeriodZ0Z_0\
        );

    \I__3243\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24815\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__24815\,
            I => \sEEPeriod_i_0\
        );

    \I__3241\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__24809\,
            I => \sEEPeriodZ0Z_1\
        );

    \I__3239\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24803\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__24803\,
            I => \sEEPeriod_i_1\
        );

    \I__3237\ : InMux
    port map (
            O => \N__24800\,
            I => \N__24797\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__24797\,
            I => \sEEPeriodZ0Z_2\
        );

    \I__3235\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24791\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__24791\,
            I => \sEEPeriod_i_2\
        );

    \I__3233\ : InMux
    port map (
            O => \N__24788\,
            I => \N__24785\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__24785\,
            I => \sEEPeriodZ0Z_3\
        );

    \I__3231\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24779\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__24779\,
            I => \sDAC_dataZ0Z_0\
        );

    \I__3229\ : InMux
    port map (
            O => \N__24776\,
            I => \N__24773\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__24773\,
            I => \sDAC_dataZ0Z_1\
        );

    \I__3227\ : InMux
    port map (
            O => \N__24770\,
            I => \N__24767\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__24767\,
            I => \sDAC_dataZ0Z_11\
        );

    \I__3225\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24761\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__24761\,
            I => \sDAC_dataZ0Z_12\
        );

    \I__3223\ : InMux
    port map (
            O => \N__24758\,
            I => \N__24755\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__24755\,
            I => \sDAC_dataZ0Z_13\
        );

    \I__3221\ : InMux
    port map (
            O => \N__24752\,
            I => \N__24749\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__24749\,
            I => \sDAC_dataZ0Z_14\
        );

    \I__3219\ : InMux
    port map (
            O => \N__24746\,
            I => \N__24743\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__24743\,
            I => \sDAC_dataZ0Z_15\
        );

    \I__3217\ : CEMux
    port map (
            O => \N__24740\,
            I => \N__24737\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__24737\,
            I => \N__24734\
        );

    \I__3215\ : Span4Mux_v
    port map (
            O => \N__24734\,
            I => \N__24731\
        );

    \I__3214\ : Span4Mux_v
    port map (
            O => \N__24731\,
            I => \N__24728\
        );

    \I__3213\ : Odrv4
    port map (
            O => \N__24728\,
            I => \sAddress_RNIA6242Z0Z_0\
        );

    \I__3212\ : IoInMux
    port map (
            O => \N__24725\,
            I => \N__24722\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__24722\,
            I => \N__24719\
        );

    \I__3210\ : Span4Mux_s3_v
    port map (
            O => \N__24719\,
            I => \N__24716\
        );

    \I__3209\ : Span4Mux_v
    port map (
            O => \N__24716\,
            I => \N__24713\
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__24713\,
            I => \LED3_c_i\
        );

    \I__3207\ : InMux
    port map (
            O => \N__24710\,
            I => \N__24707\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__24707\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15\
        );

    \I__3205\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24701\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__24701\,
            I => \N__24697\
        );

    \I__3203\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24694\
        );

    \I__3202\ : Span4Mux_h
    port map (
            O => \N__24697\,
            I => \N__24686\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__24694\,
            I => \N__24686\
        );

    \I__3200\ : InMux
    port map (
            O => \N__24693\,
            I => \N__24683\
        );

    \I__3199\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24677\
        );

    \I__3198\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24677\
        );

    \I__3197\ : Span4Mux_h
    port map (
            O => \N__24686\,
            I => \N__24672\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__24683\,
            I => \N__24672\
        );

    \I__3195\ : InMux
    port map (
            O => \N__24682\,
            I => \N__24669\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__24677\,
            I => \N__24664\
        );

    \I__3193\ : Span4Mux_h
    port map (
            O => \N__24672\,
            I => \N__24659\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__24669\,
            I => \N__24659\
        );

    \I__3191\ : InMux
    port map (
            O => \N__24668\,
            I => \N__24656\
        );

    \I__3190\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24653\
        );

    \I__3189\ : Span4Mux_h
    port map (
            O => \N__24664\,
            I => \N__24646\
        );

    \I__3188\ : Span4Mux_v
    port map (
            O => \N__24659\,
            I => \N__24643\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__24656\,
            I => \N__24638\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__24653\,
            I => \N__24638\
        );

    \I__3185\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24633\
        );

    \I__3184\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24633\
        );

    \I__3183\ : InMux
    port map (
            O => \N__24650\,
            I => \N__24630\
        );

    \I__3182\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24627\
        );

    \I__3181\ : Odrv4
    port map (
            O => \N__24646\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__3180\ : Odrv4
    port map (
            O => \N__24643\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__3179\ : Odrv12
    port map (
            O => \N__24638\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__24633\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__24630\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__24627\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__3175\ : InMux
    port map (
            O => \N__24614\,
            I => \N__24611\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__3173\ : Odrv12
    port map (
            O => \N__24608\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15\
        );

    \I__3172\ : CEMux
    port map (
            O => \N__24605\,
            I => \N__24602\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__24602\,
            I => \N__24599\
        );

    \I__3170\ : Span4Mux_v
    port map (
            O => \N__24599\,
            I => \N__24596\
        );

    \I__3169\ : Odrv4
    port map (
            O => \N__24596\,
            I => \sAddress_RNIA6242_4Z0Z_0\
        );

    \I__3168\ : CEMux
    port map (
            O => \N__24593\,
            I => \N__24590\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__24590\,
            I => \N__24587\
        );

    \I__3166\ : Span4Mux_v
    port map (
            O => \N__24587\,
            I => \N__24584\
        );

    \I__3165\ : Span4Mux_h
    port map (
            O => \N__24584\,
            I => \N__24581\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__24581\,
            I => \sDAC_mem_31_1_sqmuxa\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__24578\,
            I => \spi_slave_inst.un23_i_ssn_cascade_\
        );

    \I__3162\ : InMux
    port map (
            O => \N__24575\,
            I => \N__24572\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__24572\,
            I => \N__24569\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__24569\,
            I => g0_10
        );

    \I__3159\ : InMux
    port map (
            O => \N__24566\,
            I => \N__24563\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__24563\,
            I => g0_10_0
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__24560\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2_cascade_\
        );

    \I__3156\ : InMux
    port map (
            O => \N__24557\,
            I => \N__24554\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__24554\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2\
        );

    \I__3154\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24547\
        );

    \I__3153\ : InMux
    port map (
            O => \N__24550\,
            I => \N__24544\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__24547\,
            I => \N__24538\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__24544\,
            I => \N__24538\
        );

    \I__3150\ : InMux
    port map (
            O => \N__24543\,
            I => \N__24535\
        );

    \I__3149\ : Span4Mux_v
    port map (
            O => \N__24538\,
            I => \N__24530\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__24535\,
            I => \N__24530\
        );

    \I__3147\ : Span4Mux_h
    port map (
            O => \N__24530\,
            I => \N__24527\
        );

    \I__3146\ : Span4Mux_h
    port map (
            O => \N__24527\,
            I => \N__24524\
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__24524\,
            I => \spi_master_inst.sclk_gen_u0.N_158_7\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__24521\,
            I => \N__24517\
        );

    \I__3143\ : InMux
    port map (
            O => \N__24520\,
            I => \N__24514\
        );

    \I__3142\ : InMux
    port map (
            O => \N__24517\,
            I => \N__24509\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__24514\,
            I => \N__24506\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__24513\,
            I => \N__24503\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__24512\,
            I => \N__24500\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__24509\,
            I => \N__24496\
        );

    \I__3137\ : Span4Mux_v
    port map (
            O => \N__24506\,
            I => \N__24492\
        );

    \I__3136\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24489\
        );

    \I__3135\ : InMux
    port map (
            O => \N__24500\,
            I => \N__24486\
        );

    \I__3134\ : InMux
    port map (
            O => \N__24499\,
            I => \N__24483\
        );

    \I__3133\ : Span4Mux_h
    port map (
            O => \N__24496\,
            I => \N__24480\
        );

    \I__3132\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24477\
        );

    \I__3131\ : Span4Mux_h
    port map (
            O => \N__24492\,
            I => \N__24474\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__24489\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__24486\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__24483\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__24480\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__24477\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__24474\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\
        );

    \I__3124\ : InMux
    port map (
            O => \N__24461\,
            I => \N__24456\
        );

    \I__3123\ : InMux
    port map (
            O => \N__24460\,
            I => \N__24451\
        );

    \I__3122\ : InMux
    port map (
            O => \N__24459\,
            I => \N__24448\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__24456\,
            I => \N__24445\
        );

    \I__3120\ : InMux
    port map (
            O => \N__24455\,
            I => \N__24442\
        );

    \I__3119\ : InMux
    port map (
            O => \N__24454\,
            I => \N__24439\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__24451\,
            I => \N__24434\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__24448\,
            I => \N__24434\
        );

    \I__3116\ : Span4Mux_h
    port map (
            O => \N__24445\,
            I => \N__24431\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__24442\,
            I => \N__24428\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__24439\,
            I => \N__24425\
        );

    \I__3113\ : Span4Mux_h
    port map (
            O => \N__24434\,
            I => \N__24422\
        );

    \I__3112\ : Span4Mux_h
    port map (
            O => \N__24431\,
            I => \N__24419\
        );

    \I__3111\ : Span4Mux_v
    port map (
            O => \N__24428\,
            I => \N__24416\
        );

    \I__3110\ : Span4Mux_v
    port map (
            O => \N__24425\,
            I => \N__24413\
        );

    \I__3109\ : Span4Mux_h
    port map (
            O => \N__24422\,
            I => \N__24410\
        );

    \I__3108\ : Span4Mux_v
    port map (
            O => \N__24419\,
            I => \N__24407\
        );

    \I__3107\ : Span4Mux_v
    port map (
            O => \N__24416\,
            I => \N__24404\
        );

    \I__3106\ : Span4Mux_h
    port map (
            O => \N__24413\,
            I => \N__24399\
        );

    \I__3105\ : Span4Mux_v
    port map (
            O => \N__24410\,
            I => \N__24399\
        );

    \I__3104\ : Odrv4
    port map (
            O => \N__24407\,
            I => \spi_master_inst.sclk_gen_u0.spi_start_iZ0\
        );

    \I__3103\ : Odrv4
    port map (
            O => \N__24404\,
            I => \spi_master_inst.sclk_gen_u0.spi_start_iZ0\
        );

    \I__3102\ : Odrv4
    port map (
            O => \N__24399\,
            I => \spi_master_inst.sclk_gen_u0.spi_start_iZ0\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__24392\,
            I => \spi_master_inst.sclk_gen_u0.N_158_7_cascade_\
        );

    \I__3100\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24382\
        );

    \I__3099\ : InMux
    port map (
            O => \N__24388\,
            I => \N__24379\
        );

    \I__3098\ : CascadeMux
    port map (
            O => \N__24387\,
            I => \N__24375\
        );

    \I__3097\ : InMux
    port map (
            O => \N__24386\,
            I => \N__24372\
        );

    \I__3096\ : InMux
    port map (
            O => \N__24385\,
            I => \N__24369\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__24382\,
            I => \N__24366\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__24379\,
            I => \N__24363\
        );

    \I__3093\ : InMux
    port map (
            O => \N__24378\,
            I => \N__24360\
        );

    \I__3092\ : InMux
    port map (
            O => \N__24375\,
            I => \N__24357\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__24372\,
            I => \N__24354\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__24369\,
            I => \N__24349\
        );

    \I__3089\ : Span4Mux_v
    port map (
            O => \N__24366\,
            I => \N__24349\
        );

    \I__3088\ : Span12Mux_h
    port map (
            O => \N__24363\,
            I => \N__24346\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__24360\,
            I => \N__24339\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__24357\,
            I => \N__24339\
        );

    \I__3085\ : Span4Mux_h
    port map (
            O => \N__24354\,
            I => \N__24339\
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__24349\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\
        );

    \I__3083\ : Odrv12
    port map (
            O => \N__24346\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__24339\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\
        );

    \I__3081\ : InMux
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__24329\,
            I => \N__24326\
        );

    \I__3079\ : Span4Mux_h
    port map (
            O => \N__24326\,
            I => \N__24323\
        );

    \I__3078\ : Span4Mux_v
    port map (
            O => \N__24323\,
            I => \N__24320\
        );

    \I__3077\ : Span4Mux_h
    port map (
            O => \N__24320\,
            I => \N__24317\
        );

    \I__3076\ : Odrv4
    port map (
            O => \N__24317\,
            I => \spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0\
        );

    \I__3075\ : InMux
    port map (
            O => \N__24314\,
            I => \N__24311\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__24311\,
            I => g2_6
        );

    \I__3073\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24305\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__24305\,
            I => \N__24301\
        );

    \I__3071\ : InMux
    port map (
            O => \N__24304\,
            I => \N__24298\
        );

    \I__3070\ : Span4Mux_h
    port map (
            O => \N__24301\,
            I => \N__24295\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__24298\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__24295\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__3067\ : InMux
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__24287\,
            I => \N__24283\
        );

    \I__3065\ : InMux
    port map (
            O => \N__24286\,
            I => \N__24280\
        );

    \I__3064\ : Span4Mux_h
    port map (
            O => \N__24283\,
            I => \N__24277\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__24280\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__3062\ : Odrv4
    port map (
            O => \N__24277\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__3061\ : InMux
    port map (
            O => \N__24272\,
            I => \N__24269\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__24269\,
            I => \N__24266\
        );

    \I__3059\ : Span4Mux_v
    port map (
            O => \N__24266\,
            I => \N__24263\
        );

    \I__3058\ : Span4Mux_h
    port map (
            O => \N__24263\,
            I => \N__24260\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__24260\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_i6_3\
        );

    \I__3056\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24251\
        );

    \I__3055\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24248\
        );

    \I__3054\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24243\
        );

    \I__3053\ : InMux
    port map (
            O => \N__24254\,
            I => \N__24243\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__24251\,
            I => \N__24240\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__24248\,
            I => \N__24235\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__24243\,
            I => \N__24235\
        );

    \I__3049\ : Span4Mux_h
    port map (
            O => \N__24240\,
            I => \N__24232\
        );

    \I__3048\ : Span12Mux_h
    port map (
            O => \N__24235\,
            I => \N__24227\
        );

    \I__3047\ : Sp12to4
    port map (
            O => \N__24232\,
            I => \N__24227\
        );

    \I__3046\ : Odrv12
    port map (
            O => \N__24227\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_i6\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__24224\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__24221\,
            I => \N__24217\
        );

    \I__3043\ : InMux
    port map (
            O => \N__24220\,
            I => \N__24214\
        );

    \I__3042\ : InMux
    port map (
            O => \N__24217\,
            I => \N__24211\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__24214\,
            I => \N__24206\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__24211\,
            I => \N__24206\
        );

    \I__3039\ : Span4Mux_h
    port map (
            O => \N__24206\,
            I => \N__24203\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__24203\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_3\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__24200\,
            I => \spi_slave_inst.un23_i_ssn_3_cascade_\
        );

    \I__3036\ : InMux
    port map (
            O => \N__24197\,
            I => \N__24194\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__24194\,
            I => \N__24191\
        );

    \I__3034\ : Span4Mux_v
    port map (
            O => \N__24191\,
            I => \N__24188\
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__24188\,
            I => un21_trig_prev_21_5
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__24185\,
            I => \op_gt_op_gt_un13_striginternallto23_5_cascade_\
        );

    \I__3031\ : InMux
    port map (
            O => \N__24182\,
            I => \N__24179\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__24179\,
            I => \N__24176\
        );

    \I__3029\ : Odrv12
    port map (
            O => \N__24176\,
            I => un1_reset_rpi_inv_2_0_o2_2
        );

    \I__3028\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24170\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__24170\,
            I => g0_13_0
        );

    \I__3026\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24164\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__24164\,
            I => un21_trig_prev_21_4
        );

    \I__3024\ : InMux
    port map (
            O => \N__24161\,
            I => \N__24158\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__24158\,
            I => g0_6
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__24155\,
            I => \N__24152\
        );

    \I__3021\ : InMux
    port map (
            O => \N__24152\,
            I => \N__24149\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__24149\,
            I => \N__24146\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__24146\,
            I => \N_99\
        );

    \I__3018\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24140\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__24140\,
            I => op_gt_op_gt_un13_striginternallto23_3
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__24137\,
            I => \N__24133\
        );

    \I__3015\ : InMux
    port map (
            O => \N__24136\,
            I => \N__24130\
        );

    \I__3014\ : InMux
    port map (
            O => \N__24133\,
            I => \N__24127\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__24130\,
            I => \N__24124\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__24127\,
            I => \N_831_16\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__24124\,
            I => \N_831_16\
        );

    \I__3010\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24116\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__24116\,
            I => op_gt_op_gt_un13_striginternallto23_6
        );

    \I__3008\ : CEMux
    port map (
            O => \N__24113\,
            I => \N__24110\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__24110\,
            I => \sDAC_mem_15_1_sqmuxa\
        );

    \I__3006\ : CEMux
    port map (
            O => \N__24107\,
            I => \N__24104\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__24104\,
            I => \N__24101\
        );

    \I__3004\ : Span4Mux_v
    port map (
            O => \N__24101\,
            I => \N__24098\
        );

    \I__3003\ : Span4Mux_h
    port map (
            O => \N__24098\,
            I => \N__24095\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__24095\,
            I => \sAddress_RNI9IH12_1Z0Z_2\
        );

    \I__3001\ : CEMux
    port map (
            O => \N__24092\,
            I => \N__24089\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__24089\,
            I => \N__24086\
        );

    \I__2999\ : Span4Mux_v
    port map (
            O => \N__24086\,
            I => \N__24083\
        );

    \I__2998\ : Span4Mux_h
    port map (
            O => \N__24083\,
            I => \N__24080\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__24080\,
            I => \sDAC_mem_14_1_sqmuxa\
        );

    \I__2996\ : CEMux
    port map (
            O => \N__24077\,
            I => \N__24074\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__24074\,
            I => \N__24071\
        );

    \I__2994\ : Span4Mux_h
    port map (
            O => \N__24071\,
            I => \N__24068\
        );

    \I__2993\ : Span4Mux_h
    port map (
            O => \N__24068\,
            I => \N__24065\
        );

    \I__2992\ : Odrv4
    port map (
            O => \N__24065\,
            I => \sAddress_RNI9IH12Z0Z_0\
        );

    \I__2991\ : CEMux
    port map (
            O => \N__24062\,
            I => \N__24059\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__24059\,
            I => \N__24056\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__24056\,
            I => \sDAC_mem_42_1_sqmuxa\
        );

    \I__2988\ : InMux
    port map (
            O => \N__24053\,
            I => \N__24050\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__24050\,
            I => \N__24047\
        );

    \I__2986\ : Span4Mux_h
    port map (
            O => \N__24047\,
            I => \N__24044\
        );

    \I__2985\ : Odrv4
    port map (
            O => \N__24044\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_11\
        );

    \I__2984\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24038\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__24038\,
            I => \N__24035\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__24035\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_13\
        );

    \I__2981\ : InMux
    port map (
            O => \N__24032\,
            I => \N__24029\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__24029\,
            I => \N__24026\
        );

    \I__2979\ : Odrv4
    port map (
            O => \N__24026\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_14\
        );

    \I__2978\ : InMux
    port map (
            O => \N__24023\,
            I => \N__24020\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__24020\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_15\
        );

    \I__2976\ : InMux
    port map (
            O => \N__24017\,
            I => \bfn_9_20_0_\
        );

    \I__2975\ : IoInMux
    port map (
            O => \N__24014\,
            I => \N__24011\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__24008\
        );

    \I__2973\ : Span12Mux_s0_h
    port map (
            O => \N__24008\,
            I => \N__24005\
        );

    \I__2972\ : Span12Mux_h
    port map (
            O => \N__24005\,
            I => \N__24002\
        );

    \I__2971\ : Odrv12
    port map (
            O => \N__24002\,
            I => \pon_obuf_RNOZ0\
        );

    \I__2970\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23996\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__23996\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10\
        );

    \I__2968\ : InMux
    port map (
            O => \N__23993\,
            I => \N__23990\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__23990\,
            I => \N__23987\
        );

    \I__2966\ : Odrv12
    port map (
            O => \N__23987\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_0\
        );

    \I__2965\ : InMux
    port map (
            O => \N__23984\,
            I => \N__23981\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__23981\,
            I => \N__23978\
        );

    \I__2963\ : Odrv12
    port map (
            O => \N__23978\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_1\
        );

    \I__2962\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23972\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__23972\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_10\
        );

    \I__2960\ : InMux
    port map (
            O => \N__23969\,
            I => \N__23966\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__23966\,
            I => \sEEPonZ0Z_4\
        );

    \I__2958\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23960\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__23960\,
            I => \sEEPon_i_4\
        );

    \I__2956\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23954\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__23954\,
            I => \sEEPonZ0Z_5\
        );

    \I__2954\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23948\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__23948\,
            I => \sEEPon_i_5\
        );

    \I__2952\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23942\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__23942\,
            I => \sEEPonZ0Z_6\
        );

    \I__2950\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23936\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__23936\,
            I => \sEEPon_i_6\
        );

    \I__2948\ : InMux
    port map (
            O => \N__23933\,
            I => \N__23930\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__23930\,
            I => \sEEPonZ0Z_7\
        );

    \I__2946\ : InMux
    port map (
            O => \N__23927\,
            I => \N__23924\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__23924\,
            I => \sEEPon_i_7\
        );

    \I__2944\ : CEMux
    port map (
            O => \N__23921\,
            I => \N__23918\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__23918\,
            I => \N__23915\
        );

    \I__2942\ : Sp12to4
    port map (
            O => \N__23915\,
            I => \N__23912\
        );

    \I__2941\ : Odrv12
    port map (
            O => \N__23912\,
            I => \sDAC_mem_30_1_sqmuxa\
        );

    \I__2940\ : InMux
    port map (
            O => \N__23909\,
            I => \N__23906\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__23906\,
            I => \sEEPonZ0Z_0\
        );

    \I__2938\ : CascadeMux
    port map (
            O => \N__23903\,
            I => \N__23900\
        );

    \I__2937\ : InMux
    port map (
            O => \N__23900\,
            I => \N__23897\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__23897\,
            I => \sEEPon_i_0\
        );

    \I__2935\ : InMux
    port map (
            O => \N__23894\,
            I => \N__23891\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__23891\,
            I => \sEEPonZ0Z_1\
        );

    \I__2933\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__23885\,
            I => \sEEPon_i_1\
        );

    \I__2931\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__23879\,
            I => \sEEPonZ0Z_2\
        );

    \I__2929\ : InMux
    port map (
            O => \N__23876\,
            I => \N__23873\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__23873\,
            I => \sEEPon_i_2\
        );

    \I__2927\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23867\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__23867\,
            I => \sEEPonZ0Z_3\
        );

    \I__2925\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23861\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__23861\,
            I => \sEEPon_i_3\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__23858\,
            I => \N__23855\
        );

    \I__2922\ : InMux
    port map (
            O => \N__23855\,
            I => \N__23852\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__23852\,
            I => g0_13_1
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__23849\,
            I => \N__23846\
        );

    \I__2919\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23843\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__23843\,
            I => g0_17_0
        );

    \I__2917\ : InMux
    port map (
            O => \N__23840\,
            I => \N__23837\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__23837\,
            I => \N__23831\
        );

    \I__2915\ : InMux
    port map (
            O => \N__23836\,
            I => \N__23828\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__23835\,
            I => \N__23825\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__23834\,
            I => \N__23820\
        );

    \I__2912\ : Span4Mux_v
    port map (
            O => \N__23831\,
            I => \N__23817\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__23828\,
            I => \N__23814\
        );

    \I__2910\ : InMux
    port map (
            O => \N__23825\,
            I => \N__23805\
        );

    \I__2909\ : InMux
    port map (
            O => \N__23824\,
            I => \N__23805\
        );

    \I__2908\ : InMux
    port map (
            O => \N__23823\,
            I => \N__23805\
        );

    \I__2907\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23805\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__23817\,
            I => \N_326\
        );

    \I__2905\ : Odrv12
    port map (
            O => \N__23814\,
            I => \N_326\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__23805\,
            I => \N_326\
        );

    \I__2903\ : InMux
    port map (
            O => \N__23798\,
            I => \N__23795\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__23795\,
            I => g0_16_0
        );

    \I__2901\ : InMux
    port map (
            O => \N__23792\,
            I => \N__23789\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__23789\,
            I => g1_i_a4_6
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__23786\,
            I => \g1_i_a4_5_cascade_\
        );

    \I__2898\ : InMux
    port map (
            O => \N__23783\,
            I => \N__23780\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__23780\,
            I => \N__23777\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__23777\,
            I => un1_reset_rpi_inv_2_0_o2_5
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__23774\,
            I => \g1_i_a4_9_cascade_\
        );

    \I__2894\ : InMux
    port map (
            O => \N__23771\,
            I => \N__23768\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__23768\,
            I => \N__23765\
        );

    \I__2892\ : Odrv4
    port map (
            O => \N__23765\,
            I => \sEETrigInternal_prev_RNIH3OJZ0Z1\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__23762\,
            I => \N__23759\
        );

    \I__2890\ : InMux
    port map (
            O => \N__23759\,
            I => \N__23756\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__23756\,
            I => \N__23753\
        );

    \I__2888\ : Span4Mux_h
    port map (
            O => \N__23753\,
            I => \N__23750\
        );

    \I__2887\ : Odrv4
    port map (
            O => \N__23750\,
            I => g0_0_1
        );

    \I__2886\ : InMux
    port map (
            O => \N__23747\,
            I => \N__23744\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__23744\,
            I => g0_16
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__23741\,
            I => \N__23738\
        );

    \I__2883\ : InMux
    port map (
            O => \N__23738\,
            I => \N__23735\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__23735\,
            I => \N__23732\
        );

    \I__2881\ : Span4Mux_v
    port map (
            O => \N__23732\,
            I => \N__23729\
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__23729\,
            I => g0_11
        );

    \I__2879\ : InMux
    port map (
            O => \N__23726\,
            I => \N__23723\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__23723\,
            I => g0_14
        );

    \I__2877\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23715\
        );

    \I__2876\ : InMux
    port map (
            O => \N__23719\,
            I => \N__23712\
        );

    \I__2875\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23708\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__23715\,
            I => \N__23699\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__23712\,
            I => \N__23699\
        );

    \I__2872\ : InMux
    port map (
            O => \N__23711\,
            I => \N__23696\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__23708\,
            I => \N__23693\
        );

    \I__2870\ : InMux
    port map (
            O => \N__23707\,
            I => \N__23688\
        );

    \I__2869\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23688\
        );

    \I__2868\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23683\
        );

    \I__2867\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23683\
        );

    \I__2866\ : Sp12to4
    port map (
            O => \N__23699\,
            I => \N__23678\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__23696\,
            I => \N__23678\
        );

    \I__2864\ : Span4Mux_v
    port map (
            O => \N__23693\,
            I => \N__23675\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__23688\,
            I => \sEETrigInternalZ0\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__23683\,
            I => \sEETrigInternalZ0\
        );

    \I__2861\ : Odrv12
    port map (
            O => \N__23678\,
            I => \sEETrigInternalZ0\
        );

    \I__2860\ : Odrv4
    port map (
            O => \N__23675\,
            I => \sEETrigInternalZ0\
        );

    \I__2859\ : InMux
    port map (
            O => \N__23666\,
            I => \N__23663\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__23663\,
            I => \N__23660\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__23660\,
            I => g3_0
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__23657\,
            I => \N__23652\
        );

    \I__2855\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23649\
        );

    \I__2854\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23646\
        );

    \I__2853\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23642\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__23649\,
            I => \N__23637\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__23646\,
            I => \N__23637\
        );

    \I__2850\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23634\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__23642\,
            I => \N__23631\
        );

    \I__2848\ : Sp12to4
    port map (
            O => \N__23637\,
            I => \N__23628\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__23634\,
            I => \N__23623\
        );

    \I__2846\ : Span4Mux_h
    port map (
            O => \N__23631\,
            I => \N__23623\
        );

    \I__2845\ : Odrv12
    port map (
            O => \N__23628\,
            I => \sEETrigInternal_prevZ0\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__23623\,
            I => \sEETrigInternal_prevZ0\
        );

    \I__2843\ : IoInMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__2841\ : Span4Mux_s1_h
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__2840\ : Span4Mux_h
    port map (
            O => \N__23609\,
            I => \N__23603\
        );

    \I__2839\ : InMux
    port map (
            O => \N__23608\,
            I => \N__23598\
        );

    \I__2838\ : InMux
    port map (
            O => \N__23607\,
            I => \N__23598\
        );

    \I__2837\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23595\
        );

    \I__2836\ : Sp12to4
    port map (
            O => \N__23603\,
            I => \N__23592\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__23598\,
            I => \N__23589\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__23595\,
            I => \N__23586\
        );

    \I__2833\ : Span12Mux_v
    port map (
            O => \N__23592\,
            I => \N__23583\
        );

    \I__2832\ : Span4Mux_h
    port map (
            O => \N__23589\,
            I => \N__23580\
        );

    \I__2831\ : Span4Mux_h
    port map (
            O => \N__23586\,
            I => \N__23577\
        );

    \I__2830\ : Odrv12
    port map (
            O => \N__23583\,
            I => \LED_MODE_c\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__23580\,
            I => \LED_MODE_c\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__23577\,
            I => \LED_MODE_c\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__23570\,
            I => \N_831_16_cascade_\
        );

    \I__2826\ : InMux
    port map (
            O => \N__23567\,
            I => \N__23562\
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__23566\,
            I => \N__23558\
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__23565\,
            I => \N__23555\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__23562\,
            I => \N__23551\
        );

    \I__2822\ : InMux
    port map (
            O => \N__23561\,
            I => \N__23547\
        );

    \I__2821\ : InMux
    port map (
            O => \N__23558\,
            I => \N__23542\
        );

    \I__2820\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23542\
        );

    \I__2819\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23539\
        );

    \I__2818\ : Span4Mux_h
    port map (
            O => \N__23551\,
            I => \N__23536\
        );

    \I__2817\ : InMux
    port map (
            O => \N__23550\,
            I => \N__23533\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__23547\,
            I => \N__23528\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__23542\,
            I => \N__23528\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__23539\,
            I => \N_319\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__23536\,
            I => \N_319\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__23533\,
            I => \N_319\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__23528\,
            I => \N_319\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__23519\,
            I => \g0_13_cascade_\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__23516\,
            I => \N__23513\
        );

    \I__2808\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23510\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__23510\,
            I => g0_1_0
        );

    \I__2806\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23504\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__23504\,
            I => g0_15_0
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__23501\,
            I => \sAddress_RNIAM2A_0Z0Z_1_cascade_\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__23498\,
            I => \N_445_cascade_\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__23495\,
            I => \N__23491\
        );

    \I__2801\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23485\
        );

    \I__2800\ : InMux
    port map (
            O => \N__23491\,
            I => \N__23485\
        );

    \I__2799\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23482\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__23485\,
            I => \N__23479\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__23482\,
            I => \sAddress_RNI6VH7_5Z0Z_1\
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__23479\,
            I => \sAddress_RNI6VH7_5Z0Z_1\
        );

    \I__2795\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23471\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__23471\,
            I => \N_445\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__23468\,
            I => \N__23465\
        );

    \I__2792\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23458\
        );

    \I__2791\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23455\
        );

    \I__2790\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23452\
        );

    \I__2789\ : InMux
    port map (
            O => \N__23462\,
            I => \N__23449\
        );

    \I__2788\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23446\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__23458\,
            I => \N__23434\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__23455\,
            I => \N__23434\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__23452\,
            I => \N__23434\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__23449\,
            I => \N__23434\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__23446\,
            I => \N__23434\
        );

    \I__2782\ : InMux
    port map (
            O => \N__23445\,
            I => \N__23431\
        );

    \I__2781\ : Span4Mux_v
    port map (
            O => \N__23434\,
            I => \N__23428\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__23431\,
            I => \N_316\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__23428\,
            I => \N_316\
        );

    \I__2778\ : CEMux
    port map (
            O => \N__23423\,
            I => \N__23419\
        );

    \I__2777\ : CEMux
    port map (
            O => \N__23422\,
            I => \N__23414\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__23419\,
            I => \N__23410\
        );

    \I__2775\ : CEMux
    port map (
            O => \N__23418\,
            I => \N__23406\
        );

    \I__2774\ : CEMux
    port map (
            O => \N__23417\,
            I => \N__23403\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__23414\,
            I => \N__23400\
        );

    \I__2772\ : CEMux
    port map (
            O => \N__23413\,
            I => \N__23397\
        );

    \I__2771\ : Span4Mux_v
    port map (
            O => \N__23410\,
            I => \N__23394\
        );

    \I__2770\ : CEMux
    port map (
            O => \N__23409\,
            I => \N__23391\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__23406\,
            I => \N__23388\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__23403\,
            I => \N__23385\
        );

    \I__2767\ : Span4Mux_h
    port map (
            O => \N__23400\,
            I => \N__23382\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__23397\,
            I => \N__23379\
        );

    \I__2765\ : Span4Mux_h
    port map (
            O => \N__23394\,
            I => \N__23374\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__23391\,
            I => \N__23374\
        );

    \I__2763\ : Span4Mux_v
    port map (
            O => \N__23388\,
            I => \N__23371\
        );

    \I__2762\ : Span4Mux_h
    port map (
            O => \N__23385\,
            I => \N__23368\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__23382\,
            I => \N__23365\
        );

    \I__2760\ : Span4Mux_v
    port map (
            O => \N__23379\,
            I => \N__23362\
        );

    \I__2759\ : Span4Mux_h
    port map (
            O => \N__23374\,
            I => \N__23359\
        );

    \I__2758\ : Span4Mux_h
    port map (
            O => \N__23371\,
            I => \N__23354\
        );

    \I__2757\ : Span4Mux_h
    port map (
            O => \N__23368\,
            I => \N__23354\
        );

    \I__2756\ : Odrv4
    port map (
            O => \N__23365\,
            I => un1_spointer11_0
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__23362\,
            I => un1_spointer11_0
        );

    \I__2754\ : Odrv4
    port map (
            O => \N__23359\,
            I => un1_spointer11_0
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__23354\,
            I => un1_spointer11_0
        );

    \I__2752\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23341\
        );

    \I__2751\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23337\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__23341\,
            I => \N__23334\
        );

    \I__2749\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23331\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__23337\,
            I => \N__23328\
        );

    \I__2747\ : Span4Mux_h
    port map (
            O => \N__23334\,
            I => \N__23325\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__23331\,
            I => \sAddress_RNI6VH7_2Z0Z_1\
        );

    \I__2745\ : Odrv4
    port map (
            O => \N__23328\,
            I => \sAddress_RNI6VH7_2Z0Z_1\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__23325\,
            I => \sAddress_RNI6VH7_2Z0Z_1\
        );

    \I__2743\ : IoInMux
    port map (
            O => \N__23318\,
            I => \N__23315\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__2741\ : Span12Mux_s0_h
    port map (
            O => \N__23312\,
            I => \N__23309\
        );

    \I__2740\ : Span12Mux_v
    port map (
            O => \N__23309\,
            I => \N__23306\
        );

    \I__2739\ : Span12Mux_h
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__2738\ : Odrv12
    port map (
            O => \N__23303\,
            I => \LED_ACQ_obuf_RNOZ0\
        );

    \I__2737\ : InMux
    port map (
            O => \N__23300\,
            I => \N__23295\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__23299\,
            I => \N__23290\
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__23298\,
            I => \N__23287\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__23295\,
            I => \N__23284\
        );

    \I__2733\ : InMux
    port map (
            O => \N__23294\,
            I => \N__23281\
        );

    \I__2732\ : InMux
    port map (
            O => \N__23293\,
            I => \N__23274\
        );

    \I__2731\ : InMux
    port map (
            O => \N__23290\,
            I => \N__23274\
        );

    \I__2730\ : InMux
    port map (
            O => \N__23287\,
            I => \N__23274\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__23284\,
            I => \sAddress_RNI6VH7_3Z0Z_1\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__23281\,
            I => \sAddress_RNI6VH7_3Z0Z_1\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__23274\,
            I => \sAddress_RNI6VH7_3Z0Z_1\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__23267\,
            I => \sAddress_RNI6VH7_3Z0Z_1_cascade_\
        );

    \I__2725\ : CEMux
    port map (
            O => \N__23264\,
            I => \N__23261\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__23261\,
            I => \N__23258\
        );

    \I__2723\ : Span4Mux_h
    port map (
            O => \N__23258\,
            I => \N__23255\
        );

    \I__2722\ : Span4Mux_h
    port map (
            O => \N__23255\,
            I => \N__23252\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__23252\,
            I => \sDAC_mem_10_1_sqmuxa\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__23249\,
            I => \N_326_cascade_\
        );

    \I__2719\ : CEMux
    port map (
            O => \N__23246\,
            I => \N__23243\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__23243\,
            I => \N__23240\
        );

    \I__2717\ : Span4Mux_v
    port map (
            O => \N__23240\,
            I => \N__23237\
        );

    \I__2716\ : Odrv4
    port map (
            O => \N__23237\,
            I => \sDAC_mem_38_1_sqmuxa\
        );

    \I__2715\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23231\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__23231\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4\
        );

    \I__2713\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23225\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__23225\,
            I => \N__23222\
        );

    \I__2711\ : Odrv12
    port map (
            O => \N__23222\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12\
        );

    \I__2710\ : InMux
    port map (
            O => \N__23219\,
            I => \N__23216\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__23216\,
            I => \N__23213\
        );

    \I__2708\ : Span4Mux_h
    port map (
            O => \N__23213\,
            I => \N__23210\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__23210\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10\
        );

    \I__2706\ : CEMux
    port map (
            O => \N__23207\,
            I => \N__23204\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__23204\,
            I => \N__23201\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__23201\,
            I => \N__23198\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__23198\,
            I => \sEEPon_1_sqmuxa\
        );

    \I__2702\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23192\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__23192\,
            I => \spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0\
        );

    \I__2700\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23183\
        );

    \I__2699\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23183\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__23183\,
            I => \spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0\
        );

    \I__2697\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23177\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__23177\,
            I => \N__23174\
        );

    \I__2695\ : Span4Mux_h
    port map (
            O => \N__23174\,
            I => \N__23171\
        );

    \I__2694\ : Span4Mux_v
    port map (
            O => \N__23171\,
            I => \N__23167\
        );

    \I__2693\ : InMux
    port map (
            O => \N__23170\,
            I => \N__23164\
        );

    \I__2692\ : Odrv4
    port map (
            O => \N__23167\,
            I => \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__23164\,
            I => \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0\
        );

    \I__2690\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23156\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__23156\,
            I => \spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0\
        );

    \I__2688\ : CEMux
    port map (
            O => \N__23153\,
            I => \N__23150\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__23150\,
            I => \N__23146\
        );

    \I__2686\ : CEMux
    port map (
            O => \N__23149\,
            I => \N__23143\
        );

    \I__2685\ : Span4Mux_h
    port map (
            O => \N__23146\,
            I => \N__23140\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__23143\,
            I => \N__23137\
        );

    \I__2683\ : Odrv4
    port map (
            O => \N__23140\,
            I => \sDAC_mem_29_1_sqmuxa\
        );

    \I__2682\ : Odrv12
    port map (
            O => \N__23137\,
            I => \sDAC_mem_29_1_sqmuxa\
        );

    \I__2681\ : InMux
    port map (
            O => \N__23132\,
            I => \un1_sTrigCounter_cry_11\
        );

    \I__2680\ : InMux
    port map (
            O => \N__23129\,
            I => \N__23125\
        );

    \I__2679\ : InMux
    port map (
            O => \N__23128\,
            I => \N__23122\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__23125\,
            I => \sTrigCounterZ0Z_13\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__23122\,
            I => \sTrigCounterZ0Z_13\
        );

    \I__2676\ : InMux
    port map (
            O => \N__23117\,
            I => \un1_sTrigCounter_cry_12\
        );

    \I__2675\ : InMux
    port map (
            O => \N__23114\,
            I => \N__23110\
        );

    \I__2674\ : InMux
    port map (
            O => \N__23113\,
            I => \N__23107\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__23110\,
            I => \sTrigCounterZ0Z_14\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__23107\,
            I => \sTrigCounterZ0Z_14\
        );

    \I__2671\ : InMux
    port map (
            O => \N__23102\,
            I => \un1_sTrigCounter_cry_13\
        );

    \I__2670\ : InMux
    port map (
            O => \N__23099\,
            I => \un1_sTrigCounter_cry_14\
        );

    \I__2669\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23092\
        );

    \I__2668\ : InMux
    port map (
            O => \N__23095\,
            I => \N__23089\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__23092\,
            I => \sTrigCounterZ0Z_15\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__23089\,
            I => \sTrigCounterZ0Z_15\
        );

    \I__2665\ : SRMux
    port map (
            O => \N__23084\,
            I => \N__23080\
        );

    \I__2664\ : SRMux
    port map (
            O => \N__23083\,
            I => \N__23077\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__23080\,
            I => \N_82_i\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__23077\,
            I => \N_82_i\
        );

    \I__2661\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23068\
        );

    \I__2660\ : InMux
    port map (
            O => \N__23071\,
            I => \N__23065\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__23068\,
            I => \sTrigCounterZ0Z_4\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__23065\,
            I => \sTrigCounterZ0Z_4\
        );

    \I__2657\ : InMux
    port map (
            O => \N__23060\,
            I => \un1_sTrigCounter_cry_3\
        );

    \I__2656\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23053\
        );

    \I__2655\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23050\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__23053\,
            I => \sTrigCounterZ0Z_5\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__23050\,
            I => \sTrigCounterZ0Z_5\
        );

    \I__2652\ : InMux
    port map (
            O => \N__23045\,
            I => \un1_sTrigCounter_cry_4\
        );

    \I__2651\ : InMux
    port map (
            O => \N__23042\,
            I => \N__23038\
        );

    \I__2650\ : InMux
    port map (
            O => \N__23041\,
            I => \N__23035\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__23038\,
            I => \sTrigCounterZ0Z_6\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__23035\,
            I => \sTrigCounterZ0Z_6\
        );

    \I__2647\ : InMux
    port map (
            O => \N__23030\,
            I => \un1_sTrigCounter_cry_5\
        );

    \I__2646\ : InMux
    port map (
            O => \N__23027\,
            I => \N__23023\
        );

    \I__2645\ : InMux
    port map (
            O => \N__23026\,
            I => \N__23020\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__23023\,
            I => \sTrigCounterZ0Z_7\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__23020\,
            I => \sTrigCounterZ0Z_7\
        );

    \I__2642\ : InMux
    port map (
            O => \N__23015\,
            I => \un1_sTrigCounter_cry_6\
        );

    \I__2641\ : InMux
    port map (
            O => \N__23012\,
            I => \N__23008\
        );

    \I__2640\ : InMux
    port map (
            O => \N__23011\,
            I => \N__23005\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__23008\,
            I => \sTrigCounterZ0Z_8\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__23005\,
            I => \sTrigCounterZ0Z_8\
        );

    \I__2637\ : InMux
    port map (
            O => \N__23000\,
            I => \bfn_8_14_0_\
        );

    \I__2636\ : InMux
    port map (
            O => \N__22997\,
            I => \N__22993\
        );

    \I__2635\ : InMux
    port map (
            O => \N__22996\,
            I => \N__22990\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__22993\,
            I => \sTrigCounterZ0Z_9\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__22990\,
            I => \sTrigCounterZ0Z_9\
        );

    \I__2632\ : InMux
    port map (
            O => \N__22985\,
            I => \un1_sTrigCounter_cry_8\
        );

    \I__2631\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22978\
        );

    \I__2630\ : InMux
    port map (
            O => \N__22981\,
            I => \N__22975\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__22978\,
            I => \sTrigCounterZ0Z_10\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__22975\,
            I => \sTrigCounterZ0Z_10\
        );

    \I__2627\ : InMux
    port map (
            O => \N__22970\,
            I => \un1_sTrigCounter_cry_9\
        );

    \I__2626\ : InMux
    port map (
            O => \N__22967\,
            I => \N__22963\
        );

    \I__2625\ : InMux
    port map (
            O => \N__22966\,
            I => \N__22960\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__22963\,
            I => \sTrigCounterZ0Z_11\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__22960\,
            I => \sTrigCounterZ0Z_11\
        );

    \I__2622\ : InMux
    port map (
            O => \N__22955\,
            I => \un1_sTrigCounter_cry_10\
        );

    \I__2621\ : InMux
    port map (
            O => \N__22952\,
            I => \N__22948\
        );

    \I__2620\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22945\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__22948\,
            I => \sTrigCounterZ0Z_12\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__22945\,
            I => \sTrigCounterZ0Z_12\
        );

    \I__2617\ : InMux
    port map (
            O => \N__22940\,
            I => \N__22931\
        );

    \I__2616\ : InMux
    port map (
            O => \N__22939\,
            I => \N__22931\
        );

    \I__2615\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22931\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__22931\,
            I => \N__22928\
        );

    \I__2613\ : Odrv4
    port map (
            O => \N__22928\,
            I => \un10_trig_prev_cry_15_THRU_CO\
        );

    \I__2612\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22922\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__22922\,
            I => \N_178\
        );

    \I__2610\ : InMux
    port map (
            O => \N__22919\,
            I => \N__22916\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__22916\,
            I => \N__22913\
        );

    \I__2608\ : Span4Mux_h
    port map (
            O => \N__22913\,
            I => \N__22910\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__22910\,
            I => un1_scounter_i_0
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__22907\,
            I => \N_178_cascade_\
        );

    \I__2605\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22901\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__22901\,
            I => \N_96\
        );

    \I__2603\ : CascadeMux
    port map (
            O => \N__22898\,
            I => \N_77_cascade_\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__22895\,
            I => \N__22890\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__22894\,
            I => \N__22887\
        );

    \I__2600\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22880\
        );

    \I__2599\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22880\
        );

    \I__2598\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22880\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__22880\,
            I => \sPeriod_prevZ0\
        );

    \I__2596\ : CascadeMux
    port map (
            O => \N__22877\,
            I => \N__22873\
        );

    \I__2595\ : InMux
    port map (
            O => \N__22876\,
            I => \N__22870\
        );

    \I__2594\ : InMux
    port map (
            O => \N__22873\,
            I => \N__22867\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__22870\,
            I => un1_reset_rpi_inv_2_0
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__22867\,
            I => un1_reset_rpi_inv_2_0
        );

    \I__2591\ : InMux
    port map (
            O => \N__22862\,
            I => \un1_sTrigCounter_cry_0\
        );

    \I__2590\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22855\
        );

    \I__2589\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22852\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__22855\,
            I => \sTrigCounterZ0Z_2\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__22852\,
            I => \sTrigCounterZ0Z_2\
        );

    \I__2586\ : InMux
    port map (
            O => \N__22847\,
            I => \un1_sTrigCounter_cry_1\
        );

    \I__2585\ : InMux
    port map (
            O => \N__22844\,
            I => \N__22840\
        );

    \I__2584\ : InMux
    port map (
            O => \N__22843\,
            I => \N__22837\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__22840\,
            I => \sTrigCounterZ0Z_3\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__22837\,
            I => \sTrigCounterZ0Z_3\
        );

    \I__2581\ : InMux
    port map (
            O => \N__22832\,
            I => \un1_sTrigCounter_cry_2\
        );

    \I__2580\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22824\
        );

    \I__2579\ : InMux
    port map (
            O => \N__22828\,
            I => \N__22821\
        );

    \I__2578\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22818\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__22824\,
            I => \N__22813\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__22821\,
            I => \N__22813\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__22818\,
            I => \N__22810\
        );

    \I__2574\ : Span4Mux_v
    port map (
            O => \N__22813\,
            I => \N__22807\
        );

    \I__2573\ : Span12Mux_v
    port map (
            O => \N__22810\,
            I => \N__22802\
        );

    \I__2572\ : Sp12to4
    port map (
            O => \N__22807\,
            I => \N__22802\
        );

    \I__2571\ : Odrv12
    port map (
            O => \N__22802\,
            I => trig_rpi_c
        );

    \I__2570\ : InMux
    port map (
            O => \N__22799\,
            I => \N__22795\
        );

    \I__2569\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22792\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__22795\,
            I => \N__22789\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__22792\,
            I => \N__22786\
        );

    \I__2566\ : Span4Mux_v
    port map (
            O => \N__22789\,
            I => \N__22782\
        );

    \I__2565\ : Span4Mux_v
    port map (
            O => \N__22786\,
            I => \N__22779\
        );

    \I__2564\ : InMux
    port map (
            O => \N__22785\,
            I => \N__22776\
        );

    \I__2563\ : Sp12to4
    port map (
            O => \N__22782\,
            I => \N__22769\
        );

    \I__2562\ : Sp12to4
    port map (
            O => \N__22779\,
            I => \N__22769\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__22776\,
            I => \N__22769\
        );

    \I__2560\ : Odrv12
    port map (
            O => \N__22769\,
            I => trig_ext_c
        );

    \I__2559\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22763\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__22763\,
            I => \N__22759\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__22762\,
            I => \N__22755\
        );

    \I__2556\ : Span4Mux_v
    port map (
            O => \N__22759\,
            I => \N__22752\
        );

    \I__2555\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22749\
        );

    \I__2554\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22746\
        );

    \I__2553\ : Sp12to4
    port map (
            O => \N__22752\,
            I => \N__22739\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__22749\,
            I => \N__22739\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__22746\,
            I => \N__22739\
        );

    \I__2550\ : Span12Mux_h
    port map (
            O => \N__22739\,
            I => \N__22736\
        );

    \I__2549\ : Span12Mux_v
    port map (
            O => \N__22736\,
            I => \N__22733\
        );

    \I__2548\ : Span12Mux_h
    port map (
            O => \N__22733\,
            I => \N__22730\
        );

    \I__2547\ : Odrv12
    port map (
            O => \N__22730\,
            I => trig_ft_c
        );

    \I__2546\ : InMux
    port map (
            O => \N__22727\,
            I => \N__22723\
        );

    \I__2545\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22720\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__22723\,
            I => \N__22717\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__22720\,
            I => \N__22711\
        );

    \I__2542\ : Span4Mux_v
    port map (
            O => \N__22717\,
            I => \N__22711\
        );

    \I__2541\ : InMux
    port map (
            O => \N__22716\,
            I => \N__22708\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__22711\,
            I => \trig_prevZ0\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__22708\,
            I => \trig_prevZ0\
        );

    \I__2538\ : CascadeMux
    port map (
            O => \N__22703\,
            I => \g3_0_cascade_\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__22700\,
            I => \sAddress_RNI70I7Z0Z_1_cascade_\
        );

    \I__2536\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22694\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__22694\,
            I => g1_i_a4_0_0
        );

    \I__2534\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22688\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__22688\,
            I => \N_8_mux\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__22685\,
            I => \N_319_cascade_\
        );

    \I__2531\ : CEMux
    port map (
            O => \N__22682\,
            I => \N__22679\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__2529\ : Span4Mux_v
    port map (
            O => \N__22676\,
            I => \N__22673\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__22673\,
            I => \sAddress_RNI9IH12_2Z0Z_1\
        );

    \I__2527\ : InMux
    port map (
            O => \N__22670\,
            I => \N__22667\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__22667\,
            I => \N__22664\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__22664\,
            I => \N__22659\
        );

    \I__2524\ : InMux
    port map (
            O => \N__22663\,
            I => \N__22656\
        );

    \I__2523\ : InMux
    port map (
            O => \N__22662\,
            I => \N__22653\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__22659\,
            I => \spi_slave_inst.rx_done_reg2_iZ0\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__22656\,
            I => \spi_slave_inst.rx_done_reg2_iZ0\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__22653\,
            I => \spi_slave_inst.rx_done_reg2_iZ0\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__22646\,
            I => \N__22643\
        );

    \I__2518\ : InMux
    port map (
            O => \N__22643\,
            I => \N__22640\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__22640\,
            I => \N__22637\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__22637\,
            I => \spi_slave_inst.rx_done_reg3_iZ0\
        );

    \I__2515\ : InMux
    port map (
            O => \N__22634\,
            I => \N__22631\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__22631\,
            I => \N__22628\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__22628\,
            I => \spi_slave_inst.rx_ready_i_RNOZ0Z_0\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__22625\,
            I => \sPointer_RNI5LBD1Z0Z_0_cascade_\
        );

    \I__2511\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22616\
        );

    \I__2510\ : InMux
    port map (
            O => \N__22621\,
            I => \N__22616\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__22616\,
            I => \sDAC_mem_17_1_sqmuxa_0_a2_0_a2_1_0\
        );

    \I__2508\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22604\
        );

    \I__2507\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22604\
        );

    \I__2506\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22599\
        );

    \I__2505\ : InMux
    port map (
            O => \N__22610\,
            I => \N__22599\
        );

    \I__2504\ : InMux
    port map (
            O => \N__22609\,
            I => \N__22596\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__22604\,
            I => \sAddressZ0Z_4\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__22599\,
            I => \sAddressZ0Z_4\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__22596\,
            I => \sAddressZ0Z_4\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__22589\,
            I => \sAddress_RNIP2UK1Z0Z_4_cascade_\
        );

    \I__2499\ : InMux
    port map (
            O => \N__22586\,
            I => \N__22583\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__22583\,
            I => \N__22580\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__22580\,
            I => \N__22577\
        );

    \I__2496\ : Span4Mux_v
    port map (
            O => \N__22577\,
            I => \N__22573\
        );

    \I__2495\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22570\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__22573\,
            I => \spi_slave_inst.rx_done_neg_sclk_iZ0\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__22570\,
            I => \spi_slave_inst.rx_done_neg_sclk_iZ0\
        );

    \I__2492\ : CEMux
    port map (
            O => \N__22565\,
            I => \N__22562\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__22562\,
            I => \N__22559\
        );

    \I__2490\ : Odrv12
    port map (
            O => \N__22559\,
            I => \spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541\
        );

    \I__2489\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22550\
        );

    \I__2488\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22550\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__22550\,
            I => \spi_slave_inst.rx_done_reg1_iZ0\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__22547\,
            I => \N_344_cascade_\
        );

    \I__2485\ : CEMux
    port map (
            O => \N__22544\,
            I => \N__22541\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__22541\,
            I => \N__22538\
        );

    \I__2483\ : Span4Mux_h
    port map (
            O => \N__22538\,
            I => \N__22535\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__22535\,
            I => \sDAC_mem_35_1_sqmuxa\
        );

    \I__2481\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22529\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__22529\,
            I => \sEESingleCont_RNOZ0Z_0\
        );

    \I__2479\ : InMux
    port map (
            O => \N__22526\,
            I => \N__22523\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__22523\,
            I => \N__22519\
        );

    \I__2477\ : InMux
    port map (
            O => \N__22522\,
            I => \N__22516\
        );

    \I__2476\ : Span4Mux_v
    port map (
            O => \N__22519\,
            I => \N__22513\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__22516\,
            I => \sEESingleContZ0\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__22513\,
            I => \sEESingleContZ0\
        );

    \I__2473\ : InMux
    port map (
            O => \N__22508\,
            I => \N__22505\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__22505\,
            I => \N_1631\
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__2470\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__22496\,
            I => \sEETrigInternal_3_iv_0_0_i_0\
        );

    \I__2468\ : CEMux
    port map (
            O => \N__22493\,
            I => \N__22490\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__22490\,
            I => \N__22487\
        );

    \I__2466\ : Odrv12
    port map (
            O => \N__22487\,
            I => \sDAC_mem_11_1_sqmuxa\
        );

    \I__2465\ : InMux
    port map (
            O => \N__22484\,
            I => \N__22481\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__22481\,
            I => \N__22477\
        );

    \I__2463\ : InMux
    port map (
            O => \N__22480\,
            I => \N__22474\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__22477\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__22474\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0\
        );

    \I__2460\ : InMux
    port map (
            O => \N__22469\,
            I => \N__22466\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__22466\,
            I => \N__22462\
        );

    \I__2458\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22459\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__22462\,
            I => \N__22454\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__22459\,
            I => \N__22454\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__22454\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1\
        );

    \I__2454\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22447\
        );

    \I__2453\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22444\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__22447\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__22444\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2\
        );

    \I__2450\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22435\
        );

    \I__2449\ : InMux
    port map (
            O => \N__22438\,
            I => \N__22432\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__22435\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__22432\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3\
        );

    \I__2446\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22423\
        );

    \I__2445\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22420\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__22423\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__22420\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4\
        );

    \I__2442\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22411\
        );

    \I__2441\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22408\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__22411\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__22408\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5\
        );

    \I__2438\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22399\
        );

    \I__2437\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22396\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__22399\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__22396\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6\
        );

    \I__2434\ : InMux
    port map (
            O => \N__22391\,
            I => \N__22388\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__22388\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__22385\,
            I => \N__22382\
        );

    \I__2431\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22378\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__22381\,
            I => \N__22375\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__22378\,
            I => \N__22372\
        );

    \I__2428\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22369\
        );

    \I__2427\ : Odrv4
    port map (
            O => \N__22372\,
            I => un3_trig_0
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__22369\,
            I => un3_trig_0
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__22364\,
            I => \N__22361\
        );

    \I__2424\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22358\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__22358\,
            I => \sEEADC_freqZ0Z_5\
        );

    \I__2422\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__22352\,
            I => \N__22349\
        );

    \I__2420\ : Span4Mux_v
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__2419\ : Sp12to4
    port map (
            O => \N__22346\,
            I => \N__22343\
        );

    \I__2418\ : Span12Mux_h
    port map (
            O => \N__22343\,
            I => \N__22340\
        );

    \I__2417\ : Odrv12
    port map (
            O => \N__22340\,
            I => spi_mosi_rpi_c
        );

    \I__2416\ : InMux
    port map (
            O => \N__22337\,
            I => \N__22334\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__2414\ : Span4Mux_v
    port map (
            O => \N__22331\,
            I => \N__22328\
        );

    \I__2413\ : Span4Mux_h
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__2412\ : Sp12to4
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__2411\ : Span12Mux_h
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__2410\ : Odrv12
    port map (
            O => \N__22319\,
            I => spi_mosi_ft_c
        );

    \I__2409\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__22313\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__2406\ : InMux
    port map (
            O => \N__22307\,
            I => \N__22304\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__22304\,
            I => un10_trig_prev_14
        );

    \I__2404\ : InMux
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__22298\,
            I => \sTrigCounter_i_14\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__22295\,
            I => \N__22292\
        );

    \I__2401\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22289\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__22289\,
            I => un10_trig_prev_15
        );

    \I__2399\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22283\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__22283\,
            I => \sTrigCounter_i_15\
        );

    \I__2397\ : InMux
    port map (
            O => \N__22280\,
            I => \bfn_7_14_0_\
        );

    \I__2396\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__22274\,
            I => \N_173\
        );

    \I__2394\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22268\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__22268\,
            I => \sEEADC_freqZ0Z_4\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__22265\,
            I => \N__22262\
        );

    \I__2391\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__22259\,
            I => un10_trig_prev_6
        );

    \I__2389\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22253\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__22253\,
            I => \sTrigCounter_i_6\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__2386\ : InMux
    port map (
            O => \N__22247\,
            I => \N__22244\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__22244\,
            I => un10_trig_prev_7
        );

    \I__2384\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22238\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__22238\,
            I => \sTrigCounter_i_7\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__22235\,
            I => \N__22232\
        );

    \I__2381\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22229\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__22229\,
            I => un10_trig_prev_8
        );

    \I__2379\ : InMux
    port map (
            O => \N__22226\,
            I => \N__22223\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__22223\,
            I => \sTrigCounter_i_8\
        );

    \I__2377\ : CascadeMux
    port map (
            O => \N__22220\,
            I => \N__22217\
        );

    \I__2376\ : InMux
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__22214\,
            I => un10_trig_prev_9
        );

    \I__2374\ : InMux
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__22208\,
            I => \sTrigCounter_i_9\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__2371\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__22199\,
            I => un10_trig_prev_10
        );

    \I__2369\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__22193\,
            I => \sTrigCounter_i_10\
        );

    \I__2367\ : CascadeMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__2366\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__22184\,
            I => un10_trig_prev_11
        );

    \I__2364\ : InMux
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__22178\,
            I => \sTrigCounter_i_11\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__2361\ : InMux
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__22169\,
            I => un10_trig_prev_12
        );

    \I__2359\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22163\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__22163\,
            I => \sTrigCounter_i_12\
        );

    \I__2357\ : CascadeMux
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__2356\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22154\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__22154\,
            I => un10_trig_prev_13
        );

    \I__2354\ : InMux
    port map (
            O => \N__22151\,
            I => \N__22148\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__22148\,
            I => \sTrigCounter_i_13\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__22145\,
            I => \N__22141\
        );

    \I__2351\ : InMux
    port map (
            O => \N__22144\,
            I => \N__22138\
        );

    \I__2350\ : InMux
    port map (
            O => \N__22141\,
            I => \N__22135\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__22138\,
            I => un8_trig_prev_0
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__22135\,
            I => un8_trig_prev_0
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__22130\,
            I => \N__22127\
        );

    \I__2346\ : InMux
    port map (
            O => \N__22127\,
            I => \N__22124\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__22124\,
            I => un10_trig_prev_0
        );

    \I__2344\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22118\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__22118\,
            I => \sTrigCounter_i_0\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__22115\,
            I => \N__22112\
        );

    \I__2341\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22109\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__22109\,
            I => un10_trig_prev_1
        );

    \I__2339\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22103\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__22103\,
            I => \sTrigCounter_i_1\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__2336\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22094\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__22094\,
            I => un10_trig_prev_2
        );

    \I__2334\ : InMux
    port map (
            O => \N__22091\,
            I => \N__22088\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__22088\,
            I => \sTrigCounter_i_2\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__2331\ : InMux
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__22079\,
            I => un10_trig_prev_3
        );

    \I__2329\ : InMux
    port map (
            O => \N__22076\,
            I => \N__22073\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__22073\,
            I => \sTrigCounter_i_3\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__22070\,
            I => \N__22067\
        );

    \I__2326\ : InMux
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__22064\,
            I => un10_trig_prev_4
        );

    \I__2324\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22058\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__22058\,
            I => \sTrigCounter_i_4\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__22055\,
            I => \N__22052\
        );

    \I__2321\ : InMux
    port map (
            O => \N__22052\,
            I => \N__22049\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__22049\,
            I => un10_trig_prev_5
        );

    \I__2319\ : InMux
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__22043\,
            I => \sTrigCounter_i_5\
        );

    \I__2317\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22036\
        );

    \I__2316\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22033\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__22036\,
            I => \N__22030\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__22033\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2313\ : Odrv4
    port map (
            O => \N__22030\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2312\ : InMux
    port map (
            O => \N__22025\,
            I => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1\
        );

    \I__2311\ : InMux
    port map (
            O => \N__22022\,
            I => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2\
        );

    \I__2310\ : InMux
    port map (
            O => \N__22019\,
            I => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3\
        );

    \I__2309\ : InMux
    port map (
            O => \N__22016\,
            I => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4\
        );

    \I__2308\ : InMux
    port map (
            O => \N__22013\,
            I => \N__22009\
        );

    \I__2307\ : InMux
    port map (
            O => \N__22012\,
            I => \N__22006\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__22009\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__22006\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__2304\ : InMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__2302\ : Span4Mux_h
    port map (
            O => \N__21995\,
            I => \N__21988\
        );

    \I__2301\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21983\
        );

    \I__2300\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21983\
        );

    \I__2299\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21978\
        );

    \I__2298\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21978\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__21988\,
            I => spi_mosi_ready
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__21983\,
            I => spi_mosi_ready
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__21978\,
            I => spi_mosi_ready
        );

    \I__2294\ : InMux
    port map (
            O => \N__21971\,
            I => \N__21967\
        );

    \I__2293\ : InMux
    port map (
            O => \N__21970\,
            I => \N__21964\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__21967\,
            I => \spi_mosi_ready_prevZ0\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__21964\,
            I => \spi_mosi_ready_prevZ0\
        );

    \I__2290\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21955\
        );

    \I__2289\ : InMux
    port map (
            O => \N__21958\,
            I => \N__21952\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__21955\,
            I => \spi_mosi_ready_prevZ0Z2\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__21952\,
            I => \spi_mosi_ready_prevZ0Z2\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__2285\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__21941\,
            I => \spi_mosi_ready_prevZ0Z3\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__21938\,
            I => \N_346_i_cascade_\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__21935\,
            I => \un1_spointer11_8_0_0_a2_1_cascade_\
        );

    \I__2281\ : CEMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__2279\ : Span4Mux_v
    port map (
            O => \N__21926\,
            I => \N__21923\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__21923\,
            I => \sAddress_RNI7G5E2Z0Z_6\
        );

    \I__2277\ : InMux
    port map (
            O => \N__21920\,
            I => \N__21910\
        );

    \I__2276\ : InMux
    port map (
            O => \N__21919\,
            I => \N__21910\
        );

    \I__2275\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21910\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__21917\,
            I => \N__21907\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__21910\,
            I => \N__21904\
        );

    \I__2272\ : InMux
    port map (
            O => \N__21907\,
            I => \N__21901\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__21904\,
            I => \N__21896\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__21901\,
            I => \N__21896\
        );

    \I__2269\ : Span4Mux_h
    port map (
            O => \N__21896\,
            I => \N__21893\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__21893\,
            I => \sAddressZ0Z_7\
        );

    \I__2267\ : InMux
    port map (
            O => \N__21890\,
            I => \N__21881\
        );

    \I__2266\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21881\
        );

    \I__2265\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21881\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__21881\,
            I => \N__21877\
        );

    \I__2263\ : InMux
    port map (
            O => \N__21880\,
            I => \N__21874\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__21877\,
            I => \N__21869\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__21874\,
            I => \N__21869\
        );

    \I__2260\ : Span4Mux_h
    port map (
            O => \N__21869\,
            I => \N__21866\
        );

    \I__2259\ : Odrv4
    port map (
            O => \N__21866\,
            I => \sAddressZ0Z_6\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__21863\,
            I => \N__21860\
        );

    \I__2257\ : InMux
    port map (
            O => \N__21860\,
            I => \N__21856\
        );

    \I__2256\ : InMux
    port map (
            O => \N__21859\,
            I => \N__21853\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__21856\,
            I => \N__21850\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__21853\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__21850\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__2252\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21841\
        );

    \I__2251\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21838\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__21841\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__21838\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__2248\ : InMux
    port map (
            O => \N__21833\,
            I => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__21830\,
            I => \N_316_cascade_\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__21827\,
            I => \N_317_cascade_\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__21824\,
            I => \sAddress_RNI8U0V1Z0Z_1_cascade_\
        );

    \I__2244\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21818\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__21818\,
            I => \sAddress_RNI8U0V1Z0Z_1\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__21815\,
            I => \N_454_cascade_\
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__2240\ : InMux
    port map (
            O => \N__21809\,
            I => \N__21806\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__21806\,
            I => \sEETrigCounterZ0Z_9\
        );

    \I__2238\ : InMux
    port map (
            O => \N__21803\,
            I => \N__21800\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__21800\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11\
        );

    \I__2236\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__2234\ : Span4Mux_v
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__21788\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1\
        );

    \I__2232\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__21782\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5\
        );

    \I__2230\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__21776\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13\
        );

    \I__2228\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__21770\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14\
        );

    \I__2226\ : InMux
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__21761\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0\
        );

    \I__2223\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__21755\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_6\
        );

    \I__2221\ : InMux
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__21749\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_5\
        );

    \I__2219\ : InMux
    port map (
            O => \N__21746\,
            I => un8_trig_prev_0_cry_13
        );

    \I__2218\ : InMux
    port map (
            O => \N__21743\,
            I => un8_trig_prev_0_cry_14
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__2216\ : InMux
    port map (
            O => \N__21737\,
            I => \N__21734\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__21734\,
            I => \sEETrigCounterZ0Z_10\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__2213\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21725\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__21725\,
            I => \sEETrigCounterZ0Z_11\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__21722\,
            I => \N__21719\
        );

    \I__2210\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21716\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__21716\,
            I => \sEETrigCounterZ0Z_12\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__21713\,
            I => \N__21710\
        );

    \I__2207\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21707\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__21707\,
            I => \sEETrigCounterZ0Z_13\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__2204\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__21698\,
            I => \sEETrigCounterZ0Z_14\
        );

    \I__2202\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21692\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__21692\,
            I => \sEETrigCounterZ0Z_15\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__21689\,
            I => \N__21686\
        );

    \I__2199\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21683\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__21683\,
            I => \sEETrigCounterZ0Z_8\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__2196\ : InMux
    port map (
            O => \N__21677\,
            I => \N__21674\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__21674\,
            I => \sEETrigCounterZ0Z_5\
        );

    \I__2194\ : InMux
    port map (
            O => \N__21671\,
            I => un8_trig_prev_0_cry_4
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__2192\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__21662\,
            I => \sEETrigCounterZ0Z_6\
        );

    \I__2190\ : InMux
    port map (
            O => \N__21659\,
            I => un8_trig_prev_0_cry_5
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__2188\ : InMux
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__21650\,
            I => \sEETrigCounterZ0Z_7\
        );

    \I__2186\ : InMux
    port map (
            O => \N__21647\,
            I => un8_trig_prev_0_cry_6
        );

    \I__2185\ : InMux
    port map (
            O => \N__21644\,
            I => \bfn_6_13_0_\
        );

    \I__2184\ : InMux
    port map (
            O => \N__21641\,
            I => un8_trig_prev_0_cry_8
        );

    \I__2183\ : InMux
    port map (
            O => \N__21638\,
            I => un8_trig_prev_0_cry_9
        );

    \I__2182\ : InMux
    port map (
            O => \N__21635\,
            I => un8_trig_prev_0_cry_10
        );

    \I__2181\ : InMux
    port map (
            O => \N__21632\,
            I => un8_trig_prev_0_cry_11
        );

    \I__2180\ : InMux
    port map (
            O => \N__21629\,
            I => un8_trig_prev_0_cry_12
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__21626\,
            I => \N__21623\
        );

    \I__2178\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21620\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__21620\,
            I => \sEETrigCounterZ0Z_1\
        );

    \I__2176\ : InMux
    port map (
            O => \N__21617\,
            I => un8_trig_prev_0_cry_0
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__2174\ : InMux
    port map (
            O => \N__21611\,
            I => \N__21608\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__21608\,
            I => \sEETrigCounterZ0Z_2\
        );

    \I__2172\ : InMux
    port map (
            O => \N__21605\,
            I => un8_trig_prev_0_cry_1
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__21602\,
            I => \N__21599\
        );

    \I__2170\ : InMux
    port map (
            O => \N__21599\,
            I => \N__21596\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__21596\,
            I => \sEETrigCounterZ0Z_3\
        );

    \I__2168\ : InMux
    port map (
            O => \N__21593\,
            I => un8_trig_prev_0_cry_2
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__21590\,
            I => \N__21587\
        );

    \I__2166\ : InMux
    port map (
            O => \N__21587\,
            I => \N__21584\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__21584\,
            I => \sEETrigCounterZ0Z_4\
        );

    \I__2164\ : InMux
    port map (
            O => \N__21581\,
            I => un8_trig_prev_0_cry_3
        );

    \I__2163\ : InMux
    port map (
            O => \N__21578\,
            I => \N__21574\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__21577\,
            I => \N__21571\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__21574\,
            I => \N__21567\
        );

    \I__2160\ : InMux
    port map (
            O => \N__21571\,
            I => \N__21564\
        );

    \I__2159\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21560\
        );

    \I__2158\ : Span4Mux_v
    port map (
            O => \N__21567\,
            I => \N__21555\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__21564\,
            I => \N__21555\
        );

    \I__2156\ : InMux
    port map (
            O => \N__21563\,
            I => \N__21552\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__21560\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__21555\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__21552\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__2152\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21541\
        );

    \I__2151\ : InMux
    port map (
            O => \N__21544\,
            I => \N__21538\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__21541\,
            I => \N__21535\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__21538\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__2148\ : Odrv12
    port map (
            O => \N__21535\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__21530\,
            I => \N__21527\
        );

    \I__2146\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21523\
        );

    \I__2145\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21520\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__21523\,
            I => \N__21517\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__21520\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__2142\ : Odrv12
    port map (
            O => \N__21517\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__2141\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21508\
        );

    \I__2140\ : InMux
    port map (
            O => \N__21511\,
            I => \N__21505\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__21508\,
            I => \N__21498\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__21505\,
            I => \N__21498\
        );

    \I__2137\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21495\
        );

    \I__2136\ : InMux
    port map (
            O => \N__21503\,
            I => \N__21491\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__21498\,
            I => \N__21486\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__21495\,
            I => \N__21486\
        );

    \I__2133\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21483\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__21491\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__2131\ : Odrv4
    port map (
            O => \N__21486\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__21483\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__2129\ : InMux
    port map (
            O => \N__21476\,
            I => \N__21472\
        );

    \I__2128\ : InMux
    port map (
            O => \N__21475\,
            I => \N__21469\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__21472\,
            I => \N__21466\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__21469\,
            I => \N__21463\
        );

    \I__2125\ : Odrv4
    port map (
            O => \N__21466\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__21463\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3\
        );

    \I__2123\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21454\
        );

    \I__2122\ : InMux
    port map (
            O => \N__21457\,
            I => \N__21451\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__21454\,
            I => \spi_mosi_ready64_prevZ0Z2\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__21451\,
            I => \spi_mosi_ready64_prevZ0Z2\
        );

    \I__2119\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21442\
        );

    \I__2118\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21439\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__21442\,
            I => \spi_mosi_ready64_prevZ0\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__21439\,
            I => \spi_mosi_ready64_prevZ0\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__21434\,
            I => \N__21431\
        );

    \I__2114\ : InMux
    port map (
            O => \N__21431\,
            I => \N__21428\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__21428\,
            I => \spi_mosi_ready64_prevZ0Z3\
        );

    \I__2112\ : CascadeMux
    port map (
            O => \N__21425\,
            I => \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_\
        );

    \I__2111\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21418\
        );

    \I__2110\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21412\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__21418\,
            I => \N__21409\
        );

    \I__2108\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21406\
        );

    \I__2107\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21403\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__21415\,
            I => \N__21397\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__21412\,
            I => \N__21394\
        );

    \I__2104\ : Span4Mux_h
    port map (
            O => \N__21409\,
            I => \N__21387\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__21406\,
            I => \N__21387\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__21403\,
            I => \N__21387\
        );

    \I__2101\ : InMux
    port map (
            O => \N__21402\,
            I => \N__21384\
        );

    \I__2100\ : InMux
    port map (
            O => \N__21401\,
            I => \N__21379\
        );

    \I__2099\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21379\
        );

    \I__2098\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21376\
        );

    \I__2097\ : Odrv12
    port map (
            O => \N__21394\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__21387\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__21384\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__21379\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__21376\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2092\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21362\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__21362\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO\
        );

    \I__2090\ : InMux
    port map (
            O => \N__21359\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1\
        );

    \I__2089\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21353\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__21353\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO\
        );

    \I__2087\ : InMux
    port map (
            O => \N__21350\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2\
        );

    \I__2086\ : InMux
    port map (
            O => \N__21347\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3\
        );

    \I__2085\ : InMux
    port map (
            O => \N__21344\,
            I => \bfn_6_8_0_\
        );

    \I__2084\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21338\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__21338\,
            I => \N__21335\
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__21335\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__21332\,
            I => \N__21328\
        );

    \I__2080\ : InMux
    port map (
            O => \N__21331\,
            I => \N__21321\
        );

    \I__2079\ : InMux
    port map (
            O => \N__21328\,
            I => \N__21321\
        );

    \I__2078\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21316\
        );

    \I__2077\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21316\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__21321\,
            I => \N__21313\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__21316\,
            I => \N__21310\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__21313\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__21310\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__21305\,
            I => \N__21301\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__21304\,
            I => \N__21298\
        );

    \I__2070\ : InMux
    port map (
            O => \N__21301\,
            I => \N__21291\
        );

    \I__2069\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21291\
        );

    \I__2068\ : CEMux
    port map (
            O => \N__21297\,
            I => \N__21288\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__21296\,
            I => \N__21285\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__21291\,
            I => \N__21277\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__21288\,
            I => \N__21277\
        );

    \I__2064\ : InMux
    port map (
            O => \N__21285\,
            I => \N__21274\
        );

    \I__2063\ : InMux
    port map (
            O => \N__21284\,
            I => \N__21269\
        );

    \I__2062\ : InMux
    port map (
            O => \N__21283\,
            I => \N__21269\
        );

    \I__2061\ : InMux
    port map (
            O => \N__21282\,
            I => \N__21266\
        );

    \I__2060\ : Span4Mux_v
    port map (
            O => \N__21277\,
            I => \N__21263\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__21274\,
            I => \spi_master_inst.o_sclk_RNIH6AC\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__21269\,
            I => \spi_master_inst.o_sclk_RNIH6AC\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__21266\,
            I => \spi_master_inst.o_sclk_RNIH6AC\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__21263\,
            I => \spi_master_inst.o_sclk_RNIH6AC\
        );

    \I__2055\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21250\
        );

    \I__2054\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21247\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__21250\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__21247\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2\
        );

    \I__2051\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21239\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__21239\,
            I => \spi_master_inst.spi_data_path_u1.N_1411\
        );

    \I__2049\ : InMux
    port map (
            O => \N__21236\,
            I => \N__21233\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__21233\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13\
        );

    \I__2047\ : InMux
    port map (
            O => \N__21230\,
            I => \N__21227\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__21227\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14\
        );

    \I__2045\ : InMux
    port map (
            O => \N__21224\,
            I => \N__21221\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__21221\,
            I => \spi_master_inst.spi_data_path_u1.N_1418\
        );

    \I__2043\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21212\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__21212\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6\
        );

    \I__2040\ : InMux
    port map (
            O => \N__21209\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0\
        );

    \I__2039\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21202\
        );

    \I__2038\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21199\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__21202\,
            I => \N__21194\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__21199\,
            I => \N__21194\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__21194\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6\
        );

    \I__2034\ : InMux
    port map (
            O => \N__21191\,
            I => \N__21187\
        );

    \I__2033\ : InMux
    port map (
            O => \N__21190\,
            I => \N__21184\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__21187\,
            I => \N__21181\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__21184\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__21181\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__21176\,
            I => \N__21173\
        );

    \I__2028\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21169\
        );

    \I__2027\ : InMux
    port map (
            O => \N__21172\,
            I => \N__21166\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__21169\,
            I => \N__21163\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__21166\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7\
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__21163\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7\
        );

    \I__2023\ : InMux
    port map (
            O => \N__21158\,
            I => \N__21154\
        );

    \I__2022\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21151\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__21154\,
            I => \N__21148\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__21151\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__21148\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4\
        );

    \I__2018\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__21140\,
            I => \N__21136\
        );

    \I__2016\ : InMux
    port map (
            O => \N__21139\,
            I => \N__21133\
        );

    \I__2015\ : Span4Mux_h
    port map (
            O => \N__21136\,
            I => \N__21130\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__21133\,
            I => \N__21127\
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__21130\,
            I => \spi_master_inst.sclk_gen_u0.N_1737\
        );

    \I__2012\ : Odrv12
    port map (
            O => \N__21127\,
            I => \spi_master_inst.sclk_gen_u0.N_1737\
        );

    \I__2011\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21119\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__2009\ : Span4Mux_h
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__21113\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__21110\,
            I => \spi_master_inst.sclk_gen_u0.N_1737_cascade_\
        );

    \I__2006\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21104\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__21104\,
            I => \N__21100\
        );

    \I__2004\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21097\
        );

    \I__2003\ : Span4Mux_h
    port map (
            O => \N__21100\,
            I => \N__21094\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__21097\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0\
        );

    \I__2001\ : Odrv4
    port map (
            O => \N__21094\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0\
        );

    \I__2000\ : InMux
    port map (
            O => \N__21089\,
            I => \N__21083\
        );

    \I__1999\ : InMux
    port map (
            O => \N__21088\,
            I => \N__21083\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__21083\,
            I => \N__21080\
        );

    \I__1997\ : Odrv12
    port map (
            O => \N__21080\,
            I => \spi_master_inst.sclk_gen_u0.N_1540\
        );

    \I__1996\ : InMux
    port map (
            O => \N__21077\,
            I => \N__21073\
        );

    \I__1995\ : InMux
    port map (
            O => \N__21076\,
            I => \N__21070\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__21073\,
            I => \N__21067\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__21070\,
            I => \N__21059\
        );

    \I__1992\ : Span12Mux_s8_h
    port map (
            O => \N__21067\,
            I => \N__21059\
        );

    \I__1991\ : InMux
    port map (
            O => \N__21066\,
            I => \N__21056\
        );

    \I__1990\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21051\
        );

    \I__1989\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21051\
        );

    \I__1988\ : Odrv12
    port map (
            O => \N__21059\,
            I => \spi_master_inst.ss_start_i\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__21056\,
            I => \spi_master_inst.ss_start_i\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__21051\,
            I => \spi_master_inst.ss_start_i\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__21044\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__21041\,
            I => \spi_master_inst.spi_data_path_u1.N_1421_cascade_\
        );

    \I__1983\ : InMux
    port map (
            O => \N__21038\,
            I => \N__21035\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__21035\,
            I => \spi_master_inst.spi_data_path_u1.N_1422\
        );

    \I__1981\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21029\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__21029\,
            I => \N__21024\
        );

    \I__1979\ : InMux
    port map (
            O => \N__21028\,
            I => \N__21021\
        );

    \I__1978\ : InMux
    port map (
            O => \N__21027\,
            I => \N__21018\
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__21024\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__21021\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__21018\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2\
        );

    \I__1974\ : InMux
    port map (
            O => \N__21011\,
            I => \N__21007\
        );

    \I__1973\ : InMux
    port map (
            O => \N__21010\,
            I => \N__21003\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__21007\,
            I => \N__21000\
        );

    \I__1971\ : InMux
    port map (
            O => \N__21006\,
            I => \N__20997\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__21003\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__21000\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__20997\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__1966\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__20984\,
            I => \N__20979\
        );

    \I__1964\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20976\
        );

    \I__1963\ : InMux
    port map (
            O => \N__20982\,
            I => \N__20973\
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__20979\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__20976\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__20973\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3\
        );

    \I__1959\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20962\
        );

    \I__1958\ : InMux
    port map (
            O => \N__20965\,
            I => \N__20958\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__20962\,
            I => \N__20955\
        );

    \I__1956\ : InMux
    port map (
            O => \N__20961\,
            I => \N__20952\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__20958\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__20955\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__20952\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4\
        );

    \I__1952\ : InMux
    port map (
            O => \N__20945\,
            I => \N__20942\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__20942\,
            I => \spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1\
        );

    \I__1950\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20936\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__20936\,
            I => \N__20932\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__20935\,
            I => \N__20928\
        );

    \I__1947\ : Span4Mux_h
    port map (
            O => \N__20932\,
            I => \N__20925\
        );

    \I__1946\ : InMux
    port map (
            O => \N__20931\,
            I => \N__20922\
        );

    \I__1945\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20919\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__20925\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__20922\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__20919\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7\
        );

    \I__1941\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20909\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__1939\ : Span4Mux_h
    port map (
            O => \N__20906\,
            I => \N__20901\
        );

    \I__1938\ : InMux
    port map (
            O => \N__20905\,
            I => \N__20898\
        );

    \I__1937\ : InMux
    port map (
            O => \N__20904\,
            I => \N__20895\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__20901\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__20898\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__20895\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6\
        );

    \I__1933\ : IoInMux
    port map (
            O => \N__20888\,
            I => \N__20885\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__20885\,
            I => \N__20882\
        );

    \I__1931\ : Span4Mux_s2_v
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__1930\ : Sp12to4
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__1929\ : Span12Mux_s8_h
    port map (
            O => \N__20876\,
            I => \N__20872\
        );

    \I__1928\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20869\
        );

    \I__1927\ : Odrv12
    port map (
            O => \N__20872\,
            I => \DAC_sclk_c\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__20869\,
            I => \DAC_sclk_c\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__20864\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_cascade_\
        );

    \I__1924\ : InMux
    port map (
            O => \N__20861\,
            I => \N__20857\
        );

    \I__1923\ : InMux
    port map (
            O => \N__20860\,
            I => \N__20854\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__20857\,
            I => \spi_master_inst.sclk_gen_u0.N_36\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__20854\,
            I => \spi_master_inst.sclk_gen_u0.N_36\
        );

    \I__1920\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__20846\,
            I => \spi_master_inst.sclk_gen_u0.N_5\
        );

    \I__1918\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20839\
        );

    \I__1917\ : InMux
    port map (
            O => \N__20842\,
            I => \N__20835\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__20839\,
            I => \N__20832\
        );

    \I__1915\ : InMux
    port map (
            O => \N__20838\,
            I => \N__20829\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__20835\,
            I => \spi_master_inst.sclk_gen_u0.N_150_0\
        );

    \I__1913\ : Odrv4
    port map (
            O => \N__20832\,
            I => \spi_master_inst.sclk_gen_u0.N_150_0\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__20829\,
            I => \spi_master_inst.sclk_gen_u0.N_150_0\
        );

    \I__1911\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20819\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__20819\,
            I => \spi_master_inst.sclk_gen_u0.N_48\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__20816\,
            I => \spi_master_inst.spi_data_path_u1.N_1414_cascade_\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__20813\,
            I => \spi_master_inst.spi_data_path_u1.N_1415_cascade_\
        );

    \I__1907\ : IoInMux
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__20807\,
            I => \N__20804\
        );

    \I__1905\ : IoSpan4Mux
    port map (
            O => \N__20804\,
            I => \N__20801\
        );

    \I__1904\ : Span4Mux_s3_v
    port map (
            O => \N__20801\,
            I => \N__20798\
        );

    \I__1903\ : Span4Mux_v
    port map (
            O => \N__20798\,
            I => \N__20795\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__20795\,
            I => \DAC_mosi_c\
        );

    \I__1901\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20789\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__20789\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1\
        );

    \I__1899\ : InMux
    port map (
            O => \N__20786\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_4\
        );

    \I__1898\ : InMux
    port map (
            O => \N__20783\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_5\
        );

    \I__1897\ : InMux
    port map (
            O => \N__20780\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_6\
        );

    \I__1896\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__20774\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3\
        );

    \I__1894\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20766\
        );

    \I__1893\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20763\
        );

    \I__1892\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20760\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__20766\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__20763\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__20760\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3\
        );

    \I__1888\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20747\
        );

    \I__1887\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20744\
        );

    \I__1886\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20739\
        );

    \I__1885\ : InMux
    port map (
            O => \N__20750\,
            I => \N__20739\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__20747\,
            I => \spi_master_inst.sclk_gen_u0.N_1531\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__20744\,
            I => \spi_master_inst.sclk_gen_u0.N_1531\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__20739\,
            I => \spi_master_inst.sclk_gen_u0.N_1531\
        );

    \I__1881\ : InMux
    port map (
            O => \N__20732\,
            I => \N__20728\
        );

    \I__1880\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20725\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__20728\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_start_iZ0\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__20725\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_start_iZ0\
        );

    \I__1877\ : InMux
    port map (
            O => \N__20720\,
            I => \N__20711\
        );

    \I__1876\ : InMux
    port map (
            O => \N__20719\,
            I => \N__20711\
        );

    \I__1875\ : InMux
    port map (
            O => \N__20718\,
            I => \N__20711\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__20711\,
            I => \N__20703\
        );

    \I__1873\ : InMux
    port map (
            O => \N__20710\,
            I => \N__20692\
        );

    \I__1872\ : InMux
    port map (
            O => \N__20709\,
            I => \N__20692\
        );

    \I__1871\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20692\
        );

    \I__1870\ : InMux
    port map (
            O => \N__20707\,
            I => \N__20692\
        );

    \I__1869\ : InMux
    port map (
            O => \N__20706\,
            I => \N__20692\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__20703\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_start_i_i\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__20692\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_start_i_i\
        );

    \I__1866\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20682\
        );

    \I__1865\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20677\
        );

    \I__1864\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20677\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__20682\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__20677\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0\
        );

    \I__1861\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20667\
        );

    \I__1860\ : InMux
    port map (
            O => \N__20671\,
            I => \N__20664\
        );

    \I__1859\ : InMux
    port map (
            O => \N__20670\,
            I => \N__20661\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__20667\,
            I => \N__20658\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__20664\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__20661\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__20658\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__20651\,
            I => \N__20646\
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__20650\,
            I => \N__20643\
        );

    \I__1852\ : InMux
    port map (
            O => \N__20649\,
            I => \N__20640\
        );

    \I__1851\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20637\
        );

    \I__1850\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20634\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__20640\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__20637\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__20634\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3\
        );

    \I__1846\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20622\
        );

    \I__1845\ : InMux
    port map (
            O => \N__20626\,
            I => \N__20619\
        );

    \I__1844\ : InMux
    port map (
            O => \N__20625\,
            I => \N__20616\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__20622\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__20619\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__20616\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__20609\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__20606\,
            I => \spi_master_inst.sclk_gen_u0.N_48_cascade_\
        );

    \I__1838\ : InMux
    port map (
            O => \N__20603\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6\
        );

    \I__1837\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20597\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__20597\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_s_1\
        );

    \I__1835\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20590\
        );

    \I__1834\ : InMux
    port map (
            O => \N__20593\,
            I => \N__20587\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__20590\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__20587\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__20582\,
            I => \N__20579\
        );

    \I__1830\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20572\
        );

    \I__1829\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20572\
        );

    \I__1828\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20568\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__20572\,
            I => \N__20565\
        );

    \I__1826\ : InMux
    port map (
            O => \N__20571\,
            I => \N__20562\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__20568\,
            I => \N__20559\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__20565\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__20562\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0\
        );

    \I__1822\ : Odrv12
    port map (
            O => \N__20559\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0\
        );

    \I__1821\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__20549\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_s_0\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__20546\,
            I => \N__20542\
        );

    \I__1818\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20533\
        );

    \I__1817\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20530\
        );

    \I__1816\ : InMux
    port map (
            O => \N__20541\,
            I => \N__20523\
        );

    \I__1815\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20523\
        );

    \I__1814\ : InMux
    port map (
            O => \N__20539\,
            I => \N__20523\
        );

    \I__1813\ : InMux
    port map (
            O => \N__20538\,
            I => \N__20516\
        );

    \I__1812\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20516\
        );

    \I__1811\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20516\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__20533\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__20530\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__20523\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__20516\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i\
        );

    \I__1806\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20500\
        );

    \I__1805\ : InMux
    port map (
            O => \N__20506\,
            I => \N__20500\
        );

    \I__1804\ : InMux
    port map (
            O => \N__20505\,
            I => \N__20497\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__20500\,
            I => \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__20497\,
            I => \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i\
        );

    \I__1801\ : InMux
    port map (
            O => \N__20492\,
            I => \N__20489\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__20489\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0\
        );

    \I__1799\ : InMux
    port map (
            O => \N__20486\,
            I => \bfn_3_8_0_\
        );

    \I__1798\ : InMux
    port map (
            O => \N__20483\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_0\
        );

    \I__1797\ : InMux
    port map (
            O => \N__20480\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_1\
        );

    \I__1796\ : InMux
    port map (
            O => \N__20477\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_2\
        );

    \I__1795\ : InMux
    port map (
            O => \N__20474\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_3\
        );

    \I__1794\ : IoInMux
    port map (
            O => \N__20471\,
            I => \N__20468\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__20468\,
            I => \N__20465\
        );

    \I__1792\ : Span4Mux_s3_v
    port map (
            O => \N__20465\,
            I => \N__20462\
        );

    \I__1791\ : Span4Mux_h
    port map (
            O => \N__20462\,
            I => \N__20459\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__20459\,
            I => \DAC_cs_c\
        );

    \I__1789\ : InMux
    port map (
            O => \N__20456\,
            I => \bfn_3_6_0_\
        );

    \I__1788\ : InMux
    port map (
            O => \N__20453\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0\
        );

    \I__1787\ : InMux
    port map (
            O => \N__20450\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1\
        );

    \I__1786\ : InMux
    port map (
            O => \N__20447\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2\
        );

    \I__1785\ : InMux
    port map (
            O => \N__20444\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3\
        );

    \I__1784\ : InMux
    port map (
            O => \N__20441\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4\
        );

    \I__1783\ : InMux
    port map (
            O => \N__20438\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__20435\,
            I => \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1_cascade_\
        );

    \I__1781\ : CascadeMux
    port map (
            O => \N__20432\,
            I => \spi_master_inst.sclk_gen_u0.N_1531_cascade_\
        );

    \I__1780\ : CascadeMux
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__1779\ : InMux
    port map (
            O => \N__20426\,
            I => \N__20417\
        );

    \I__1778\ : InMux
    port map (
            O => \N__20425\,
            I => \N__20417\
        );

    \I__1777\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20417\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__20417\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1\
        );

    \I__1775\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__1773\ : Span12Mux_h
    port map (
            O => \N__20408\,
            I => \N__20405\
        );

    \I__1772\ : Span12Mux_v
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__1771\ : Odrv12
    port map (
            O => \N__20402\,
            I => button_mode_c
        );

    \I__1770\ : IoInMux
    port map (
            O => \N__20399\,
            I => \N__20396\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__1768\ : Odrv12
    port map (
            O => \N__20393\,
            I => \button_mode_ibuf_RNIN5KZ0Z7\
        );

    \I__1767\ : InMux
    port map (
            O => \N__20390\,
            I => \sRAM_pointer_write_cry_10\
        );

    \I__1766\ : InMux
    port map (
            O => \N__20387\,
            I => \sRAM_pointer_write_cry_11\
        );

    \I__1765\ : InMux
    port map (
            O => \N__20384\,
            I => \sRAM_pointer_write_cry_12\
        );

    \I__1764\ : InMux
    port map (
            O => \N__20381\,
            I => \sRAM_pointer_write_cry_13\
        );

    \I__1763\ : InMux
    port map (
            O => \N__20378\,
            I => \sRAM_pointer_write_cry_14\
        );

    \I__1762\ : InMux
    port map (
            O => \N__20375\,
            I => \bfn_1_13_0_\
        );

    \I__1761\ : InMux
    port map (
            O => \N__20372\,
            I => \sRAM_pointer_write_cry_16\
        );

    \I__1760\ : InMux
    port map (
            O => \N__20369\,
            I => \sRAM_pointer_write_cry_17\
        );

    \I__1759\ : CEMux
    port map (
            O => \N__20366\,
            I => \N__20357\
        );

    \I__1758\ : CEMux
    port map (
            O => \N__20365\,
            I => \N__20357\
        );

    \I__1757\ : CEMux
    port map (
            O => \N__20364\,
            I => \N__20357\
        );

    \I__1756\ : GlobalMux
    port map (
            O => \N__20357\,
            I => \N__20354\
        );

    \I__1755\ : gio2CtrlBuf
    port map (
            O => \N__20354\,
            I => \N_1487_g\
        );

    \I__1754\ : InMux
    port map (
            O => \N__20351\,
            I => \sRAM_pointer_write_cry_1\
        );

    \I__1753\ : InMux
    port map (
            O => \N__20348\,
            I => \sRAM_pointer_write_cry_2\
        );

    \I__1752\ : InMux
    port map (
            O => \N__20345\,
            I => \sRAM_pointer_write_cry_3\
        );

    \I__1751\ : InMux
    port map (
            O => \N__20342\,
            I => \sRAM_pointer_write_cry_4\
        );

    \I__1750\ : InMux
    port map (
            O => \N__20339\,
            I => \sRAM_pointer_write_cry_5\
        );

    \I__1749\ : InMux
    port map (
            O => \N__20336\,
            I => \sRAM_pointer_write_cry_6\
        );

    \I__1748\ : InMux
    port map (
            O => \N__20333\,
            I => \bfn_1_12_0_\
        );

    \I__1747\ : InMux
    port map (
            O => \N__20330\,
            I => \sRAM_pointer_write_cry_8\
        );

    \I__1746\ : InMux
    port map (
            O => \N__20327\,
            I => \sRAM_pointer_write_cry_9\
        );

    \I__1745\ : InMux
    port map (
            O => \N__20324\,
            I => \bfn_1_11_0_\
        );

    \I__1744\ : InMux
    port map (
            O => \N__20321\,
            I => \sRAM_pointer_write_cry_0\
        );

    \I__1743\ : IoInMux
    port map (
            O => \N__20318\,
            I => \N__20315\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__20315\,
            I => \N__20312\
        );

    \I__1741\ : Span4Mux_s0_h
    port map (
            O => \N__20312\,
            I => \N__20309\
        );

    \I__1740\ : Span4Mux_h
    port map (
            O => \N__20309\,
            I => \N__20306\
        );

    \I__1739\ : Sp12to4
    port map (
            O => \N__20306\,
            I => \N__20303\
        );

    \I__1738\ : Span12Mux_v
    port map (
            O => \N__20303\,
            I => \N__20300\
        );

    \I__1737\ : Span12Mux_h
    port map (
            O => \N__20300\,
            I => \N__20297\
        );

    \I__1736\ : Odrv12
    port map (
            O => \N__20297\,
            I => \pll128M2_inst.pll_clk128\
        );

    \I__1735\ : IoInMux
    port map (
            O => \N__20294\,
            I => \N__20291\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__20291\,
            I => \N__20288\
        );

    \I__1733\ : Span4Mux_s2_h
    port map (
            O => \N__20288\,
            I => \N__20285\
        );

    \I__1732\ : Span4Mux_v
    port map (
            O => \N__20285\,
            I => \N__20282\
        );

    \I__1731\ : Sp12to4
    port map (
            O => \N__20282\,
            I => \N__20279\
        );

    \I__1730\ : Span12Mux_s11_h
    port map (
            O => \N__20279\,
            I => \N__20276\
        );

    \I__1729\ : Span12Mux_h
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__1728\ : Odrv12
    port map (
            O => \N__20273\,
            I => cs_rpi2flash_c
        );

    \I__1727\ : IoInMux
    port map (
            O => \N__20270\,
            I => \N__20267\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__20267\,
            I => \N__20264\
        );

    \I__1725\ : Span4Mux_s3_v
    port map (
            O => \N__20264\,
            I => \N__20261\
        );

    \I__1724\ : Sp12to4
    port map (
            O => \N__20261\,
            I => \N__20258\
        );

    \I__1723\ : Span12Mux_h
    port map (
            O => \N__20258\,
            I => \N__20255\
        );

    \I__1722\ : Span12Mux_v
    port map (
            O => \N__20255\,
            I => \N__20252\
        );

    \I__1721\ : Odrv12
    port map (
            O => \N__20252\,
            I => clk_c
        );

    \I__1720\ : IoInMux
    port map (
            O => \N__20249\,
            I => \N__20246\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__20246\,
            I => \N__20243\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__20243\,
            I => \pll128M2_inst.pll_clk64_0\
        );

    \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C\ : INV
    port map (
            O => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            I => \N__48262\
        );

    \INVspi_slave_inst.rx_done_neg_sclk_iC\ : INV
    port map (
            O => \INVspi_slave_inst.rx_done_neg_sclk_iC_net\,
            I => \N__48265\
        );

    \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C\ : INV
    port map (
            O => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            I => \N__48261\
        );

    \IN_MUX_bfv_6_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_12_0_\
        );

    \IN_MUX_bfv_6_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un8_trig_prev_0_cry_7,
            carryinitout => \bfn_6_13_0_\
        );

    \IN_MUX_bfv_20_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_10_0_\
        );

    \IN_MUX_bfv_20_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_scounterdac_cry_8,
            carryinitout => \bfn_20_11_0_\
        );

    \IN_MUX_bfv_13_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_14_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_sacqtime_cry_7,
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_sacqtime_cry_15,
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_sacqtime_cry_23,
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_16_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_13_0_\
        );

    \IN_MUX_bfv_16_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_button_debounce_counter_cry_8,
            carryinitout => \bfn_16_14_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_button_debounce_counter_cry_16,
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO\,
            carryinitout => \bfn_6_8_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un7_spon_cry_7,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un7_spon_cry_15,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un7_spon_cry_23,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_sdacdyn_cry_7,
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_sdacdyn_cry_15,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_sdacdyn_cry_23,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_spoff_cry_7,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_spoff_cry_15,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_spoff_cry_23,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_speriod_cry_7,
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_speriod_cry_15,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_speriod_cry_23,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_sacqtime_cry_7,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_sacqtime_cry_15,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_sacqtime_cry_23,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_spoff_cry_7,
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_spoff_cry_15,
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_spoff_cry_23,
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un10_trig_prev_cry_7,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un10_trig_prev_cry_15,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_22_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_7_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_3_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_6_0_\
        );

    \IN_MUX_bfv_3_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_8_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_sTrigCounter_cry_7\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sRAM_pointer_write_cry_7\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sRAM_pointer_write_cry_15\,
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sRAM_pointer_read_cry_7\,
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sRAM_pointer_read_cry_15\,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sCounter_cry_7\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sCounter_cry_15\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_15_0_\
        );

    \reset_rpi_ibuf_RNIIUT3_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__24725\,
            GLOBALBUFFEROUTPUT => \LED3_c_i_g\
        );

    \un4_sacqtime_cry_23_c_RNI2CQM_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__26744\,
            GLOBALBUFFEROUTPUT => \N_1487_g\
        );

    \pll128M2_inst.PLLOUTCOREB_derived_clock_RNI5L14\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__20249\,
            GLOBALBUFFEROUTPUT => pll_clk64_0_g
        );

    \spi_sclk_inferred_clock_RNIH8F3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__25799\,
            GLOBALBUFFEROUTPUT => spi_sclk_g
        );

    \sSPI_MSB0LSB1_RNILL2C1_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__39191\,
            GLOBALBUFFEROUTPUT => \N_28_g\
        );

    \sCounterDAC_RNIBR1C_0_5\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__48179\,
            GLOBALBUFFEROUTPUT => op_eq_scounterdac10_g
        );

    \pll128M2_inst.PLLOUTCOREA_derived_clock_RNI4765\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__20318\,
            GLOBALBUFFEROUTPUT => pll_clk128_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \button_mode_ibuf_RNIN5K7_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__20399\,
            GLOBALBUFFEROUTPUT => \N_3154_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \sRAM_pointer_write_0_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39407\,
            in1 => \N__35872\,
            in2 => \_gnd_net_\,
            in3 => \N__20324\,
            lcout => \sRAM_pointer_writeZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \sRAM_pointer_write_cry_0\,
            clk => \N__52346\,
            ce => \N__20364\,
            sr => \N__51801\
        );

    \sRAM_pointer_write_1_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39399\,
            in1 => \N__36058\,
            in2 => \_gnd_net_\,
            in3 => \N__20321\,
            lcout => \sRAM_pointer_writeZ0Z_1\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_0\,
            carryout => \sRAM_pointer_write_cry_1\,
            clk => \N__52346\,
            ce => \N__20364\,
            sr => \N__51801\
        );

    \sRAM_pointer_write_2_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39408\,
            in1 => \N__36100\,
            in2 => \_gnd_net_\,
            in3 => \N__20351\,
            lcout => \sRAM_pointer_writeZ0Z_2\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_1\,
            carryout => \sRAM_pointer_write_cry_2\,
            clk => \N__52346\,
            ce => \N__20364\,
            sr => \N__51801\
        );

    \sRAM_pointer_write_3_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39400\,
            in1 => \N__43510\,
            in2 => \_gnd_net_\,
            in3 => \N__20348\,
            lcout => \sRAM_pointer_writeZ0Z_3\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_2\,
            carryout => \sRAM_pointer_write_cry_3\,
            clk => \N__52346\,
            ce => \N__20364\,
            sr => \N__51801\
        );

    \sRAM_pointer_write_4_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39409\,
            in1 => \N__43573\,
            in2 => \_gnd_net_\,
            in3 => \N__20345\,
            lcout => \sRAM_pointer_writeZ0Z_4\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_3\,
            carryout => \sRAM_pointer_write_cry_4\,
            clk => \N__52346\,
            ce => \N__20364\,
            sr => \N__51801\
        );

    \sRAM_pointer_write_5_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39401\,
            in1 => \N__35227\,
            in2 => \_gnd_net_\,
            in3 => \N__20342\,
            lcout => \sRAM_pointer_writeZ0Z_5\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_4\,
            carryout => \sRAM_pointer_write_cry_5\,
            clk => \N__52346\,
            ce => \N__20364\,
            sr => \N__51801\
        );

    \sRAM_pointer_write_6_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39410\,
            in1 => \N__36001\,
            in2 => \_gnd_net_\,
            in3 => \N__20339\,
            lcout => \sRAM_pointer_writeZ0Z_6\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_5\,
            carryout => \sRAM_pointer_write_cry_6\,
            clk => \N__52346\,
            ce => \N__20364\,
            sr => \N__51801\
        );

    \sRAM_pointer_write_7_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39402\,
            in1 => \N__36181\,
            in2 => \_gnd_net_\,
            in3 => \N__20336\,
            lcout => \sRAM_pointer_writeZ0Z_7\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_6\,
            carryout => \sRAM_pointer_write_cry_7\,
            clk => \N__52346\,
            ce => \N__20364\,
            sr => \N__51801\
        );

    \sRAM_pointer_write_8_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39406\,
            in1 => \N__43645\,
            in2 => \_gnd_net_\,
            in3 => \N__20333\,
            lcout => \sRAM_pointer_writeZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \sRAM_pointer_write_cry_8\,
            clk => \N__52348\,
            ce => \N__20365\,
            sr => \N__51788\
        );

    \sRAM_pointer_write_9_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39359\,
            in1 => \N__36250\,
            in2 => \_gnd_net_\,
            in3 => \N__20330\,
            lcout => \sRAM_pointer_writeZ0Z_9\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_8\,
            carryout => \sRAM_pointer_write_cry_9\,
            clk => \N__52348\,
            ce => \N__20365\,
            sr => \N__51788\
        );

    \sRAM_pointer_write_10_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39403\,
            in1 => \N__35809\,
            in2 => \_gnd_net_\,
            in3 => \N__20327\,
            lcout => \sRAM_pointer_writeZ0Z_10\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_9\,
            carryout => \sRAM_pointer_write_cry_10\,
            clk => \N__52348\,
            ce => \N__20365\,
            sr => \N__51788\
        );

    \sRAM_pointer_write_11_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39356\,
            in1 => \N__35737\,
            in2 => \_gnd_net_\,
            in3 => \N__20390\,
            lcout => \sRAM_pointer_writeZ0Z_11\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_10\,
            carryout => \sRAM_pointer_write_cry_11\,
            clk => \N__52348\,
            ce => \N__20365\,
            sr => \N__51788\
        );

    \sRAM_pointer_write_12_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39404\,
            in1 => \N__35689\,
            in2 => \_gnd_net_\,
            in3 => \N__20387\,
            lcout => \sRAM_pointer_writeZ0Z_12\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_11\,
            carryout => \sRAM_pointer_write_cry_12\,
            clk => \N__52348\,
            ce => \N__20365\,
            sr => \N__51788\
        );

    \sRAM_pointer_write_13_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39357\,
            in1 => \N__35605\,
            in2 => \_gnd_net_\,
            in3 => \N__20384\,
            lcout => \sRAM_pointer_writeZ0Z_13\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_12\,
            carryout => \sRAM_pointer_write_cry_13\,
            clk => \N__52348\,
            ce => \N__20365\,
            sr => \N__51788\
        );

    \sRAM_pointer_write_14_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39405\,
            in1 => \N__35560\,
            in2 => \_gnd_net_\,
            in3 => \N__20381\,
            lcout => \sRAM_pointer_writeZ0Z_14\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_13\,
            carryout => \sRAM_pointer_write_cry_14\,
            clk => \N__52348\,
            ce => \N__20365\,
            sr => \N__51788\
        );

    \sRAM_pointer_write_15_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39358\,
            in1 => \N__35464\,
            in2 => \_gnd_net_\,
            in3 => \N__20378\,
            lcout => \sRAM_pointer_writeZ0Z_15\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_14\,
            carryout => \sRAM_pointer_write_cry_15\,
            clk => \N__52348\,
            ce => \N__20365\,
            sr => \N__51788\
        );

    \sRAM_pointer_write_16_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39397\,
            in1 => \N__35395\,
            in2 => \_gnd_net_\,
            in3 => \N__20375\,
            lcout => \sRAM_pointer_writeZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \sRAM_pointer_write_cry_16\,
            clk => \N__52349\,
            ce => \N__20366\,
            sr => \N__51776\
        );

    \sRAM_pointer_write_17_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39396\,
            in1 => \N__36388\,
            in2 => \_gnd_net_\,
            in3 => \N__20372\,
            lcout => \sRAM_pointer_writeZ0Z_17\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_16\,
            carryout => \sRAM_pointer_write_cry_17\,
            clk => \N__52349\,
            ce => \N__20366\,
            sr => \N__51776\
        );

    \sRAM_pointer_write_18_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39398\,
            in1 => \N__36322\,
            in2 => \_gnd_net_\,
            in3 => \N__20369\,
            lcout => \sRAM_pointer_writeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52349\,
            ce => \N__20366\,
            sr => \N__51776\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_start_i_RNIPPNJ2_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20577\,
            in2 => \_gnd_net_\,
            in3 => \N__20505\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIIUTC1_7_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20904\,
            in1 => \N__21006\,
            in2 => \N__20935\,
            in3 => \N__20961\,
            lcout => OPEN,
            ltout => \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIL2KE2_1_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__21027\,
            in1 => \N__20982\,
            in2 => \N__20435\,
            in3 => \N__20593\,
            lcout => \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4D3E3_1_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20672\,
            in1 => \N__20777\,
            in2 => \N__20650\,
            in3 => \N__21139\,
            lcout => \spi_master_inst.sclk_gen_u0.N_1531\,
            ltout => \spi_master_inst.sclk_gen_u0.N_1531_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0RFT3_1_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20769\,
            in2 => \N__20432\,
            in3 => \N__20424\,
            lcout => \spi_master_inst.sclk_gen_u0.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_1_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__20751\,
            in1 => \N__24378\,
            in2 => \N__20429\,
            in3 => \N__24551\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48488\,
            ce => 'H',
            sr => \N__51818\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI1JPL3_1_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20425\,
            in2 => \_gnd_net_\,
            in3 => \N__20750\,
            lcout => \spi_master_inst.sclk_gen_u0.N_1540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_start_i_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000011101111"
        )
    port map (
            in0 => \N__20732\,
            in1 => \N__24550\,
            in2 => \N__24387\,
            in3 => \N__20849\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_start_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48489\,
            ce => 'H',
            sr => \N__51810\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_3_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110010100000"
        )
    port map (
            in0 => \N__24460\,
            in1 => \N__20753\,
            in2 => \N__24513\,
            in3 => \N__20771\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48489\,
            ce => 'H',
            sr => \N__51810\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_start_i_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__20571\,
            in1 => \N__20842\,
            in2 => \N__24512\,
            in3 => \N__20861\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48489\,
            ce => 'H',
            sr => \N__51810\
        );

    \button_mode_ibuf_RNIN5K7_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__20414\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49445\,
            lcout => \button_mode_ibuf_RNIN5KZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_12_7_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50027\,
            lcout => \sDAC_mem_12Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52341\,
            ce => \N__36959\,
            sr => \N__51789\
        );

    \spi_master_inst.o_slave_csn_0_LC_3_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21077\,
            lcout => \DAC_cs_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48464\,
            ce => 'H',
            sr => \N__51827\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_0_LC_3_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20492\,
            in2 => \_gnd_net_\,
            in3 => \N__20456\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_i_s_0\,
            ltout => OPEN,
            carryin => \bfn_3_6_0_\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_1_LC_3_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20594\,
            in2 => \_gnd_net_\,
            in3 => \N__20453\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_i_s_1\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_2_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20536\,
            in1 => \N__21028\,
            in2 => \_gnd_net_\,
            in3 => \N__20450\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2\,
            clk => \N__48478\,
            ce => 'H',
            sr => \N__51822\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_3_LC_3_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20539\,
            in1 => \N__20983\,
            in2 => \_gnd_net_\,
            in3 => \N__20447\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3\,
            clk => \N__48478\,
            ce => 'H',
            sr => \N__51822\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_4_LC_3_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20537\,
            in1 => \N__20965\,
            in2 => \_gnd_net_\,
            in3 => \N__20444\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4\,
            clk => \N__48478\,
            ce => 'H',
            sr => \N__51822\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_5_LC_3_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20540\,
            in1 => \N__21010\,
            in2 => \_gnd_net_\,
            in3 => \N__20441\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5\,
            clk => \N__48478\,
            ce => 'H',
            sr => \N__51822\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_6_LC_3_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20538\,
            in1 => \N__20905\,
            in2 => \_gnd_net_\,
            in3 => \N__20438\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6\,
            clk => \N__48478\,
            ce => 'H',
            sr => \N__51822\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_7_LC_3_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20541\,
            in1 => \N__20931\,
            in2 => \_gnd_net_\,
            in3 => \N__20603\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48478\,
            ce => 'H',
            sr => \N__51822\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_1_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111110101010"
        )
    port map (
            in0 => \N__20600\,
            in1 => \N__20507\,
            in2 => \N__20582\,
            in3 => \N__20545\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48482\,
            ce => 'H',
            sr => \N__51819\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_0_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__20578\,
            in1 => \N__20552\,
            in2 => \N__20546\,
            in3 => \N__20506\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48482\,
            ce => 'H',
            sr => \N__51819\
        );

    \spi_master_inst.sclk_gen_u0.falling_count_start_i_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__27943\,
            in1 => \N__24332\,
            in2 => \_gnd_net_\,
            in3 => \N__20843\,
            lcout => \spi_master_inst.sclk_gen_u0.falling_count_start_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48482\,
            ce => 'H',
            sr => \N__51819\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_0_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101111101110"
        )
    port map (
            in0 => \N__20706\,
            in1 => \N__20687\,
            in2 => \_gnd_net_\,
            in3 => \N__20486\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_3_8_0_\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_0\,
            clk => \N__48485\,
            ce => 'H',
            sr => \N__51811\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_1_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20718\,
            in1 => \N__20671\,
            in2 => \_gnd_net_\,
            in3 => \N__20483\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_0\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_1\,
            clk => \N__48485\,
            ce => 'H',
            sr => \N__51811\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_2_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20707\,
            in1 => \N__20627\,
            in2 => \_gnd_net_\,
            in3 => \N__20480\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_1\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_2\,
            clk => \N__48485\,
            ce => 'H',
            sr => \N__51811\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_3_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20719\,
            in1 => \N__20649\,
            in2 => \_gnd_net_\,
            in3 => \N__20477\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_2\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_3\,
            clk => \N__48485\,
            ce => 'H',
            sr => \N__51811\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_4_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20708\,
            in1 => \N__21157\,
            in2 => \_gnd_net_\,
            in3 => \N__20474\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_3\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_4\,
            clk => \N__48485\,
            ce => 'H',
            sr => \N__51811\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_5_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20720\,
            in1 => \N__21190\,
            in2 => \_gnd_net_\,
            in3 => \N__20786\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_4\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_5\,
            clk => \N__48485\,
            ce => 'H',
            sr => \N__51811\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_6_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20709\,
            in1 => \N__21206\,
            in2 => \_gnd_net_\,
            in3 => \N__20783\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_5\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_6\,
            clk => \N__48485\,
            ce => 'H',
            sr => \N__51811\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_7_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21172\,
            in1 => \N__20710\,
            in2 => \_gnd_net_\,
            in3 => \N__20780\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48485\,
            ce => 'H',
            sr => \N__51811\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4MGR_0_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20625\,
            in2 => \_gnd_net_\,
            in3 => \N__20685\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI3LPL3_3_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20770\,
            in2 => \_gnd_net_\,
            in3 => \N__20752\,
            lcout => \spi_master_inst.sclk_gen_u0.N_150_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNI6TQC_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20731\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_start_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_RNIAE1N1_0_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__20686\,
            in1 => \N__20670\,
            in2 => \N__20651\,
            in3 => \N__20626\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4\,
            ltout => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0IPL3_0_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21107\,
            in2 => \N__20609\,
            in3 => \N__21143\,
            lcout => \spi_master_inst.sclk_gen_u0.N_48\,
            ltout => \spi_master_inst.sclk_gen_u0.N_48_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNO_0_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__24495\,
            in1 => \N__24459\,
            in2 => \N__20606\,
            in3 => \N__20860\,
            lcout => \spi_master_inst.sclk_gen_u0.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_2_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__24385\,
            in1 => \N__24543\,
            in2 => \_gnd_net_\,
            in3 => \N__20838\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48490\,
            ce => 'H',
            sr => \N__51790\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_4_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__24499\,
            in1 => \N__24461\,
            in2 => \_gnd_net_\,
            in3 => \N__20822\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48490\,
            ce => 'H',
            sr => \N__51790\
        );

    \sAddress_7_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__26198\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49929\,
            lcout => \sAddressZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52332\,
            ce => \N__23423\,
            sr => \N__51777\
        );

    \sAddress_6_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50327\,
            in2 => \_gnd_net_\,
            in3 => \N__26197\,
            lcout => \sAddressZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52332\,
            ce => \N__23423\,
            sr => \N__51777\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI73G42_2_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21421\,
            in1 => \N__21236\,
            in2 => \_gnd_net_\,
            in3 => \N__20792\,
            lcout => OPEN,
            ltout => \spi_master_inst.spi_data_path_u1.N_1414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI60IB4_1_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__21512\,
            in1 => \_gnd_net_\,
            in2 => \N__20816\,
            in3 => \N__21242\,
            lcout => OPEN,
            ltout => \spi_master_inst.spi_data_path_u1.N_1415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI70MD9_0_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__21578\,
            in1 => \N__21038\,
            in2 => \N__20813\,
            in3 => \N__21076\,
            lcout => \DAC_mosi_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01_1_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25748\,
            in1 => \N__21797\,
            in2 => \_gnd_net_\,
            in3 => \N__24668\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01_0_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47567\,
            in1 => \N__21767\,
            in2 => \_gnd_net_\,
            in3 => \N__24667\,
            lcout => OPEN,
            ltout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI3VF42_2_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23228\,
            in2 => \N__21044\,
            in3 => \N__21416\,
            lcout => OPEN,
            ltout => \spi_master_inst.spi_data_path_u1.N_1421_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIUNHB4_1_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__21224\,
            in1 => \_gnd_net_\,
            in2 => \N__21041\,
            in3 => \N__21511\,
            lcout => \spi_master_inst.spi_data_path_u1.N_1422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.o_sclk_RNIH6AC_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__27989\,
            in1 => \N__24386\,
            in2 => \_gnd_net_\,
            in3 => \N__20875\,
            lcout => \spi_master_inst.o_sclk_RNIH6AC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.div_clk_i_RNO_0_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21032\,
            in1 => \N__21011\,
            in2 => \N__20990\,
            in3 => \N__20966\,
            lcout => \spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.div_clk_i_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__20945\,
            in1 => \N__20939\,
            in2 => \_gnd_net_\,
            in3 => \N__20912\,
            lcout => \spi_master_inst.sclk_gen_u0.div_clk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48474\,
            ce => 'H',
            sr => \N__51802\
        );

    \spi_master_inst.sclk_gen_u0.o_sclk_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27993\,
            in2 => \_gnd_net_\,
            in3 => \N__24389\,
            lcout => \DAC_sclk_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48474\,
            ce => 'H',
            sr => \N__51802\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_2_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001101000101010"
        )
    port map (
            in0 => \N__21401\,
            in1 => \N__21331\,
            in2 => \N__21296\,
            in3 => \N__21365\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48474\,
            ce => 'H',
            sr => \N__51802\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIL1LO1_2_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21476\,
            in1 => \N__21400\,
            in2 => \_gnd_net_\,
            in3 => \N__24651\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6\,
            ltout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_i_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101011100010"
        )
    port map (
            in0 => \N__23170\,
            in1 => \N__21284\,
            in2 => \N__20864\,
            in3 => \N__21066\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48474\,
            ce => 'H',
            sr => \N__51802\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_3_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100011001001100"
        )
    port map (
            in0 => \N__21283\,
            in1 => \N__24652\,
            in2 => \N__21332\,
            in3 => \N__21356\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48474\,
            ce => 'H',
            sr => \N__51802\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_RNIQU1N1_7_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21205\,
            in1 => \N__21191\,
            in2 => \N__21176\,
            in3 => \N__21158\,
            lcout => \spi_master_inst.sclk_gen_u0.N_1737\,
            ltout => \spi_master_inst.sclk_gen_u0.N_1737_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_0_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__21089\,
            in1 => \N__21122\,
            in2 => \N__21110\,
            in3 => \N__21103\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48479\,
            ce => 'H',
            sr => \N__51791\
        );

    \spi_master_inst.sclk_gen_u0.o_ss_start_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100111010"
        )
    port map (
            in0 => \N__21065\,
            in1 => \N__24454\,
            in2 => \N__24521\,
            in3 => \N__21088\,
            lcout => \spi_master_inst.ss_start_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48479\,
            ce => 'H',
            sr => \N__51791\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52_2_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__24649\,
            in1 => \N__21064\,
            in2 => \N__21415\,
            in3 => \N__21475\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_mosi_ready64_prev_e_0_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22001\,
            lcout => \spi_mosi_ready64_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52340\,
            ce => \N__49426\,
            sr => \_gnd_net_\
        );

    \spi_mosi_ready64_prev2_e_0_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21446\,
            lcout => \spi_mosi_ready64_prevZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52331\,
            ce => \N__49441\,
            sr => \_gnd_net_\
        );

    \spi_mosi_ready64_prev3_e_0_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21458\,
            lcout => \spi_mosi_ready64_prevZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52331\,
            ce => \N__49441\,
            sr => \_gnd_net_\
        );

    \sSingleCont_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26399\,
            in2 => \_gnd_net_\,
            in3 => \N__22526\,
            lcout => \LED_MODE_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48491\,
            ce => 'H',
            sr => \N__51736\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIMGLT1_2_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21803\,
            in1 => \N__24614\,
            in2 => \_gnd_net_\,
            in3 => \N__21422\,
            lcout => \spi_master_inst.spi_data_path_u1.N_1411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4Q_14_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21218\,
            in1 => \N__21773\,
            in2 => \_gnd_net_\,
            in3 => \N__24693\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4Q_13_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24682\,
            in1 => \N__21785\,
            in2 => \_gnd_net_\,
            in3 => \N__21779\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIICLT1_2_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21417\,
            in1 => \N__21230\,
            in2 => \_gnd_net_\,
            in3 => \N__23219\,
            lcout => \spi_master_inst.spi_data_path_u1.N_1418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_6_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21758\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48465\,
            ce => 'H',
            sr => \N__51803\
        );

    \spi_master_inst.sclk_gen_u0.delay_clk_i_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28000\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_clk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48465\,
            ce => 'H',
            sr => \N__51803\
        );

    \sDAC_mem_29_5_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44952\,
            lcout => \sDAC_mem_29Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52347\,
            ce => \N__23153\,
            sr => \N__51792\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_c_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21253\,
            in2 => \N__21577\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_LUT4_0_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21504\,
            in2 => \_gnd_net_\,
            in3 => \N__21209\,
            lcout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_LUT4_0_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21402\,
            in2 => \_gnd_net_\,
            in3 => \N__21359\,
            lcout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_LUT4_0_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24650\,
            in2 => \_gnd_net_\,
            in3 => \N__21350\,
            lcout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_4_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21282\,
            in1 => \N__21526\,
            in2 => \_gnd_net_\,
            in3 => \N__21347\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4\,
            clk => \N__48467\,
            ce => 'H',
            sr => \N__51778\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_0_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52738\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_1_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__52782\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_2_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52742\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_5_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21544\,
            in2 => \_gnd_net_\,
            in3 => \N__21344\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48471\,
            ce => \N__21297\,
            sr => \N__51763\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_1_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001111101000000"
        )
    port map (
            in0 => \N__21327\,
            in1 => \N__21341\,
            in2 => \N__21305\,
            in3 => \N__21503\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48475\,
            ce => 'H',
            sr => \N__51751\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_0_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001110001001100"
        )
    port map (
            in0 => \N__21326\,
            in1 => \N__21570\,
            in2 => \N__21304\,
            in3 => \N__21254\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48475\,
            ce => 'H',
            sr => \N__51751\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_RNI06S51_5_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__21563\,
            in1 => \N__21545\,
            in2 => \N__21530\,
            in3 => \N__21494\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_mosi_ready64_prev3_e_0_RNICM2C1_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21457\,
            in1 => \N__21445\,
            in2 => \N__21434\,
            in3 => \N__21991\,
            lcout => \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1\,
            ltout => \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sPointer_RNI85NC1_0_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21425\,
            in3 => \N__26098\,
            lcout => un1_spointer11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_mosi_ready_prev3_RNILKER_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21958\,
            in1 => \N__21970\,
            in2 => \N__21947\,
            in3 => \N__21992\,
            lcout => \spi_mosi_ready_prev3_RNILKERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_RNICMDR1_5_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22040\,
            in1 => \N__21844\,
            in2 => \N__21863\,
            in3 => \N__22012\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_i6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_0_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46324\,
            lcout => un8_trig_prev_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52302\,
            ce => \N__22682\,
            sr => \N__51724\
        );

    \sEETrigCounter_1_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50984\,
            lcout => \sEETrigCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52302\,
            ce => \N__22682\,
            sr => \N__51724\
        );

    \sEETrigCounter_2_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47413\,
            lcout => \sEETrigCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52302\,
            ce => \N__22682\,
            sr => \N__51724\
        );

    \sEETrigCounter_3_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46840\,
            lcout => \sEETrigCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52302\,
            ce => \N__22682\,
            sr => \N__51724\
        );

    \sEETrigCounter_4_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45554\,
            lcout => \sEETrigCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52302\,
            ce => \N__22682\,
            sr => \N__51724\
        );

    \sEETrigCounter_5_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45000\,
            lcout => \sEETrigCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52302\,
            ce => \N__22682\,
            sr => \N__51724\
        );

    \sEETrigCounter_6_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50328\,
            lcout => \sEETrigCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52302\,
            ce => \N__22682\,
            sr => \N__51724\
        );

    \sEETrigCounter_7_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50023\,
            lcout => \sEETrigCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52302\,
            ce => \N__22682\,
            sr => \N__51724\
        );

    \un8_trig_prev_0_cry_0_c_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22145\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_12_0_\,
            carryout => un8_trig_prev_0_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_trig_prev_0_cry_0_c_RNILB0M_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52763\,
            in2 => \N__21626\,
            in3 => \N__21617\,
            lcout => un10_trig_prev_1,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_0,
            carryout => un8_trig_prev_0_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_trig_prev_0_cry_1_c_RNINE1M_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52779\,
            in2 => \N__21614\,
            in3 => \N__21605\,
            lcout => un10_trig_prev_2,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_1,
            carryout => un8_trig_prev_0_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_trig_prev_0_cry_2_c_RNIPH2M_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52764\,
            in2 => \N__21602\,
            in3 => \N__21593\,
            lcout => un10_trig_prev_3,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_2,
            carryout => un8_trig_prev_0_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_trig_prev_0_cry_3_c_RNIRK3M_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52780\,
            in2 => \N__21590\,
            in3 => \N__21581\,
            lcout => un10_trig_prev_4,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_3,
            carryout => un8_trig_prev_0_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_trig_prev_0_cry_4_c_RNITN4M_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52765\,
            in2 => \N__21680\,
            in3 => \N__21671\,
            lcout => un10_trig_prev_5,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_4,
            carryout => un8_trig_prev_0_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_trig_prev_0_cry_5_c_RNIVQ5M_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52781\,
            in2 => \N__21668\,
            in3 => \N__21659\,
            lcout => un10_trig_prev_6,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_5,
            carryout => un8_trig_prev_0_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_trig_prev_0_cry_6_c_RNI1U6M_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52766\,
            in2 => \N__21656\,
            in3 => \N__21647\,
            lcout => un10_trig_prev_7,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_6,
            carryout => un8_trig_prev_0_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_trig_prev_0_cry_7_c_RNI318M_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52789\,
            in2 => \N__21689\,
            in3 => \N__21644\,
            lcout => un10_trig_prev_8,
            ltout => OPEN,
            carryin => \bfn_6_13_0_\,
            carryout => un8_trig_prev_0_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_trig_prev_0_cry_8_c_RNI549M_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52769\,
            in2 => \N__21812\,
            in3 => \N__21641\,
            lcout => un10_trig_prev_9,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_8,
            carryout => un8_trig_prev_0_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_trig_prev_0_cry_9_c_RNIEEGI_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52790\,
            in2 => \N__21740\,
            in3 => \N__21638\,
            lcout => un10_trig_prev_10,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_9,
            carryout => un8_trig_prev_0_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNINORL_11_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52767\,
            in2 => \N__21731\,
            in3 => \N__21635\,
            lcout => un10_trig_prev_11,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_10,
            carryout => un8_trig_prev_0_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIPRSL_12_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52787\,
            in2 => \N__21722\,
            in3 => \N__21632\,
            lcout => un10_trig_prev_12,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_11,
            carryout => un8_trig_prev_0_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIRUTL_13_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52768\,
            in2 => \N__21713\,
            in3 => \N__21629\,
            lcout => un10_trig_prev_13,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_12,
            carryout => un8_trig_prev_0_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIT1VL_14_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52788\,
            in2 => \N__21704\,
            in3 => \N__21746\,
            lcout => un10_trig_prev_14,
            ltout => OPEN,
            carryin => un8_trig_prev_0_cry_13,
            carryout => un8_trig_prev_0_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIV40M_15_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21695\,
            in2 => \_gnd_net_\,
            in3 => \N__21743\,
            lcout => un10_trig_prev_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_10_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47480\,
            lcout => \sEETrigCounterZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52333\,
            ce => \N__21932\,
            sr => \N__51695\
        );

    \sEETrigCounter_11_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46919\,
            lcout => \sEETrigCounterZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52333\,
            ce => \N__21932\,
            sr => \N__51695\
        );

    \sEETrigCounter_12_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45601\,
            lcout => \sEETrigCounterZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52333\,
            ce => \N__21932\,
            sr => \N__51695\
        );

    \sEETrigCounter_13_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45117\,
            lcout => \sEETrigCounterZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52333\,
            ce => \N__21932\,
            sr => \N__51695\
        );

    \sEETrigCounter_14_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50378\,
            lcout => \sEETrigCounterZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52333\,
            ce => \N__21932\,
            sr => \N__51695\
        );

    \sEETrigCounter_15_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50049\,
            lcout => \sEETrigCounterZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52333\,
            ce => \N__21932\,
            sr => \N__51695\
        );

    \sEETrigCounter_8_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46281\,
            lcout => \sEETrigCounterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52333\,
            ce => \N__21932\,
            sr => \N__51695\
        );

    \sEETrigCounter_9_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51068\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEETrigCounterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52333\,
            ce => \N__21932\,
            sr => \N__51695\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4Q_11_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25790\,
            in1 => \N__22316\,
            in2 => \_gnd_net_\,
            in3 => \N__24700\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_1_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23984\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48459\,
            ce => 'H',
            sr => \N__51804\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_5_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21752\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48459\,
            ce => 'H',
            sr => \N__51804\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_13_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24041\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48459\,
            ce => 'H',
            sr => \N__51804\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_14_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24032\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48459\,
            ce => 'H',
            sr => \N__51804\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_0_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23993\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48459\,
            ce => 'H',
            sr => \N__51804\
        );

    \spi_master_inst.spi_data_path_u1.data_in_6_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27170\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48461\,
            ce => \N__43902\,
            sr => \N__51793\
        );

    \spi_master_inst.spi_data_path_u1.data_in_5_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37127\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48461\,
            ce => \N__43902\,
            sr => \N__51793\
        );

    \sDAC_mem_35_0_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46130\,
            lcout => \sDAC_mem_35Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52342\,
            ce => \N__22544\,
            sr => \N__51779\
        );

    \sDAC_mem_35_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50717\,
            lcout => \sDAC_mem_35Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52342\,
            ce => \N__22544\,
            sr => \N__51779\
        );

    \sDAC_mem_35_2_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47120\,
            lcout => \sDAC_mem_35Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52342\,
            ce => \N__22544\,
            sr => \N__51779\
        );

    \sDAC_mem_35_3_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46520\,
            lcout => \sDAC_mem_35Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52342\,
            ce => \N__22544\,
            sr => \N__51779\
        );

    \sDAC_mem_35_4_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45225\,
            lcout => \sDAC_mem_35Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52342\,
            ce => \N__22544\,
            sr => \N__51779\
        );

    \sDAC_mem_35_5_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44732\,
            lcout => \sDAC_mem_35Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52342\,
            ce => \N__22544\,
            sr => \N__51779\
        );

    \sDAC_mem_35_6_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50169\,
            lcout => \sDAC_mem_35Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52342\,
            ce => \N__22544\,
            sr => \N__51779\
        );

    \sDAC_mem_35_7_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49671\,
            lcout => \sDAC_mem_35Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52342\,
            ce => \N__22544\,
            sr => \N__51779\
        );

    \sDAC_mem_22_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46042\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_22Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52334\,
            ce => \N__33883\,
            sr => \N__51764\
        );

    \sDAC_mem_22_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50903\,
            lcout => \sDAC_mem_22Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52334\,
            ce => \N__33883\,
            sr => \N__51764\
        );

    \sDAC_mem_22_2_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47202\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_22Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52334\,
            ce => \N__33883\,
            sr => \N__51764\
        );

    \sDAC_mem_22_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46604\,
            lcout => \sDAC_mem_22Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52334\,
            ce => \N__33883\,
            sr => \N__51764\
        );

    \sDAC_mem_22_7_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49726\,
            lcout => \sDAC_mem_22Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52334\,
            ce => \N__33883\,
            sr => \N__51764\
        );

    \sAddress_RNIQ63A_6_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__21880\,
            in1 => \N__40861\,
            in2 => \N__21917\,
            in3 => \N__22609\,
            lcout => \N_316\,
            ltout => \N_316_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIUTJC_3_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__40269\,
            in1 => \_gnd_net_\,
            in2 => \N__21830\,
            in3 => \_gnd_net_\,
            lcout => \N_317\,
            ltout => \N_317_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI8U0V1_1_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__40632\,
            in1 => \N__40533\,
            in2 => \N__21827\,
            in3 => \N__33754\,
            lcout => \sAddress_RNI8U0V1Z0Z_1\,
            ltout => \sAddress_RNI8U0V1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIETI62_1_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__23836\,
            in1 => \_gnd_net_\,
            in2 => \N__21824\,
            in3 => \_gnd_net_\,
            lcout => \sAddress_RNIETI62Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__40180\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21821\,
            lcout => \sAddress_RNI9IH12Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPointerReset_RNO_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__33755\,
            in1 => \N__23345\,
            in2 => \N__49352\,
            in3 => \N__27092\,
            lcout => OPEN,
            ltout => \N_454_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPointerReset_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001011111110"
        )
    port map (
            in0 => \N__39225\,
            in1 => \N__26006\,
            in2 => \N__21815\,
            in3 => \N__25952\,
            lcout => \sEEPointerResetZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIBH15_4_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40871\,
            in2 => \_gnd_net_\,
            in3 => \N__22610\,
            lcout => OPEN,
            ltout => \N_346_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIUTJC_6_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40410\,
            in1 => \N__21920\,
            in2 => \N__21938\,
            in3 => \N__21890\,
            lcout => OPEN,
            ltout => \un1_spointer11_8_0_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI7G5E2_6_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__23554\,
            in1 => \N__27093\,
            in2 => \N__21935\,
            in3 => \N__33747\,
            lcout => \sAddress_RNI7G5E2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_4_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45387\,
            in2 => \_gnd_net_\,
            in3 => \N__26166\,
            lcout => \sAddressZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52312\,
            ce => \N__23417\,
            sr => \N__51738\
        );

    \sAddress_5_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__26167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45037\,
            lcout => \sAddressZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52312\,
            ce => \N__23417\,
            sr => \N__51738\
        );

    \sAddress_RNIQ63A_0_6_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__22611\,
            in1 => \N__21919\,
            in2 => \N__40900\,
            in3 => \N__21889\,
            lcout => \sEEPonPoff_1_sqmuxa_0_a3_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIFL15_6_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21918\,
            in2 => \_gnd_net_\,
            in3 => \N__21888\,
            lcout => \sDAC_mem_17_1_sqmuxa_0_a2_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_0_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24254\,
            in1 => \N__21859\,
            in2 => \N__24221\,
            in3 => \N__24220\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0\,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51725\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24256\,
            in1 => \N__21845\,
            in2 => \_gnd_net_\,
            in3 => \N__21833\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0\,
            carryout => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1\,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51725\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_2_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24255\,
            in1 => \N__22039\,
            in2 => \_gnd_net_\,
            in3 => \N__22025\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1\,
            carryout => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2\,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51725\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_3_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24286\,
            in2 => \_gnd_net_\,
            in3 => \N__22022\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2\,
            carryout => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3\,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51725\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_4_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24304\,
            in2 => \_gnd_net_\,
            in3 => \N__22019\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3\,
            carryout => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4\,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51725\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_5_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22013\,
            in2 => \_gnd_net_\,
            in3 => \N__22016\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51725\
        );

    \spi_slave_inst.rx_ready_i_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111111101100"
        )
    port map (
            in0 => \N__51223\,
            in1 => \N__22634\,
            in2 => \N__49353\,
            in3 => \N__21993\,
            lcout => spi_mosi_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52292\,
            ce => 'H',
            sr => \N__51714\
        );

    \spi_mosi_ready_prev_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21994\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_mosi_ready_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52292\,
            ce => 'H',
            sr => \N__51714\
        );

    \spi_mosi_ready_prev2_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21971\,
            lcout => \spi_mosi_ready_prevZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52292\,
            ce => 'H',
            sr => \N__51714\
        );

    \spi_mosi_ready_prev3_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21959\,
            lcout => \spi_mosi_ready_prevZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52292\,
            ce => 'H',
            sr => \N__51714\
        );

    \trig_prev_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__22798\,
            in1 => \N__22828\,
            in2 => \_gnd_net_\,
            in3 => \N__22758\,
            lcout => \trig_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52292\,
            ce => 'H',
            sr => \N__51714\
        );

    \sEETrigCounter_RNIR6CE_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22144\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un10_trig_prev_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_done_reg3_i_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22670\,
            lcout => \spi_slave_inst.rx_done_reg3_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52292\,
            ce => 'H',
            sr => \N__51714\
        );

    \un10_trig_prev_cry_0_c_inv_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22121\,
            in2 => \N__22130\,
            in3 => \N__26562\,
            lcout => \sTrigCounter_i_0\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => un10_trig_prev_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_1_c_inv_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22106\,
            in2 => \N__22115\,
            in3 => \N__26949\,
            lcout => \sTrigCounter_i_1\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_0,
            carryout => un10_trig_prev_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_2_c_inv_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22091\,
            in2 => \N__22100\,
            in3 => \N__22858\,
            lcout => \sTrigCounter_i_2\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_1,
            carryout => un10_trig_prev_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_3_c_inv_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22076\,
            in2 => \N__22085\,
            in3 => \N__22843\,
            lcout => \sTrigCounter_i_3\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_2,
            carryout => un10_trig_prev_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_4_c_inv_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22061\,
            in2 => \N__22070\,
            in3 => \N__23071\,
            lcout => \sTrigCounter_i_4\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_3,
            carryout => un10_trig_prev_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_5_c_inv_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23056\,
            in1 => \N__22046\,
            in2 => \N__22055\,
            in3 => \_gnd_net_\,
            lcout => \sTrigCounter_i_5\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_4,
            carryout => un10_trig_prev_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_6_c_inv_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22256\,
            in2 => \N__22265\,
            in3 => \N__23041\,
            lcout => \sTrigCounter_i_6\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_5,
            carryout => un10_trig_prev_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_7_c_inv_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22241\,
            in2 => \N__22250\,
            in3 => \N__23026\,
            lcout => \sTrigCounter_i_7\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_6,
            carryout => un10_trig_prev_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_8_c_inv_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22226\,
            in2 => \N__22235\,
            in3 => \N__23011\,
            lcout => \sTrigCounter_i_8\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => un10_trig_prev_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_9_c_inv_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22211\,
            in2 => \N__22220\,
            in3 => \N__22996\,
            lcout => \sTrigCounter_i_9\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_8,
            carryout => un10_trig_prev_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_10_c_inv_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22981\,
            in1 => \N__22196\,
            in2 => \N__22205\,
            in3 => \_gnd_net_\,
            lcout => \sTrigCounter_i_10\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_9,
            carryout => un10_trig_prev_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_11_c_inv_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22181\,
            in2 => \N__22190\,
            in3 => \N__22966\,
            lcout => \sTrigCounter_i_11\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_10,
            carryout => un10_trig_prev_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_12_c_inv_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22951\,
            in1 => \N__22166\,
            in2 => \N__22175\,
            in3 => \_gnd_net_\,
            lcout => \sTrigCounter_i_12\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_11,
            carryout => un10_trig_prev_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_13_c_inv_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22151\,
            in2 => \N__22160\,
            in3 => \N__23128\,
            lcout => \sTrigCounter_i_13\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_12,
            carryout => un10_trig_prev_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_14_c_inv_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22301\,
            in2 => \N__22310\,
            in3 => \N__23113\,
            lcout => \sTrigCounter_i_14\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_13,
            carryout => un10_trig_prev_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_15_c_inv_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22286\,
            in2 => \N__22295\,
            in3 => \N__23095\,
            lcout => \sTrigCounter_i_15\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_14,
            carryout => un10_trig_prev_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_15_THRU_LUT4_0_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22280\,
            lcout => \un10_trig_prev_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_rpi_ibuf_RNI4GQD1_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49354\,
            in2 => \_gnd_net_\,
            in3 => \N__22277\,
            lcout => \N_82_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_prev_RNIIHS91_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110110000"
        )
    port map (
            in0 => \N__23656\,
            in1 => \N__23720\,
            in2 => \N__22381\,
            in3 => \N__22726\,
            lcout => \N_173\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_ft_ibuf_RNI4OFN_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__22785\,
            in1 => \N__22829\,
            in2 => \_gnd_net_\,
            in3 => \N__22766\,
            lcout => un3_trig_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_done_neg_sclk_i_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__51227\,
            in1 => \N__22576\,
            in2 => \_gnd_net_\,
            in3 => \N__24257\,
            lcout => \spi_slave_inst.rx_done_neg_sclk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi_slave_inst.rx_done_neg_sclk_iC_net\,
            ce => 'H',
            sr => \N__51681\
        );

    \sEEADC_freq_RNICSIA1_4_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__22271\,
            in1 => \N__43052\,
            in2 => \N__22364\,
            in3 => \N__43079\,
            lcout => \un11_sacqtime_NE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEADC_freq_4_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45576\,
            lcout => \sEEADC_freqZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52343\,
            ce => \N__49561\,
            sr => \_gnd_net_\
        );

    \sTrigInternal_RNO_2_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001111"
        )
    port map (
            in0 => \N__23655\,
            in1 => \N__23719\,
            in2 => \N__22385\,
            in3 => \N__22727\,
            lcout => un1_scounter_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEADC_freq_5_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45009\,
            lcout => \sEEADC_freqZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52343\,
            ce => \N__49561\,
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_1_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22480\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48259\,
            ce => \N__48231\,
            sr => \N__51812\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_0_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22355\,
            in1 => \N__48011\,
            in2 => \_gnd_net_\,
            in3 => \N__22337\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48259\,
            ce => \N__48231\,
            sr => \N__51812\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_11_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24053\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48455\,
            ce => 'H',
            sr => \N__51805\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_6_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22414\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48260\,
            ce => \N__48236\,
            sr => \N__51794\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_2_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22465\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48260\,
            ce => \N__48236\,
            sr => \N__51794\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_3_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22450\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48260\,
            ce => \N__48236\,
            sr => \N__51794\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_4_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22438\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48260\,
            ce => \N__48236\,
            sr => \N__51794\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_5_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22426\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48260\,
            ce => \N__48236\,
            sr => \N__51794\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_7_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22402\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48260\,
            ce => \N__48236\,
            sr => \N__51794\
        );

    \spi_slave_inst.rxdata_reg_i_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22484\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => spi_data_mosi_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52344\,
            ce => \N__22565\,
            sr => \N__51780\
        );

    \spi_slave_inst.rxdata_reg_i_1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => spi_data_mosi_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52344\,
            ce => \N__22565\,
            sr => \N__51780\
        );

    \spi_slave_inst.rxdata_reg_i_2_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22451\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => spi_data_mosi_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52344\,
            ce => \N__22565\,
            sr => \N__51780\
        );

    \spi_slave_inst.rxdata_reg_i_3_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22439\,
            lcout => spi_data_mosi_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52344\,
            ce => \N__22565\,
            sr => \N__51780\
        );

    \spi_slave_inst.rxdata_reg_i_4_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22427\,
            lcout => spi_data_mosi_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52344\,
            ce => \N__22565\,
            sr => \N__51780\
        );

    \spi_slave_inst.rxdata_reg_i_5_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22415\,
            lcout => spi_data_mosi_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52344\,
            ce => \N__22565\,
            sr => \N__51780\
        );

    \spi_slave_inst.rxdata_reg_i_6_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22403\,
            lcout => spi_data_mosi_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52344\,
            ce => \N__22565\,
            sr => \N__51780\
        );

    \spi_slave_inst.rxdata_reg_i_7_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22391\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => spi_data_mosi_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52344\,
            ce => \N__22565\,
            sr => \N__51780\
        );

    \sDAC_mem_11_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45978\,
            lcout => \sDAC_mem_11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52335\,
            ce => \N__22493\,
            sr => \N__51765\
        );

    \sDAC_mem_11_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50716\,
            lcout => \sDAC_mem_11Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52335\,
            ce => \N__22493\,
            sr => \N__51765\
        );

    \sDAC_mem_11_2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47119\,
            lcout => \sDAC_mem_11Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52335\,
            ce => \N__22493\,
            sr => \N__51765\
        );

    \sDAC_mem_11_3_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46519\,
            lcout => \sDAC_mem_11Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52335\,
            ce => \N__22493\,
            sr => \N__51765\
        );

    \sDAC_mem_11_4_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45388\,
            lcout => \sDAC_mem_11Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52335\,
            ce => \N__22493\,
            sr => \N__51765\
        );

    \sDAC_mem_11_5_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44731\,
            lcout => \sDAC_mem_11Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52335\,
            ce => \N__22493\,
            sr => \N__51765\
        );

    \sDAC_mem_11_6_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50168\,
            lcout => \sDAC_mem_11Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52335\,
            ce => \N__22493\,
            sr => \N__51765\
        );

    \sDAC_mem_11_7_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49655\,
            lcout => \sDAC_mem_11Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52335\,
            ce => \N__22493\,
            sr => \N__51765\
        );

    \sAddress_RNI9IH12_15_5_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__34857\,
            in1 => \N__40306\,
            in2 => \N__40998\,
            in3 => \N__40753\,
            lcout => \sDAC_mem_11_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_19_5_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__40751\,
            in1 => \N__40294\,
            in2 => \N__40976\,
            in3 => \N__34858\,
            lcout => \sDAC_mem_3_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_3_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46603\,
            in2 => \_gnd_net_\,
            in3 => \N__26163\,
            lcout => \sAddressZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52325\,
            ce => \N__23413\,
            sr => \N__51752\
        );

    \sEETrigInternal_RNO_2_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__40307\,
            in1 => \N__34853\,
            in2 => \_gnd_net_\,
            in3 => \N__23445\,
            lcout => OPEN,
            ltout => \N_344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigInternal_RNO_1_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001101"
        )
    port map (
            in0 => \N__26087\,
            in1 => \N__23705\,
            in2 => \N__22547\,
            in3 => \N__25945\,
            lcout => \sEETrigInternal_3_iv_0_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_6_5_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__40752\,
            in1 => \N__40295\,
            in2 => \N__40977\,
            in3 => \N__34859\,
            lcout => \sDAC_mem_35_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigInternal_RNO_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__27091\,
            in1 => \N__23704\,
            in2 => \N__34866\,
            in3 => \N__26162\,
            lcout => \N_1631\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEESingleCont_RNO_0_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__26041\,
            in1 => \N__26088\,
            in2 => \N__26184\,
            in3 => \N__27090\,
            lcout => \sEESingleCont_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEESingleCont_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__23490\,
            in1 => \N__22522\,
            in2 => \N__46211\,
            in3 => \N__22532\,
            lcout => \sEESingleContZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52313\,
            ce => 'H',
            sr => \N__51739\
        );

    \sEETrigInternal_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__22508\,
            in1 => \N__26043\,
            in2 => \N__22502\,
            in3 => \N__23706\,
            lcout => \sEETrigInternalZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52313\,
            ce => 'H',
            sr => \N__51739\
        );

    \sEETrigInternal_prev_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23707\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEETrigInternal_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52313\,
            ce => 'H',
            sr => \N__51739\
        );

    \sPointer_1_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011100000111000"
        )
    port map (
            in0 => \N__26089\,
            in1 => \N__26042\,
            in2 => \N__26193\,
            in3 => \_gnd_net_\,
            lcout => \sPointerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52313\,
            ce => 'H',
            sr => \N__51739\
        );

    \sPointer_0_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100100000"
        )
    port map (
            in0 => \N__26044\,
            in1 => \N__26174\,
            in2 => \N__25046\,
            in3 => \N__26090\,
            lcout => \sPointerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52313\,
            ce => 'H',
            sr => \N__51739\
        );

    \spi_slave_inst.rx_done_reg1_i_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51216\,
            in1 => \N__48284\,
            in2 => \_gnd_net_\,
            in3 => \N__22586\,
            lcout => \spi_slave_inst.rx_done_reg1_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52313\,
            ce => 'H',
            sr => \N__51739\
        );

    \spi_slave_inst.rx_done_reg1_i_RNID541_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22555\,
            in2 => \_gnd_net_\,
            in3 => \N__22663\,
            lcout => \spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_done_reg2_i_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22556\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_inst.rx_done_reg2_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52313\,
            ce => 'H',
            sr => \N__51739\
        );

    \sAddress_RNI9IH12_5_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__40895\,
            in1 => \_gnd_net_\,
            in2 => \N__26977\,
            in3 => \N__40744\,
            lcout => \sDAC_mem_37_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_18_5_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__40742\,
            in1 => \N__40407\,
            in2 => \N__23565\,
            in3 => \N__40894\,
            lcout => \sDAC_mem_7_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_0_3_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23340\,
            in1 => \N__40406\,
            in2 => \_gnd_net_\,
            in3 => \N__39970\,
            lcout => \sDAC_mem_32_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_7_5_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__40743\,
            in1 => \N__40409\,
            in2 => \N__23566\,
            in3 => \N__40896\,
            lcout => \sDAC_mem_39_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI6VH7_1_1_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110111"
        )
    port map (
            in0 => \N__40620\,
            in1 => \N__40500\,
            in2 => \N__40195\,
            in3 => \_gnd_net_\,
            lcout => \N_319\,
            ltout => \N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_9_3_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__39971\,
            in1 => \_gnd_net_\,
            in2 => \N__22685\,
            in3 => \N__40408\,
            lcout => \sDAC_mem_23_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_2_1_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__23561\,
            in1 => \N__27094\,
            in2 => \_gnd_net_\,
            in3 => \N__33744\,
            lcout => \sAddress_RNI9IH12_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_ready_i_RNO_0_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__22662\,
            in1 => \_gnd_net_\,
            in2 => \N__22646\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_inst.rx_ready_i_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_10_5_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__40864\,
            in1 => \N__40404\,
            in2 => \N__27061\,
            in3 => \N__40747\,
            lcout => \sDAC_mem_13_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_3_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__40405\,
            in1 => \N__27057\,
            in2 => \_gnd_net_\,
            in3 => \N__39969\,
            lcout => \sDAC_mem_29_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sPointer_RNI5LBD1_0_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__26178\,
            in1 => \N__26091\,
            in2 => \_gnd_net_\,
            in3 => \N__26027\,
            lcout => \sPointer_RNI5LBD1Z0Z_0\,
            ltout => \sPointer_RNI5LBD1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIVREN1_4_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22613\,
            in1 => \N__22622\,
            in2 => \N__22625\,
            in3 => \N__40862\,
            lcout => \sAddress_RNIVREN1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIP2UK1_4_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22621\,
            in1 => \N__22612\,
            in2 => \_gnd_net_\,
            in3 => \N__33732\,
            lcout => \sAddress_RNIP2UK1Z0Z_4\,
            ltout => \sAddress_RNIP2UK1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_11_5_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__40403\,
            in1 => \N__23344\,
            in2 => \N__22589\,
            in3 => \N__40863\,
            lcout => \sDAC_mem_16_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_1_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__40073\,
            in1 => \N__23464\,
            in2 => \_gnd_net_\,
            in3 => \N__33733\,
            lcout => \sEEPon_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_prev_RNIM2UO_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__22827\,
            in1 => \N__22799\,
            in2 => \N__22762\,
            in3 => \N__22716\,
            lcout => g3_0,
            ltout => \g3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigInternal_prev_RNIIHS91_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__23645\,
            in1 => \_gnd_net_\,
            in2 => \N__22703\,
            in3 => \N__23711\,
            lcout => g1_i_a4_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI70I7_1_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__40175\,
            in1 => \N__40402\,
            in2 => \_gnd_net_\,
            in3 => \N__40509\,
            lcout => \sAddress_RNI70I7Z0Z_1\,
            ltout => \sAddress_RNI70I7Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_5_2_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40950\,
            in1 => \N__40647\,
            in2 => \N__22700\,
            in3 => \N__40740\,
            lcout => \sDAC_mem_4_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI25GS1_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__40176\,
            in1 => \N__23461\,
            in2 => \N__40531\,
            in3 => \N__33739\,
            lcout => un1_spointer11_5_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_rpi_ibuf_RNI3E6DF_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001101"
        )
    port map (
            in0 => \N__22697\,
            in1 => \N__22691\,
            in2 => \N__23762\,
            in3 => \N__22925\,
            lcout => un1_reset_rpi_inv_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_15_c_RNIGF876_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23798\,
            in1 => \N__23507\,
            in2 => \N__23849\,
            in3 => \N__22938\,
            lcout => \N_8_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigInternal_RNO_1_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__22940\,
            in1 => \N__23608\,
            in2 => \N__31048\,
            in3 => \N__22893\,
            lcout => \N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_15_c_RNI3GF11_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23607\,
            in1 => \N__25159\,
            in2 => \N__22895\,
            in3 => \N__22939\,
            lcout => \N_178\,
            ltout => \N_178_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigInternal_RNO_0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__22919\,
            in1 => \N__29554\,
            in2 => \N__22907\,
            in3 => \N__22904\,
            lcout => OPEN,
            ltout => \N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigInternal_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110001011100"
        )
    port map (
            in0 => \N__31033\,
            in1 => \N__25206\,
            in2 => \N__22898\,
            in3 => \N__29556\,
            lcout => \sTrigInternalZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52293\,
            ce => 'H',
            sr => \N__51696\
        );

    \sPeriod_prev_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__25160\,
            in1 => \N__29555\,
            in2 => \_gnd_net_\,
            in3 => \N__31034\,
            lcout => \sPeriod_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52293\,
            ce => 'H',
            sr => \N__51696\
        );

    \sPeriod_prev_RNI43A11_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__31569\,
            in1 => \N__30674\,
            in2 => \N__22894\,
            in3 => \N__30888\,
            lcout => g0_13_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26563\,
            in2 => \N__22877\,
            in3 => \N__22876\,
            lcout => \sTrigCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \un1_sTrigCounter_cry_0\,
            clk => \N__52303\,
            ce => 'H',
            sr => \N__23084\
        );

    \sTrigCounter_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26950\,
            in2 => \_gnd_net_\,
            in3 => \N__22862\,
            lcout => \sTrigCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_0\,
            carryout => \un1_sTrigCounter_cry_1\,
            clk => \N__52303\,
            ce => 'H',
            sr => \N__23084\
        );

    \sTrigCounter_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22859\,
            in2 => \_gnd_net_\,
            in3 => \N__22847\,
            lcout => \sTrigCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_1\,
            carryout => \un1_sTrigCounter_cry_2\,
            clk => \N__52303\,
            ce => 'H',
            sr => \N__23084\
        );

    \sTrigCounter_3_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22844\,
            in2 => \_gnd_net_\,
            in3 => \N__22832\,
            lcout => \sTrigCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_2\,
            carryout => \un1_sTrigCounter_cry_3\,
            clk => \N__52303\,
            ce => 'H',
            sr => \N__23084\
        );

    \sTrigCounter_4_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23072\,
            in2 => \_gnd_net_\,
            in3 => \N__23060\,
            lcout => \sTrigCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_3\,
            carryout => \un1_sTrigCounter_cry_4\,
            clk => \N__52303\,
            ce => 'H',
            sr => \N__23084\
        );

    \sTrigCounter_5_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23057\,
            in2 => \_gnd_net_\,
            in3 => \N__23045\,
            lcout => \sTrigCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_4\,
            carryout => \un1_sTrigCounter_cry_5\,
            clk => \N__52303\,
            ce => 'H',
            sr => \N__23084\
        );

    \sTrigCounter_6_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23042\,
            in2 => \_gnd_net_\,
            in3 => \N__23030\,
            lcout => \sTrigCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_5\,
            carryout => \un1_sTrigCounter_cry_6\,
            clk => \N__52303\,
            ce => 'H',
            sr => \N__23084\
        );

    \sTrigCounter_7_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23027\,
            in2 => \_gnd_net_\,
            in3 => \N__23015\,
            lcout => \sTrigCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_6\,
            carryout => \un1_sTrigCounter_cry_7\,
            clk => \N__52303\,
            ce => 'H',
            sr => \N__23084\
        );

    \sTrigCounter_8_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23012\,
            in2 => \_gnd_net_\,
            in3 => \N__23000\,
            lcout => \sTrigCounterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \un1_sTrigCounter_cry_8\,
            clk => \N__52314\,
            ce => 'H',
            sr => \N__23083\
        );

    \sTrigCounter_9_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22997\,
            in2 => \_gnd_net_\,
            in3 => \N__22985\,
            lcout => \sTrigCounterZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_8\,
            carryout => \un1_sTrigCounter_cry_9\,
            clk => \N__52314\,
            ce => 'H',
            sr => \N__23083\
        );

    \sTrigCounter_10_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22982\,
            in2 => \_gnd_net_\,
            in3 => \N__22970\,
            lcout => \sTrigCounterZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_9\,
            carryout => \un1_sTrigCounter_cry_10\,
            clk => \N__52314\,
            ce => 'H',
            sr => \N__23083\
        );

    \sTrigCounter_11_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22967\,
            in2 => \_gnd_net_\,
            in3 => \N__22955\,
            lcout => \sTrigCounterZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_10\,
            carryout => \un1_sTrigCounter_cry_11\,
            clk => \N__52314\,
            ce => 'H',
            sr => \N__23083\
        );

    \sTrigCounter_12_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22952\,
            in2 => \_gnd_net_\,
            in3 => \N__23132\,
            lcout => \sTrigCounterZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_11\,
            carryout => \un1_sTrigCounter_cry_12\,
            clk => \N__52314\,
            ce => 'H',
            sr => \N__23083\
        );

    \sTrigCounter_13_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23129\,
            in2 => \_gnd_net_\,
            in3 => \N__23117\,
            lcout => \sTrigCounterZ0Z_13\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_12\,
            carryout => \un1_sTrigCounter_cry_13\,
            clk => \N__52314\,
            ce => 'H',
            sr => \N__23083\
        );

    \sTrigCounter_14_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23114\,
            in2 => \_gnd_net_\,
            in3 => \N__23102\,
            lcout => \sTrigCounterZ0Z_14\,
            ltout => OPEN,
            carryin => \un1_sTrigCounter_cry_13\,
            carryout => \un1_sTrigCounter_cry_14\,
            clk => \N__52314\,
            ce => 'H',
            sr => \N__23083\
        );

    \sTrigCounter_15_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23096\,
            in2 => \_gnd_net_\,
            in3 => \N__23099\,
            lcout => \sTrigCounterZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52314\,
            ce => 'H',
            sr => \N__23083\
        );

    \sDAC_mem_29_0_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46149\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_29Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52326\,
            ce => \N__23149\,
            sr => \N__51674\
        );

    \sDAC_mem_29_1_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50883\,
            lcout => \sDAC_mem_29Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52326\,
            ce => \N__23149\,
            sr => \N__51674\
        );

    \sDAC_mem_29_2_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47379\,
            lcout => \sDAC_mem_29Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52326\,
            ce => \N__23149\,
            sr => \N__51674\
        );

    \sDAC_mem_29_3_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46650\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_29Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52326\,
            ce => \N__23149\,
            sr => \N__51674\
        );

    \sDAC_mem_29_4_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45574\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_29Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52326\,
            ce => \N__23149\,
            sr => \N__51674\
        );

    \sDAC_mem_29_6_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50329\,
            lcout => \sDAC_mem_29Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52326\,
            ce => \N__23149\,
            sr => \N__51674\
        );

    \sDAC_mem_29_7_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50060\,
            lcout => \sDAC_mem_29Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52326\,
            ce => \N__23149\,
            sr => \N__51674\
        );

    \sDAC_mem_16_0_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46279\,
            lcout => \sDAC_mem_16Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52336\,
            ce => \N__33504\,
            sr => \N__51665\
        );

    \sDAC_mem_16_1_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50881\,
            lcout => \sDAC_mem_16Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52336\,
            ce => \N__33504\,
            sr => \N__51665\
        );

    \sDAC_mem_16_2_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47380\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_16Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52336\,
            ce => \N__33504\,
            sr => \N__51665\
        );

    \sEEPon_0_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46280\,
            lcout => \sEEPonZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52345\,
            ce => \N__23207\,
            sr => \N__51660\
        );

    \sEEPon_1_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50882\,
            lcout => \sEEPonZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52345\,
            ce => \N__23207\,
            sr => \N__51660\
        );

    \sEEPon_2_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47457\,
            lcout => \sEEPonZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52345\,
            ce => \N__23207\,
            sr => \N__51660\
        );

    \sEEPon_3_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46909\,
            lcout => \sEEPonZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52345\,
            ce => \N__23207\,
            sr => \N__51660\
        );

    \sEEPon_4_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45575\,
            lcout => \sEEPonZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52345\,
            ce => \N__23207\,
            sr => \N__51660\
        );

    \sEEPon_5_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45085\,
            lcout => \sEEPonZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52345\,
            ce => \N__23207\,
            sr => \N__51660\
        );

    \sEEPon_6_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50330\,
            lcout => \sEEPonZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52345\,
            ce => \N__23207\,
            sr => \N__51660\
        );

    \sEEPon_7_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49990\,
            lcout => \sEEPonZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52345\,
            ce => \N__23207\,
            sr => \N__51660\
        );

    \spi_master_inst.spi_data_path_u1.tx_ready_i_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011110100"
        )
    port map (
            in0 => \N__23195\,
            in1 => \N__23188\,
            in2 => \N__43888\,
            in3 => \N__47554\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_ready_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48451\,
            ce => 'H',
            sr => \N__51795\
        );

    \spi_master_inst.spi_data_path_u1.tx_done_reg3_i_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23189\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48451\,
            ce => 'H',
            sr => \N__51795\
        );

    \spi_master_inst.spi_data_path_u1.tx_done_reg2_i_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23159\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48451\,
            ce => 'H',
            sr => \N__51795\
        );

    \spi_master_inst.sclk_gen_u0.spi_start_i_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47555\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_master_inst.sclk_gen_u0.spi_start_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48451\,
            ce => 'H',
            sr => \N__51795\
        );

    \spi_master_inst.spi_data_path_u1.tx_done_reg1_i_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23180\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48451\,
            ce => 'H',
            sr => \N__51795\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_4_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31778\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48451\,
            ce => 'H',
            sr => \N__51795\
        );

    \reset_rpi_ibuf_RNIRGF52_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__23300\,
            in1 => \N__27106\,
            in2 => \N__49355\,
            in3 => \N__33768\,
            lcout => \sEEADC_freq_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4Q_12_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25766\,
            in1 => \N__23234\,
            in2 => \_gnd_net_\,
            in3 => \N__24692\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4Q_10_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43847\,
            in1 => \N__23999\,
            in2 => \_gnd_net_\,
            in3 => \N__24691\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_10_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45977\,
            lcout => \sDAC_mem_10Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52337\,
            ce => \N__23264\,
            sr => \N__51766\
        );

    \sDAC_mem_10_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50715\,
            lcout => \sDAC_mem_10Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52337\,
            ce => \N__23264\,
            sr => \N__51766\
        );

    \sDAC_mem_10_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47118\,
            lcout => \sDAC_mem_10Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52337\,
            ce => \N__23264\,
            sr => \N__51766\
        );

    \sDAC_mem_10_3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46518\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_10Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52337\,
            ce => \N__23264\,
            sr => \N__51766\
        );

    \sDAC_mem_10_4_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45224\,
            lcout => \sDAC_mem_10Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52337\,
            ce => \N__23264\,
            sr => \N__51766\
        );

    \sDAC_mem_10_5_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44730\,
            lcout => \sDAC_mem_10Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52337\,
            ce => \N__23264\,
            sr => \N__51766\
        );

    \sDAC_mem_10_6_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50224\,
            lcout => \sDAC_mem_10Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52337\,
            ce => \N__23264\,
            sr => \N__51766\
        );

    \sDAC_mem_10_7_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49654\,
            lcout => \sDAC_mem_10Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52337\,
            ce => \N__23264\,
            sr => \N__51766\
        );

    \sDAC_mem_38_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45979\,
            lcout => \sDAC_mem_38Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52327\,
            ce => \N__23246\,
            sr => \N__51753\
        );

    \sDAC_mem_38_1_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50718\,
            lcout => \sDAC_mem_38Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52327\,
            ce => \N__23246\,
            sr => \N__51753\
        );

    \sDAC_mem_38_2_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47121\,
            lcout => \sDAC_mem_38Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52327\,
            ce => \N__23246\,
            sr => \N__51753\
        );

    \sDAC_mem_38_3_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46521\,
            lcout => \sDAC_mem_38Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52327\,
            ce => \N__23246\,
            sr => \N__51753\
        );

    \sDAC_mem_38_4_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45226\,
            lcout => \sDAC_mem_38Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52327\,
            ce => \N__23246\,
            sr => \N__51753\
        );

    \sDAC_mem_38_5_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44733\,
            lcout => \sDAC_mem_38Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52327\,
            ce => \N__23246\,
            sr => \N__51753\
        );

    \sDAC_mem_38_6_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50170\,
            lcout => \sDAC_mem_38Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52327\,
            ce => \N__23246\,
            sr => \N__51753\
        );

    \sDAC_mem_38_7_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49672\,
            lcout => \sDAC_mem_38Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52327\,
            ce => \N__23246\,
            sr => \N__51753\
        );

    \sAddress_RNI9IH12_12_5_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__40298\,
            in1 => \N__40961\,
            in2 => \N__23298\,
            in3 => \N__40785\,
            lcout => \sDAC_mem_14_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_5_5_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__40786\,
            in1 => \N__23293\,
            in2 => \N__40995\,
            in3 => \N__40300\,
            lcout => \sDAC_mem_38_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_17_5_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40296\,
            in1 => \N__40960\,
            in2 => \N__23299\,
            in3 => \N__40784\,
            lcout => \sDAC_mem_6_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_3_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23294\,
            in1 => \N__40299\,
            in2 => \_gnd_net_\,
            in3 => \N__39997\,
            lcout => \sDAC_mem_30_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI6VH7_3_1_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40120\,
            in2 => \N__40532\,
            in3 => \N__40603\,
            lcout => \sAddress_RNI6VH7_3Z0Z_1\,
            ltout => \sAddress_RNI6VH7_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_7_3_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40297\,
            in2 => \N__23267\,
            in3 => \N__39998\,
            lcout => \sDAC_mem_22_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46015\,
            in2 => \_gnd_net_\,
            in3 => \N__26165\,
            lcout => \sAddressZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52315\,
            ce => \N__23418\,
            sr => \N__51740\
        );

    \sAddress_RNI6VH7_0_1_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111011"
        )
    port map (
            in0 => \N__40604\,
            in1 => \N__40516\,
            in2 => \N__40157\,
            in3 => \_gnd_net_\,
            lcout => \N_333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_16_5_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__40302\,
            in1 => \N__40968\,
            in2 => \N__23834\,
            in3 => \N__40794\,
            lcout => \sDAC_mem_10_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI6VH7_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__40615\,
            in1 => \N__40520\,
            in2 => \_gnd_net_\,
            in3 => \N__40139\,
            lcout => \N_326\,
            ltout => \N_326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_10_3_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40301\,
            in2 => \N__23249\,
            in3 => \N__40002\,
            lcout => \sDAC_mem_18_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_2_5_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__40796\,
            in1 => \N__23824\,
            in2 => \N__40997\,
            in3 => \N__40305\,
            lcout => \sDAC_mem_42_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_8_5_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__40304\,
            in1 => \N__40969\,
            in2 => \N__23835\,
            in3 => \N__40795\,
            lcout => \sDAC_mem_34_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_20_5_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__40793\,
            in1 => \N__23823\,
            in2 => \N__40996\,
            in3 => \N__40303\,
            lcout => \sDAC_mem_2_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_2_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47174\,
            in2 => \_gnd_net_\,
            in3 => \N__26164\,
            lcout => \sAddressZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52304\,
            ce => \N__23422\,
            sr => \N__51726\
        );

    \sAddress_RNI6VH7_5_1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__40616\,
            in1 => \N__40507\,
            in2 => \_gnd_net_\,
            in3 => \N__40158\,
            lcout => \sAddress_RNI6VH7_5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_ready_i_RNIBLID_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49365\,
            in2 => \_gnd_net_\,
            in3 => \N__44570\,
            lcout => \spi_slave_inst.un4_i_wr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_14_5_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__40746\,
            in1 => \N__40385\,
            in2 => \N__40994\,
            in3 => \N__23550\,
            lcout => \sDAC_mem_15_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_ACQ_obuf_RNO_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000100"
        )
    port map (
            in0 => \N__25158\,
            in1 => \N__49364\,
            in2 => \N__25187\,
            in3 => \N__25213\,
            lcout => \LED_ACQ_obuf_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_1_2_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__40618\,
            in1 => \N__23463\,
            in2 => \N__27023\,
            in3 => \N__33743\,
            lcout => \sAddress_RNI9IH12_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_2_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27015\,
            in1 => \N__40619\,
            in2 => \_gnd_net_\,
            in3 => \N__39973\,
            lcout => \sDAC_mem_24_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIAM2A_0_1_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__40617\,
            in1 => \N__40508\,
            in2 => \N__40377\,
            in3 => \N__40159\,
            lcout => \sAddress_RNIAM2A_0Z0Z_1\,
            ltout => \sAddress_RNIAM2A_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_3_5_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40956\,
            in2 => \N__23501\,
            in3 => \N__40745\,
            lcout => \sDAC_mem_5_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIAM2A_1_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100000"
        )
    port map (
            in0 => \N__40161\,
            in1 => \N__40334\,
            in2 => \N__40521\,
            in3 => \N__40646\,
            lcout => \N_445\,
            ltout => \N_445_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__40162\,
            in1 => \N__23462\,
            in2 => \N__23498\,
            in3 => \N__33745\,
            lcout => \sAddress_RNIA6242Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_13_5_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__40336\,
            in1 => \N__40949\,
            in2 => \N__23495\,
            in3 => \N__40741\,
            lcout => \sDAC_mem_12_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_2_3_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23494\,
            in1 => \N__40335\,
            in2 => \_gnd_net_\,
            in3 => \N__39972\,
            lcout => \sDAC_mem_28_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_4_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__40163\,
            in1 => \N__23474\,
            in2 => \N__23468\,
            in3 => \N__33746\,
            lcout => \sAddress_RNIA6242_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50851\,
            in2 => \_gnd_net_\,
            in3 => \N__26196\,
            lcout => \sAddressZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52282\,
            ce => \N__23409\,
            sr => \N__51703\
        );

    \sAddress_RNI6VH7_2_1_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__40645\,
            in1 => \N__40496\,
            in2 => \_gnd_net_\,
            in3 => \N__40160\,
            lcout => \sAddress_RNI6VH7_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIM4BU_20_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33362\,
            in1 => \N__29872\,
            in2 => \N__33165\,
            in3 => \N__29998\,
            lcout => g0_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigInternal_prev_RNIH3OJ1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000100"
        )
    port map (
            in0 => \N__23718\,
            in1 => \N__23666\,
            in2 => \N__23657\,
            in3 => \N__31029\,
            lcout => \sEETrigInternal_prev_RNIH3OJZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sSingleCont_RNIUP5M_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__49253\,
            in1 => \N__30555\,
            in2 => \_gnd_net_\,
            in3 => \N__23606\,
            lcout => g0_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_4_3_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__39991\,
            in1 => \N__40384\,
            in2 => \_gnd_net_\,
            in3 => \N__34867\,
            lcout => \sDAC_mem_27_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIUB4L_12_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31722\,
            in1 => \N__31550\,
            in2 => \N__31468\,
            in3 => \N__31643\,
            lcout => \N_831_16\,
            ltout => \N_831_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIP69T1_10_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__24182\,
            in1 => \N__33053\,
            in2 => \N__23570\,
            in3 => \N__30345\,
            lcout => un1_reset_rpi_inv_2_0_o2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_5_3_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100000"
        )
    port map (
            in0 => \N__40009\,
            in1 => \N__23567\,
            in2 => \N__40412\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_31_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIEQR21_10_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30457\,
            in1 => \N__30563\,
            in2 => \N__30361\,
            in3 => \N__30233\,
            lcout => OPEN,
            ltout => \g0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNID5AA2_5_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24161\,
            in1 => \N__30781\,
            in2 => \N__23519\,
            in3 => \N__30898\,
            lcout => g0_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIN61V1_10_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__24173\,
            in1 => \N__30346\,
            in2 => \N__23516\,
            in3 => \N__30458\,
            lcout => g0_15_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNI3LAJ2_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__24566\,
            in1 => \N__29873\,
            in2 => \N__23858\,
            in3 => \N__30111\,
            lcout => g0_17_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_6_3_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100000"
        )
    port map (
            in0 => \N__40010\,
            in1 => \N__23840\,
            in2 => \N__40411\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_26_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIDCVE1_18_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__25850\,
            in1 => \N__31163\,
            in2 => \N__32951\,
            in3 => \N__30005\,
            lcout => g0_16_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNITBBU_23_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32045\,
            in1 => \N__30667\,
            in2 => \N__31930\,
            in3 => \N__30110\,
            lcout => g1_i_a4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIES4L_0_16_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31161\,
            in1 => \N__31276\,
            in2 => \N__33276\,
            in3 => \N__31366\,
            lcout => OPEN,
            ltout => \g1_i_a4_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNI2KI53_16_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24314\,
            in1 => \N__23792\,
            in2 => \N__23786\,
            in3 => \N__25712\,
            lcout => OPEN,
            ltout => \g1_i_a4_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_rpi_ibuf_RNIUSHQ6_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010101010101"
        )
    port map (
            in0 => \N__49116\,
            in1 => \N__23783\,
            in2 => \N__23774\,
            in3 => \N__23771\,
            lcout => g0_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIRQR25_18_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24575\,
            in1 => \N__23747\,
            in2 => \N__23741\,
            in3 => \N__23726\,
            lcout => \N_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIKSV41_18_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__31160\,
            in1 => \N__24136\,
            in2 => \N__33275\,
            in3 => \N__33048\,
            lcout => g0_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_26_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46343\,
            lcout => \sDAC_mem_26Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52305\,
            ce => \N__28045\,
            sr => \N__51675\
        );

    \sDAC_mem_26_1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51069\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_26Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52305\,
            ce => \N__28045\,
            sr => \N__51675\
        );

    \sDAC_mem_26_3_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46866\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_26Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52305\,
            ce => \N__28045\,
            sr => \N__51675\
        );

    \sDAC_mem_26_4_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45577\,
            lcout => \sDAC_mem_26Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52305\,
            ce => \N__28045\,
            sr => \N__51675\
        );

    \sDAC_mem_26_6_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50495\,
            lcout => \sDAC_mem_26Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52305\,
            ce => \N__28045\,
            sr => \N__51675\
        );

    \sDAC_mem_26_7_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49875\,
            lcout => \sDAC_mem_26Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52305\,
            ce => \N__28045\,
            sr => \N__51675\
        );

    \sDAC_mem_30_0_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46148\,
            lcout => \sDAC_mem_30Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52316\,
            ce => \N__23921\,
            sr => \N__51666\
        );

    \sDAC_mem_30_1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51039\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_30Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52316\,
            ce => \N__23921\,
            sr => \N__51666\
        );

    \sDAC_mem_30_2_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47363\,
            lcout => \sDAC_mem_30Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52316\,
            ce => \N__23921\,
            sr => \N__51666\
        );

    \sDAC_mem_30_3_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46908\,
            lcout => \sDAC_mem_30Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52316\,
            ce => \N__23921\,
            sr => \N__51666\
        );

    \sDAC_mem_30_4_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45578\,
            lcout => \sDAC_mem_30Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52316\,
            ce => \N__23921\,
            sr => \N__51666\
        );

    \sDAC_mem_30_5_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45096\,
            lcout => \sDAC_mem_30Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52316\,
            ce => \N__23921\,
            sr => \N__51666\
        );

    \sDAC_mem_30_6_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50528\,
            lcout => \sDAC_mem_30Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52316\,
            ce => \N__23921\,
            sr => \N__51666\
        );

    \sDAC_mem_30_7_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49876\,
            lcout => \sDAC_mem_30Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52316\,
            ce => \N__23921\,
            sr => \N__51666\
        );

    \sCounter_RNIQB8L_23_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32046\,
            in1 => \N__33161\,
            in2 => \N__31937\,
            in3 => \N__33376\,
            lcout => un21_trig_prev_21_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_0_c_inv_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23909\,
            in1 => \N__30241\,
            in2 => \N__23903\,
            in3 => \_gnd_net_\,
            lcout => \sEEPon_i_0\,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => un7_spon_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_1_c_inv_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23888\,
            in2 => \N__30130\,
            in3 => \N__23894\,
            lcout => \sEEPon_i_1\,
            ltout => OPEN,
            carryin => un7_spon_cry_0,
            carryout => un7_spon_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_2_c_inv_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23882\,
            in1 => \N__23876\,
            in2 => \N__30013\,
            in3 => \_gnd_net_\,
            lcout => \sEEPon_i_2\,
            ltout => OPEN,
            carryin => un7_spon_cry_1,
            carryout => un7_spon_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_3_c_inv_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23870\,
            in1 => \N__23864\,
            in2 => \N__29885\,
            in3 => \_gnd_net_\,
            lcout => \sEEPon_i_3\,
            ltout => OPEN,
            carryin => un7_spon_cry_2,
            carryout => un7_spon_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_4_c_inv_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23963\,
            in2 => \N__31061\,
            in3 => \N__23969\,
            lcout => \sEEPon_i_4\,
            ltout => OPEN,
            carryin => un7_spon_cry_3,
            carryout => un7_spon_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_5_c_inv_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23957\,
            in1 => \N__23951\,
            in2 => \N__30907\,
            in3 => \_gnd_net_\,
            lcout => \sEEPon_i_5\,
            ltout => OPEN,
            carryin => un7_spon_cry_4,
            carryout => un7_spon_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_6_c_inv_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23945\,
            in1 => \N__23939\,
            in2 => \N__30790\,
            in3 => \_gnd_net_\,
            lcout => \sEEPon_i_6\,
            ltout => OPEN,
            carryin => un7_spon_cry_5,
            carryout => un7_spon_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_7_c_inv_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23933\,
            in1 => \N__23927\,
            in2 => \N__30682\,
            in3 => \_gnd_net_\,
            lcout => \sEEPon_i_7\,
            ltout => OPEN,
            carryin => un7_spon_cry_6,
            carryout => un7_spon_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_8_c_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52684\,
            in2 => \N__30575\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => un7_spon_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_9_c_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30466\,
            in2 => \N__52746\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_8,
            carryout => un7_spon_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_10_c_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52672\,
            in2 => \N__30362\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_9,
            carryout => un7_spon_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_11_c_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33058\,
            in2 => \N__52743\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_10,
            carryout => un7_spon_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_12_c_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52676\,
            in2 => \N__31748\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_11,
            carryout => un7_spon_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_13_c_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31660\,
            in2 => \N__52744\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_12,
            carryout => un7_spon_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_14_c_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52680\,
            in2 => \N__31580\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_13,
            carryout => un7_spon_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_15_c_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31480\,
            in2 => \N__52745\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_14,
            carryout => un7_spon_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_16_c_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52747\,
            in2 => \N__31393\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => un7_spon_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_17_c_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31285\,
            in2 => \N__52783\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_16,
            carryout => un7_spon_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_18_c_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52751\,
            in2 => \N__31178\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_17,
            carryout => un7_spon_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_19_c_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33277\,
            in2 => \N__52784\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_18,
            carryout => un7_spon_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_20_c_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52755\,
            in2 => \N__33389\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_19,
            carryout => un7_spon_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_21_c_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33170\,
            in2 => \N__52785\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_20,
            carryout => un7_spon_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_22_c_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52759\,
            in2 => \N__32047\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_21,
            carryout => un7_spon_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_23_c_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31934\,
            in2 => \N__52786\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_22,
            carryout => un7_spon_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pon_obuf_RNO_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__31059\,
            in1 => \N__29561\,
            in2 => \_gnd_net_\,
            in3 => \N__24017\,
            lcout => \pon_obuf_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_10_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23975\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48448\,
            ce => 'H',
            sr => \N__51781\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_15_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24023\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48448\,
            ce => 'H',
            sr => \N__51781\
        );

    \spi_master_inst.spi_data_path_u1.data_in_0_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24782\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48452\,
            ce => \N__43901\,
            sr => \N__51767\
        );

    \spi_master_inst.spi_data_path_u1.data_in_1_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24776\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48452\,
            ce => \N__43901\,
            sr => \N__51767\
        );

    \spi_master_inst.spi_data_path_u1.data_in_10_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29498\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48452\,
            ce => \N__43901\,
            sr => \N__51767\
        );

    \spi_master_inst.spi_data_path_u1.data_in_11_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24770\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48452\,
            ce => \N__43901\,
            sr => \N__51767\
        );

    \spi_master_inst.spi_data_path_u1.data_in_12_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24764\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48452\,
            ce => \N__43901\,
            sr => \N__51767\
        );

    \spi_master_inst.spi_data_path_u1.data_in_13_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24758\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48452\,
            ce => \N__43901\,
            sr => \N__51767\
        );

    \spi_master_inst.spi_data_path_u1.data_in_14_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24752\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48452\,
            ce => \N__43901\,
            sr => \N__51767\
        );

    \spi_master_inst.spi_data_path_u1.data_in_15_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24746\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48452\,
            ce => \N__43901\,
            sr => \N__51767\
        );

    \sDAC_mem_42_0_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46050\,
            lcout => \sDAC_mem_42Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52328\,
            ce => \N__24062\,
            sr => \N__51754\
        );

    \sDAC_mem_42_1_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50814\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_42Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52328\,
            ce => \N__24062\,
            sr => \N__51754\
        );

    \sDAC_mem_42_2_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47169\,
            lcout => \sDAC_mem_42Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52328\,
            ce => \N__24062\,
            sr => \N__51754\
        );

    \sDAC_mem_42_3_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46598\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_42Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52328\,
            ce => \N__24062\,
            sr => \N__51754\
        );

    \sDAC_mem_42_4_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45296\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_42Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52328\,
            ce => \N__24062\,
            sr => \N__51754\
        );

    \sDAC_mem_42_5_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44951\,
            lcout => \sDAC_mem_42Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52328\,
            ce => \N__24062\,
            sr => \N__51754\
        );

    \sDAC_mem_42_6_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50225\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_42Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52328\,
            ce => \N__24062\,
            sr => \N__51754\
        );

    \sDAC_mem_42_7_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49727\,
            lcout => \sDAC_mem_42Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52328\,
            ce => \N__24062\,
            sr => \N__51754\
        );

    \sDAC_mem_14_0_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46210\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_14Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52317\,
            ce => \N__24092\,
            sr => \N__51741\
        );

    \sDAC_mem_14_1_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50896\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_14Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52317\,
            ce => \N__24092\,
            sr => \N__51741\
        );

    \sDAC_mem_14_2_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47275\,
            lcout => \sDAC_mem_14Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52317\,
            ce => \N__24092\,
            sr => \N__51741\
        );

    \sDAC_mem_14_3_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46708\,
            lcout => \sDAC_mem_14Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52317\,
            ce => \N__24092\,
            sr => \N__51741\
        );

    \sDAC_mem_14_4_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45410\,
            lcout => \sDAC_mem_14Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52317\,
            ce => \N__24092\,
            sr => \N__51741\
        );

    \sDAC_mem_14_5_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44928\,
            lcout => \sDAC_mem_14Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52317\,
            ce => \N__24092\,
            sr => \N__51741\
        );

    \sDAC_mem_14_6_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50306\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_14Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52317\,
            ce => \N__24092\,
            sr => \N__51741\
        );

    \sDAC_mem_14_7_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49832\,
            lcout => \sDAC_mem_14Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52317\,
            ce => \N__24092\,
            sr => \N__51741\
        );

    \sEEPeriod_10_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47393\,
            lcout => \sEEPeriodZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52306\,
            ce => \N__24077\,
            sr => \N__51727\
        );

    \sEEPeriod_11_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46829\,
            lcout => \sEEPeriodZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52306\,
            ce => \N__24077\,
            sr => \N__51727\
        );

    \sEEPeriod_12_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45411\,
            lcout => \sEEPeriodZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52306\,
            ce => \N__24077\,
            sr => \N__51727\
        );

    \sEEPeriod_13_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44923\,
            lcout => \sEEPeriodZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52306\,
            ce => \N__24077\,
            sr => \N__51727\
        );

    \sEEPeriod_14_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50307\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52306\,
            ce => \N__24077\,
            sr => \N__51727\
        );

    \sEEPeriod_15_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49789\,
            lcout => \sEEPeriodZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52306\,
            ce => \N__24077\,
            sr => \N__51727\
        );

    \sEEPeriod_8_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46054\,
            lcout => \sEEPeriodZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52306\,
            ce => \N__24077\,
            sr => \N__51727\
        );

    \sEEPeriod_9_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50898\,
            lcout => \sEEPeriodZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52306\,
            ce => \N__24077\,
            sr => \N__51727\
        );

    \sEEPeriod_16_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46391\,
            lcout => \sEEPeriodZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52294\,
            ce => \N__24107\,
            sr => \N__51715\
        );

    \sEEPeriod_17_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50897\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52294\,
            ce => \N__24107\,
            sr => \N__51715\
        );

    \sEEPeriod_18_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47394\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52294\,
            ce => \N__24107\,
            sr => \N__51715\
        );

    \sEEPeriod_19_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46769\,
            lcout => \sEEPeriodZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52294\,
            ce => \N__24107\,
            sr => \N__51715\
        );

    \sEEPeriod_20_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45412\,
            lcout => \sEEPeriodZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52294\,
            ce => \N__24107\,
            sr => \N__51715\
        );

    \sEEPeriod_21_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44929\,
            lcout => \sEEPeriodZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52294\,
            ce => \N__24107\,
            sr => \N__51715\
        );

    \sEEPeriod_22_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50308\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52294\,
            ce => \N__24107\,
            sr => \N__51715\
        );

    \sEEPeriod_23_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49833\,
            lcout => \sEEPeriodZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52294\,
            ce => \N__24107\,
            sr => \N__51715\
        );

    \sDAC_mem_15_0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46375\,
            lcout => \sDAC_mem_15Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52283\,
            ce => \N__24113\,
            sr => \N__51704\
        );

    \sDAC_mem_15_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50899\,
            lcout => \sDAC_mem_15Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52283\,
            ce => \N__24113\,
            sr => \N__51704\
        );

    \sDAC_mem_15_2_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47395\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_15Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52283\,
            ce => \N__24113\,
            sr => \N__51704\
        );

    \sDAC_mem_15_3_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46852\,
            lcout => \sDAC_mem_15Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52283\,
            ce => \N__24113\,
            sr => \N__51704\
        );

    \sDAC_mem_15_4_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45413\,
            lcout => \sDAC_mem_15Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52283\,
            ce => \N__24113\,
            sr => \N__51704\
        );

    \sDAC_mem_15_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__44924\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_15Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52283\,
            ce => \N__24113\,
            sr => \N__51704\
        );

    \sDAC_mem_15_6_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_15Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52283\,
            ce => \N__24113\,
            sr => \N__51704\
        );

    \sDAC_mem_15_7_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49834\,
            lcout => \sDAC_mem_15Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52283\,
            ce => \N__24113\,
            sr => \N__51704\
        );

    \sDAC_mem_18_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46209\,
            lcout => \sDAC_mem_18Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52272\,
            ce => \N__28540\,
            sr => \N__51697\
        );

    \sDAC_mem_18_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50983\,
            lcout => \sDAC_mem_18Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52272\,
            ce => \N__28540\,
            sr => \N__51697\
        );

    \sDAC_mem_18_2_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47461\,
            lcout => \sDAC_mem_18Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52272\,
            ce => \N__28540\,
            sr => \N__51697\
        );

    \sDAC_mem_18_7_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49939\,
            lcout => \sDAC_mem_18Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52272\,
            ce => \N__28540\,
            sr => \N__51697\
        );

    \sCounter_RNI0D9U_10_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30534\,
            in1 => \N__33039\,
            in2 => \N__30446\,
            in3 => \N__30314\,
            lcout => op_gt_op_gt_un13_striginternallto23_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIQB5R1_1_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30081\,
            in1 => \N__29841\,
            in2 => \N__24155\,
            in3 => \N__29970\,
            lcout => OPEN,
            ltout => \op_gt_op_gt_un13_striginternallto23_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIVUR25_16_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24119\,
            in1 => \N__24197\,
            in2 => \N__24185\,
            in3 => \N__24167\,
            lcout => op_gt_op_gt_un13_striginternal_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNI2RIT_8_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__30204\,
            in1 => \N__30422\,
            in2 => \_gnd_net_\,
            in3 => \N__30533\,
            lcout => un1_reset_rpi_inv_2_0_o2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNI9MMP_12_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31630\,
            in1 => \N__31717\,
            in2 => \N__31467\,
            in3 => \N__30205\,
            lcout => g0_13_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIES4L_16_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31336\,
            in1 => \N__33223\,
            in2 => \N__31268\,
            in3 => \N__31123\,
            lcout => un21_trig_prev_21_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIU3NJ_1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30080\,
            in2 => \_gnd_net_\,
            in3 => \N__30634\,
            lcout => g0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNI3SIT_5_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__30675\,
            in1 => \N__30773\,
            in2 => \_gnd_net_\,
            in3 => \N__30880\,
            lcout => \N_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNITA9T1_4_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__31000\,
            in1 => \N__24143\,
            in2 => \N__24137\,
            in3 => \_gnd_net_\,
            lcout => op_gt_op_gt_un13_striginternallto23_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNIJFMR_1_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25489\,
            in2 => \_gnd_net_\,
            in3 => \N__25255\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNILEDN1_7_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25399\,
            in1 => \N__25474\,
            in2 => \N__25436\,
            in3 => \N__25417\,
            lcout => OPEN,
            ltout => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNISEQE3_0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__25460\,
            in1 => \N__25270\,
            in2 => \N__24560\,
            in3 => \N__24557\,
            lcout => \spi_master_inst.sclk_gen_u0.N_158_7\,
            ltout => \spi_master_inst.sclk_gen_u0.N_158_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNO_0_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__24520\,
            in1 => \N__24455\,
            in2 => \N__24392\,
            in3 => \N__24388\,
            lcout => \spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIS7E71_2_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30879\,
            in1 => \N__29851\,
            in2 => \N__30785\,
            in3 => \N__29983\,
            lcout => g2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_RNILK4P2_3_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__24308\,
            in1 => \N__24290\,
            in2 => \_gnd_net_\,
            in3 => \N__24272\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_i6\,
            ltout => \spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3_3_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000111"
        )
    port map (
            in0 => \N__47892\,
            in1 => \N__48006\,
            in2 => \N__24224\,
            in3 => \N__47956\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_RNICH5T1_5_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__42773\,
            in1 => \N__42683\,
            in2 => \N__42740\,
            in3 => \N__38657\,
            lcout => \spi_slave_inst.un23_i_ssn_3\,
            ltout => \spi_slave_inst.un23_i_ssn_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_RNI5DOR2_3_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__48304\,
            in1 => \_gnd_net_\,
            in2 => \N__24200\,
            in3 => \N__48329\,
            lcout => \spi_slave_inst.un23_i_ssn\,
            ltout => \spi_slave_inst.un23_i_ssn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_RNI4ODL3_3_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001101"
        )
    port map (
            in0 => \N__47957\,
            in1 => \N__48007\,
            in2 => \N__24578\,
            in3 => \N__47893\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNI4K6L_23_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31376\,
            in1 => \N__31239\,
            in2 => \N__31905\,
            in3 => \N__31990\,
            lcout => g0_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNI5I9U_16_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30769\,
            in1 => \N__31377\,
            in2 => \N__31267\,
            in3 => \N__30999\,
            lcout => g0_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_31_0_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46338\,
            lcout => \sDAC_mem_31Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52295\,
            ce => \N__24593\,
            sr => \N__51667\
        );

    \sDAC_mem_31_1_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50878\,
            lcout => \sDAC_mem_31Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52295\,
            ce => \N__24593\,
            sr => \N__51667\
        );

    \sDAC_mem_31_2_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47499\,
            lcout => \sDAC_mem_31Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52295\,
            ce => \N__24593\,
            sr => \N__51667\
        );

    \sDAC_mem_31_3_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46913\,
            lcout => \sDAC_mem_31Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52295\,
            ce => \N__24593\,
            sr => \N__51667\
        );

    \sDAC_mem_31_4_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45579\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_31Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52295\,
            ce => \N__24593\,
            sr => \N__51667\
        );

    \sDAC_mem_31_5_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45090\,
            lcout => \sDAC_mem_31Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52295\,
            ce => \N__24593\,
            sr => \N__51667\
        );

    \sDAC_mem_31_6_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50529\,
            lcout => \sDAC_mem_31Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52295\,
            ce => \N__24593\,
            sr => \N__51667\
        );

    \sDAC_mem_31_7_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50028\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_31Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52295\,
            ce => \N__24593\,
            sr => \N__51667\
        );

    \sDAC_mem_24_0_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46322\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_24Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52307\,
            ce => \N__27745\,
            sr => \N__51661\
        );

    \sDAC_mem_24_2_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47500\,
            lcout => \sDAC_mem_24Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52307\,
            ce => \N__27745\,
            sr => \N__51661\
        );

    \sDAC_mem_24_3_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46847\,
            lcout => \sDAC_mem_24Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52307\,
            ce => \N__27745\,
            sr => \N__51661\
        );

    \sDAC_mem_24_5_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45094\,
            lcout => \sDAC_mem_24Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52307\,
            ce => \N__27745\,
            sr => \N__51661\
        );

    \sDAC_mem_24_6_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50391\,
            lcout => \sDAC_mem_24Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52307\,
            ce => \N__27745\,
            sr => \N__51661\
        );

    \sDAC_mem_24_7_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50029\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_24Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52307\,
            ce => \N__27745\,
            sr => \N__51661\
        );

    \sDAC_mem_28_0_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46321\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_28Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52318\,
            ce => \N__37789\,
            sr => \N__51655\
        );

    \sDAC_mem_28_1_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51037\,
            lcout => \sDAC_mem_28Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52318\,
            ce => \N__37789\,
            sr => \N__51655\
        );

    \sDAC_mem_28_3_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46762\,
            lcout => \sDAC_mem_28Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52318\,
            ce => \N__37789\,
            sr => \N__51655\
        );

    \sDAC_mem_28_4_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45580\,
            lcout => \sDAC_mem_28Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52318\,
            ce => \N__37789\,
            sr => \N__51655\
        );

    \sEEDelayACQ_0_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52329\,
            ce => \N__24605\,
            sr => \N__51652\
        );

    \sEEDelayACQ_1_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51038\,
            lcout => \sEEDelayACQZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52329\,
            ce => \N__24605\,
            sr => \N__51652\
        );

    \sEEDelayACQ_2_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47502\,
            lcout => \sEEDelayACQZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52329\,
            ce => \N__24605\,
            sr => \N__51652\
        );

    \sEEDelayACQ_3_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46851\,
            lcout => \sEEDelayACQZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52329\,
            ce => \N__24605\,
            sr => \N__51652\
        );

    \sEEDelayACQ_4_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52329\,
            ce => \N__24605\,
            sr => \N__51652\
        );

    \sEEDelayACQ_5_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45095\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52329\,
            ce => \N__24605\,
            sr => \N__51652\
        );

    \sEEDelayACQ_6_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50392\,
            lcout => \sEEDelayACQZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52329\,
            ce => \N__24605\,
            sr => \N__51652\
        );

    \sEEDelayACQ_7_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50031\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52329\,
            ce => \N__24605\,
            sr => \N__51652\
        );

    \sEEDelayACQ_10_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47512\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52338\,
            ce => \N__24740\,
            sr => \N__51649\
        );

    \sEEDelayACQ_11_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46924\,
            lcout => \sEEDelayACQZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52338\,
            ce => \N__24740\,
            sr => \N__51649\
        );

    \sEEDelayACQ_12_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45604\,
            lcout => \sEEDelayACQZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52338\,
            ce => \N__24740\,
            sr => \N__51649\
        );

    \sEEDelayACQ_13_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45116\,
            lcout => \sEEDelayACQZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52338\,
            ce => \N__24740\,
            sr => \N__51649\
        );

    \sEEDelayACQ_14_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50467\,
            lcout => \sEEDelayACQZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52338\,
            ce => \N__24740\,
            sr => \N__51649\
        );

    \sEEDelayACQ_15_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50051\,
            lcout => \sEEDelayACQZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52338\,
            ce => \N__24740\,
            sr => \N__51649\
        );

    \sEEDelayACQ_8_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46331\,
            lcout => \sEEDelayACQZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52338\,
            ce => \N__24740\,
            sr => \N__51649\
        );

    \sEEDelayACQ_9_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51030\,
            lcout => \sEEDelayACQZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52338\,
            ce => \N__24740\,
            sr => \N__51649\
        );

    \reset_rpi_ibuf_RNIIUT3_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__49246\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LED3_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4Q_15_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24710\,
            in1 => \N__25754\,
            in2 => \_gnd_net_\,
            in3 => \N__24704\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_0_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48449\,
            ce => \N__43958\,
            sr => \N__51755\
        );

    \sDAC_data_1_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48449\,
            ce => \N__43958\,
            sr => \N__51755\
        );

    \sDAC_data_11_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48449\,
            ce => \N__43958\,
            sr => \N__51755\
        );

    \sDAC_data_12_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52649\,
            lcout => \sDAC_dataZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48449\,
            ce => \N__43958\,
            sr => \N__51755\
        );

    \sDAC_data_13_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__52650\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_dataZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48449\,
            ce => \N__43958\,
            sr => \N__51755\
        );

    \sDAC_data_14_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48449\,
            ce => \N__43958\,
            sr => \N__51755\
        );

    \sDAC_data_15_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48449\,
            ce => \N__43958\,
            sr => \N__51755\
        );

    \sEEPeriod_0_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46043\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52319\,
            ce => \N__24836\,
            sr => \N__51742\
        );

    \sEEPeriod_1_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50892\,
            lcout => \sEEPeriodZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52319\,
            ce => \N__24836\,
            sr => \N__51742\
        );

    \sEEPeriod_2_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47170\,
            lcout => \sEEPeriodZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52319\,
            ce => \N__24836\,
            sr => \N__51742\
        );

    \sEEPeriod_3_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46599\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52319\,
            ce => \N__24836\,
            sr => \N__51742\
        );

    \sEEPeriod_4_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45297\,
            lcout => \sEEPeriodZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52319\,
            ce => \N__24836\,
            sr => \N__51742\
        );

    \sEEPeriod_5_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44763\,
            lcout => \sEEPeriodZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52319\,
            ce => \N__24836\,
            sr => \N__51742\
        );

    \sEEPeriod_6_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50317\,
            lcout => \sEEPeriodZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52319\,
            ce => \N__24836\,
            sr => \N__51742\
        );

    \sEEPeriod_7_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49831\,
            lcout => \sEEPeriodZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52319\,
            ce => \N__24836\,
            sr => \N__51742\
        );

    \un4_speriod_cry_0_c_inv_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24818\,
            in2 => \N__30237\,
            in3 => \N__24824\,
            lcout => \sEEPeriod_i_0\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => un4_speriod_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_1_c_inv_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24806\,
            in2 => \N__30117\,
            in3 => \N__24812\,
            lcout => \sEEPeriod_i_1\,
            ltout => OPEN,
            carryin => un4_speriod_cry_0,
            carryout => un4_speriod_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_2_c_inv_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24794\,
            in2 => \N__30006\,
            in3 => \N__24800\,
            lcout => \sEEPeriod_i_2\,
            ltout => OPEN,
            carryin => un4_speriod_cry_1,
            carryout => un4_speriod_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_3_c_inv_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24929\,
            in2 => \N__29877\,
            in3 => \N__24788\,
            lcout => \sEEPeriod_i_3\,
            ltout => OPEN,
            carryin => un4_speriod_cry_2,
            carryout => un4_speriod_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_4_c_inv_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24917\,
            in2 => \N__31016\,
            in3 => \N__24923\,
            lcout => \sEEPeriod_i_4\,
            ltout => OPEN,
            carryin => un4_speriod_cry_3,
            carryout => un4_speriod_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_5_c_inv_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24911\,
            in1 => \N__24905\,
            in2 => \N__30899\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriod_i_5\,
            ltout => OPEN,
            carryin => un4_speriod_cry_4,
            carryout => un4_speriod_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_6_c_inv_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24893\,
            in2 => \N__30774\,
            in3 => \N__24899\,
            lcout => \sEEPeriod_i_6\,
            ltout => OPEN,
            carryin => un4_speriod_cry_5,
            carryout => un4_speriod_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_7_c_inv_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30650\,
            in2 => \N__24881\,
            in3 => \N__24887\,
            lcout => \sEEPeriod_i_7\,
            ltout => OPEN,
            carryin => un4_speriod_cry_6,
            carryout => un4_speriod_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_8_c_inv_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24866\,
            in2 => \N__30570\,
            in3 => \N__24872\,
            lcout => \sEEPeriod_i_8\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => un4_speriod_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_9_c_inv_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24854\,
            in2 => \N__30465\,
            in3 => \N__24860\,
            lcout => \sEEPeriod_i_9\,
            ltout => OPEN,
            carryin => un4_speriod_cry_8,
            carryout => un4_speriod_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_10_c_inv_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24842\,
            in2 => \N__30353\,
            in3 => \N__24848\,
            lcout => \sEEPeriod_i_10\,
            ltout => OPEN,
            carryin => un4_speriod_cry_9,
            carryout => un4_speriod_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_11_c_inv_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25019\,
            in2 => \N__33057\,
            in3 => \N__25025\,
            lcout => \sEEPeriod_i_11\,
            ltout => OPEN,
            carryin => un4_speriod_cry_10,
            carryout => un4_speriod_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_12_c_inv_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25013\,
            in1 => \N__25007\,
            in2 => \N__31733\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriod_i_12\,
            ltout => OPEN,
            carryin => un4_speriod_cry_11,
            carryout => un4_speriod_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_13_c_inv_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25001\,
            in1 => \N__24995\,
            in2 => \N__31658\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriod_i_13\,
            ltout => OPEN,
            carryin => un4_speriod_cry_12,
            carryout => un4_speriod_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_14_c_inv_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24983\,
            in2 => \N__31573\,
            in3 => \N__24989\,
            lcout => \sEEPeriod_i_14\,
            ltout => OPEN,
            carryin => un4_speriod_cry_13,
            carryout => un4_speriod_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_15_c_inv_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24977\,
            in1 => \N__24971\,
            in2 => \N__31479\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriod_i_15\,
            ltout => OPEN,
            carryin => un4_speriod_cry_14,
            carryout => un4_speriod_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_16_c_inv_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24959\,
            in2 => \N__31387\,
            in3 => \N__24965\,
            lcout => \sEEPeriod_i_16\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => un4_speriod_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_17_c_inv_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24947\,
            in2 => \N__31286\,
            in3 => \N__24953\,
            lcout => \sEEPeriod_i_17\,
            ltout => OPEN,
            carryin => un4_speriod_cry_16,
            carryout => un4_speriod_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_18_c_inv_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24935\,
            in2 => \N__31177\,
            in3 => \N__24941\,
            lcout => \sEEPeriod_i_18\,
            ltout => OPEN,
            carryin => un4_speriod_cry_17,
            carryout => un4_speriod_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_19_c_inv_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25103\,
            in2 => \N__33278\,
            in3 => \N__25109\,
            lcout => \sEEPeriod_i_19\,
            ltout => OPEN,
            carryin => un4_speriod_cry_18,
            carryout => un4_speriod_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_20_c_inv_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25091\,
            in2 => \N__33380\,
            in3 => \N__25097\,
            lcout => \sEEPeriod_i_20\,
            ltout => OPEN,
            carryin => un4_speriod_cry_19,
            carryout => un4_speriod_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_21_c_inv_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25085\,
            in1 => \N__25079\,
            in2 => \N__33166\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriod_i_21\,
            ltout => OPEN,
            carryin => un4_speriod_cry_20,
            carryout => un4_speriod_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_22_c_inv_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25067\,
            in2 => \N__32041\,
            in3 => \N__25073\,
            lcout => \sEEPeriod_i_22\,
            ltout => OPEN,
            carryin => un4_speriod_cry_21,
            carryout => un4_speriod_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_23_c_inv_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25055\,
            in2 => \N__31935\,
            in3 => \N__25061\,
            lcout => \sEEPeriod_i_23\,
            ltout => OPEN,
            carryin => un4_speriod_cry_22,
            carryout => un4_speriod_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_23_THRU_LUT4_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25049\,
            lcout => \un4_speriod_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sPointer_RNO_0_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__46770\,
            in1 => \N__25964\,
            in2 => \N__45481\,
            in3 => \N__25031\,
            lcout => un1_spointer11_2_0_0_a2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sPointer_RNO_1_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50305\,
            in2 => \_gnd_net_\,
            in3 => \N__47244\,
            lcout => un1_spointer11_2_0_0_a2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigInternal_RNIMEFL5_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001111"
        )
    port map (
            in0 => \N__25214\,
            in1 => \N__25183\,
            in2 => \N__49363\,
            in3 => \N__25152\,
            lcout => \LED_ACQ_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25347\,
            in1 => \N__30206\,
            in2 => \_gnd_net_\,
            in3 => \N__25133\,
            lcout => un7_spon_0,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \sCounter_cry_0\,
            clk => \N__52262\,
            ce => 'H',
            sr => \N__51689\
        );

    \sCounter_1_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25360\,
            in1 => \N__30089\,
            in2 => \_gnd_net_\,
            in3 => \N__25130\,
            lcout => un7_spon_1,
            ltout => OPEN,
            carryin => \sCounter_cry_0\,
            carryout => \sCounter_cry_1\,
            clk => \N__52262\,
            ce => 'H',
            sr => \N__51689\
        );

    \sCounter_2_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25348\,
            in1 => \N__29969\,
            in2 => \_gnd_net_\,
            in3 => \N__25127\,
            lcout => un7_spon_2,
            ltout => OPEN,
            carryin => \sCounter_cry_1\,
            carryout => \sCounter_cry_2\,
            clk => \N__52262\,
            ce => 'H',
            sr => \N__51689\
        );

    \sCounter_3_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25361\,
            in1 => \N__29840\,
            in2 => \_gnd_net_\,
            in3 => \N__25124\,
            lcout => un7_spon_3,
            ltout => OPEN,
            carryin => \sCounter_cry_2\,
            carryout => \sCounter_cry_3\,
            clk => \N__52262\,
            ce => 'H',
            sr => \N__51689\
        );

    \sCounter_4_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25349\,
            in1 => \N__30984\,
            in2 => \_gnd_net_\,
            in3 => \N__25121\,
            lcout => un7_spon_4,
            ltout => OPEN,
            carryin => \sCounter_cry_3\,
            carryout => \sCounter_cry_4\,
            clk => \N__52262\,
            ce => 'H',
            sr => \N__51689\
        );

    \sCounter_5_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25362\,
            in1 => \N__30863\,
            in2 => \_gnd_net_\,
            in3 => \N__25118\,
            lcout => un7_spon_5,
            ltout => OPEN,
            carryin => \sCounter_cry_4\,
            carryout => \sCounter_cry_5\,
            clk => \N__52262\,
            ce => 'H',
            sr => \N__51689\
        );

    \sCounter_6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25350\,
            in1 => \N__30752\,
            in2 => \_gnd_net_\,
            in3 => \N__25115\,
            lcout => un7_spon_6,
            ltout => OPEN,
            carryin => \sCounter_cry_5\,
            carryout => \sCounter_cry_6\,
            clk => \N__52262\,
            ce => 'H',
            sr => \N__51689\
        );

    \sCounter_7_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25363\,
            in1 => \N__30649\,
            in2 => \_gnd_net_\,
            in3 => \N__25112\,
            lcout => un7_spon_7,
            ltout => OPEN,
            carryin => \sCounter_cry_6\,
            carryout => \sCounter_cry_7\,
            clk => \N__52262\,
            ce => 'H',
            sr => \N__51689\
        );

    \sCounter_8_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25354\,
            in1 => \N__30541\,
            in2 => \_gnd_net_\,
            in3 => \N__25241\,
            lcout => un7_spon_8,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \sCounter_cry_8\,
            clk => \N__52251\,
            ce => 'H',
            sr => \N__51682\
        );

    \sCounter_9_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25367\,
            in1 => \N__30426\,
            in2 => \_gnd_net_\,
            in3 => \N__25238\,
            lcout => un7_spon_9,
            ltout => OPEN,
            carryin => \sCounter_cry_8\,
            carryout => \sCounter_cry_9\,
            clk => \N__52251\,
            ce => 'H',
            sr => \N__51682\
        );

    \sCounter_10_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25351\,
            in1 => \N__30315\,
            in2 => \_gnd_net_\,
            in3 => \N__25235\,
            lcout => un7_spon_10,
            ltout => OPEN,
            carryin => \sCounter_cry_9\,
            carryout => \sCounter_cry_10\,
            clk => \N__52251\,
            ce => 'H',
            sr => \N__51682\
        );

    \sCounter_11_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25364\,
            in1 => \N__33017\,
            in2 => \_gnd_net_\,
            in3 => \N__25232\,
            lcout => un7_spon_11,
            ltout => OPEN,
            carryin => \sCounter_cry_10\,
            carryout => \sCounter_cry_11\,
            clk => \N__52251\,
            ce => 'H',
            sr => \N__51682\
        );

    \sCounter_12_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25352\,
            in1 => \N__31718\,
            in2 => \_gnd_net_\,
            in3 => \N__25229\,
            lcout => un7_spon_12,
            ltout => OPEN,
            carryin => \sCounter_cry_11\,
            carryout => \sCounter_cry_12\,
            clk => \N__52251\,
            ce => 'H',
            sr => \N__51682\
        );

    \sCounter_13_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25365\,
            in1 => \N__31645\,
            in2 => \_gnd_net_\,
            in3 => \N__25226\,
            lcout => un7_spon_13,
            ltout => OPEN,
            carryin => \sCounter_cry_12\,
            carryout => \sCounter_cry_13\,
            clk => \N__52251\,
            ce => 'H',
            sr => \N__51682\
        );

    \sCounter_14_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25353\,
            in1 => \N__31537\,
            in2 => \_gnd_net_\,
            in3 => \N__25223\,
            lcout => un7_spon_14,
            ltout => OPEN,
            carryin => \sCounter_cry_13\,
            carryout => \sCounter_cry_14\,
            clk => \N__52251\,
            ce => 'H',
            sr => \N__51682\
        );

    \sCounter_15_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25366\,
            in1 => \N__31450\,
            in2 => \_gnd_net_\,
            in3 => \N__25220\,
            lcout => un7_spon_15,
            ltout => OPEN,
            carryin => \sCounter_cry_14\,
            carryout => \sCounter_cry_15\,
            clk => \N__52251\,
            ce => 'H',
            sr => \N__51682\
        );

    \sCounter_16_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25355\,
            in1 => \N__31337\,
            in2 => \_gnd_net_\,
            in3 => \N__25217\,
            lcout => un7_spon_16,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \sCounter_cry_16\,
            clk => \N__52263\,
            ce => 'H',
            sr => \N__51676\
        );

    \sCounter_17_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25368\,
            in1 => \N__31261\,
            in2 => \_gnd_net_\,
            in3 => \N__25388\,
            lcout => un7_spon_17,
            ltout => OPEN,
            carryin => \sCounter_cry_16\,
            carryout => \sCounter_cry_17\,
            clk => \N__52263\,
            ce => 'H',
            sr => \N__51676\
        );

    \sCounter_18_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25356\,
            in1 => \N__31124\,
            in2 => \_gnd_net_\,
            in3 => \N__25385\,
            lcout => un7_spon_18,
            ltout => OPEN,
            carryin => \sCounter_cry_17\,
            carryout => \sCounter_cry_18\,
            clk => \N__52263\,
            ce => 'H',
            sr => \N__51676\
        );

    \sCounter_19_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25369\,
            in1 => \N__33224\,
            in2 => \_gnd_net_\,
            in3 => \N__25382\,
            lcout => un7_spon_19,
            ltout => OPEN,
            carryin => \sCounter_cry_18\,
            carryout => \sCounter_cry_19\,
            clk => \N__52263\,
            ce => 'H',
            sr => \N__51676\
        );

    \sCounter_20_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25357\,
            in1 => \N__33331\,
            in2 => \_gnd_net_\,
            in3 => \N__25379\,
            lcout => un7_spon_20,
            ltout => OPEN,
            carryin => \sCounter_cry_19\,
            carryout => \sCounter_cry_20\,
            clk => \N__52263\,
            ce => 'H',
            sr => \N__51676\
        );

    \sCounter_21_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25370\,
            in1 => \N__33115\,
            in2 => \_gnd_net_\,
            in3 => \N__25376\,
            lcout => un7_spon_21,
            ltout => OPEN,
            carryin => \sCounter_cry_20\,
            carryout => \sCounter_cry_21\,
            clk => \N__52263\,
            ce => 'H',
            sr => \N__51676\
        );

    \sCounter_22_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25358\,
            in1 => \N__31991\,
            in2 => \_gnd_net_\,
            in3 => \N__25373\,
            lcout => un7_spon_22,
            ltout => OPEN,
            carryin => \sCounter_cry_21\,
            carryout => \sCounter_cry_22\,
            clk => \N__52263\,
            ce => 'H',
            sr => \N__51676\
        );

    \sCounter_23_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__31882\,
            in1 => \N__25359\,
            in2 => \_gnd_net_\,
            in3 => \N__25274\,
            lcout => un7_spon_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52263\,
            ce => 'H',
            sr => \N__51676\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27927\,
            in1 => \N__25271\,
            in2 => \_gnd_net_\,
            in3 => \N__25259\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0\,
            clk => \N__48472\,
            ce => \N__27968\,
            sr => \N__51668\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27922\,
            in1 => \N__25256\,
            in2 => \_gnd_net_\,
            in3 => \N__25244\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1\,
            clk => \N__48472\,
            ce => \N__27968\,
            sr => \N__51668\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_2_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27928\,
            in1 => \N__25490\,
            in2 => \_gnd_net_\,
            in3 => \N__25478\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2\,
            clk => \N__48472\,
            ce => \N__27968\,
            sr => \N__51668\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_3_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27923\,
            in1 => \N__25475\,
            in2 => \_gnd_net_\,
            in3 => \N__25463\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3\,
            clk => \N__48472\,
            ce => \N__27968\,
            sr => \N__51668\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_4_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27929\,
            in1 => \N__25453\,
            in2 => \_gnd_net_\,
            in3 => \N__25439\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4\,
            clk => \N__48472\,
            ce => \N__27968\,
            sr => \N__51668\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_5_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27924\,
            in1 => \N__25435\,
            in2 => \_gnd_net_\,
            in3 => \N__25421\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5\,
            clk => \N__48472\,
            ce => \N__27968\,
            sr => \N__51668\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_6_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27925\,
            in1 => \N__25418\,
            in2 => \_gnd_net_\,
            in3 => \N__25406\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6\,
            clk => \N__48472\,
            ce => \N__27968\,
            sr => \N__51668\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_7_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__25400\,
            in1 => \N__27926\,
            in2 => \_gnd_net_\,
            in3 => \N__25403\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48472\,
            ce => \N__27968\,
            sr => \N__51668\
        );

    \sEEPoff_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46342\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPoffZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52284\,
            ce => \N__25496\,
            sr => \N__51662\
        );

    \sEEPoff_1_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50879\,
            lcout => \sEEPoffZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52284\,
            ce => \N__25496\,
            sr => \N__51662\
        );

    \sEEPoff_2_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47501\,
            lcout => \sEEPoffZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52284\,
            ce => \N__25496\,
            sr => \N__51662\
        );

    \sEEPoff_3_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46914\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPoffZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52284\,
            ce => \N__25496\,
            sr => \N__51662\
        );

    \sEEPoff_4_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45567\,
            lcout => \sEEPoffZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52284\,
            ce => \N__25496\,
            sr => \N__51662\
        );

    \sEEPoff_5_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45089\,
            lcout => \sEEPoffZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52284\,
            ce => \N__25496\,
            sr => \N__51662\
        );

    \sEEPoff_6_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50530\,
            lcout => \sEEPoffZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52284\,
            ce => \N__25496\,
            sr => \N__51662\
        );

    \sEEPoff_7_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50030\,
            lcout => \sEEPoffZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52284\,
            ce => \N__25496\,
            sr => \N__51662\
        );

    \sAddress_RNIA6242_0_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__40190\,
            in1 => \N__25521\,
            in2 => \N__40669\,
            in3 => \N__40433\,
            lcout => \sAddress_RNIA6242_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_1_0_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__25520\,
            in1 => \N__40654\,
            in2 => \N__40438\,
            in3 => \N__40189\,
            lcout => \sAddress_RNIA6242_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_2_0_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__25523\,
            in1 => \N__40659\,
            in2 => \N__40199\,
            in3 => \N__40437\,
            lcout => \sAddress_RNIA6242_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_3_0_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__25522\,
            in1 => \N__40658\,
            in2 => \N__40439\,
            in3 => \N__40191\,
            lcout => \sAddress_RNIA6242_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI6VH7_4_1_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000010"
        )
    port map (
            in0 => \N__40653\,
            in1 => \N__40545\,
            in2 => \N__40198\,
            in3 => \_gnd_net_\,
            lcout => \sAddress_RNI6VH7_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPoff_10_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47459\,
            lcout => \sEEPoffZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52296\,
            ce => \N__26755\,
            sr => \N__51656\
        );

    \sbuttonModeStatus_RNO_3_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__49095\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35312\,
            lcout => \sbuttonModeStatus_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_0_c_inv_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25592\,
            in2 => \N__30229\,
            in3 => \N__25598\,
            lcout => \sEEDelayACQ_i_0\,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => un4_sacqtime_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_1_c_inv_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25586\,
            in1 => \N__25580\,
            in2 => \N__30109\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQ_i_1\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_0,
            carryout => un4_sacqtime_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_2_c_inv_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25574\,
            in1 => \N__25568\,
            in2 => \N__29996\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQ_i_2\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_1,
            carryout => un4_sacqtime_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_3_c_inv_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29867\,
            in2 => \N__25556\,
            in3 => \N__25562\,
            lcout => \sEEDelayACQ_i_3\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_2,
            carryout => un4_sacqtime_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_4_c_inv_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25541\,
            in2 => \N__31038\,
            in3 => \N__25547\,
            lcout => \sEEDelayACQ_i_4\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_3,
            carryout => un4_sacqtime_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_5_c_inv_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25529\,
            in2 => \N__30900\,
            in3 => \N__25535\,
            lcout => \sEEDelayACQ_i_5\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_4,
            carryout => un4_sacqtime_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_6_c_inv_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25691\,
            in2 => \N__30786\,
            in3 => \N__25697\,
            lcout => \sEEDelayACQ_i_6\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_5,
            carryout => un4_sacqtime_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_7_c_inv_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30651\,
            in2 => \N__25679\,
            in3 => \N__25685\,
            lcout => \sEEDelayACQ_i_7\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_6,
            carryout => un4_sacqtime_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_8_c_inv_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25664\,
            in2 => \N__30562\,
            in3 => \N__25670\,
            lcout => \sEEDelayACQ_i_8\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => un4_sacqtime_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_9_c_inv_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25652\,
            in2 => \N__30456\,
            in3 => \N__25658\,
            lcout => \sEEDelayACQ_i_9\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_8,
            carryout => un4_sacqtime_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_10_c_inv_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25640\,
            in2 => \N__30341\,
            in3 => \N__25646\,
            lcout => \sEEDelayACQ_i_10\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_9,
            carryout => un4_sacqtime_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_11_c_inv_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25628\,
            in2 => \N__33046\,
            in3 => \N__25634\,
            lcout => \sEEDelayACQ_i_11\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_10,
            carryout => un4_sacqtime_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_12_c_inv_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25622\,
            in1 => \N__25616\,
            in2 => \N__31743\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQ_i_12\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_11,
            carryout => un4_sacqtime_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_13_c_inv_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25610\,
            in1 => \N__25604\,
            in2 => \N__31659\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQ_i_13\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_12,
            carryout => un4_sacqtime_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_14_c_inv_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25733\,
            in2 => \N__31574\,
            in3 => \N__25739\,
            lcout => \sEEDelayACQ_i_14\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_13,
            carryout => un4_sacqtime_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_15_c_inv_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25727\,
            in1 => \N__31472\,
            in2 => \N__25721\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQ_i_15\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_14,
            carryout => un4_sacqtime_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_16_c_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31388\,
            in2 => \N__52709\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => un4_sacqtime_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_17_c_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31266\,
            in2 => \N__52707\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_16,
            carryout => un4_sacqtime_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_18_c_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31149\,
            in2 => \N__52710\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_17,
            carryout => un4_sacqtime_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_19_c_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33249\,
            in2 => \N__52708\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_18,
            carryout => un4_sacqtime_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_20_c_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52639\,
            in2 => \N__33381\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_19,
            carryout => un4_sacqtime_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIR3KA_20_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33150\,
            in2 => \N__52705\,
            in3 => \N__33366\,
            lcout => g1_i_a4_4,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_20,
            carryout => un4_sacqtime_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_22_c_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32020\,
            in2 => \N__52711\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_21,
            carryout => un4_sacqtime_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIV7KA_23_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31909\,
            in2 => \N__52706\,
            in3 => \N__32019\,
            lcout => g0_4_0,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_22,
            carryout => un4_sacqtime_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_23_THRU_LUT4_0_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25835\,
            lcout => \un4_sacqtime_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_sclk_inferred_clock_RNO_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48032\,
            in1 => \N__25832\,
            in2 => \_gnd_net_\,
            in3 => \N__25817\,
            lcout => spi_sclk,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_3_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31802\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48444\,
            ce => 'H',
            sr => \N__51750\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_12_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25778\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48444\,
            ce => 'H',
            sr => \N__51750\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_7_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31769\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48444\,
            ce => 'H',
            sr => \N__51750\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_9_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32120\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48444\,
            ce => 'H',
            sr => \N__51750\
        );

    \sDAC_mem_8_0_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46147\,
            lcout => \sDAC_mem_8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52320\,
            ce => \N__27116\,
            sr => \N__51737\
        );

    \sDAC_mem_8_1_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50939\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_8Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52320\,
            ce => \N__27116\,
            sr => \N__51737\
        );

    \sDAC_mem_8_2_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47251\,
            lcout => \sDAC_mem_8Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52320\,
            ce => \N__27116\,
            sr => \N__51737\
        );

    \sDAC_mem_8_3_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46707\,
            lcout => \sDAC_mem_8Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52320\,
            ce => \N__27116\,
            sr => \N__51737\
        );

    \sDAC_mem_8_4_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45397\,
            lcout => \sDAC_mem_8Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52320\,
            ce => \N__27116\,
            sr => \N__51737\
        );

    \sDAC_mem_8_5_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45005\,
            lcout => \sDAC_mem_8Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52320\,
            ce => \N__27116\,
            sr => \N__51737\
        );

    \sDAC_mem_8_6_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50413\,
            lcout => \sDAC_mem_8Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52320\,
            ce => \N__27116\,
            sr => \N__51737\
        );

    \sDAC_mem_8_7_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49893\,
            lcout => \sDAC_mem_8Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52320\,
            ce => \N__27116\,
            sr => \N__51737\
        );

    \sDAC_mem_3_3_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46689\,
            lcout => \sDAC_mem_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52308\,
            ce => \N__44238\,
            sr => \N__51723\
        );

    \sDAC_data_RNO_27_6_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42588\,
            in1 => \N__25991\,
            in2 => \N__42249\,
            in3 => \N__25877\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_6_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42229\,
            in1 => \N__25871\,
            in2 => \N__25859\,
            in3 => \N__25856\,
            lcout => \sDAC_data_RNO_15Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_6_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__25928\,
            in1 => \N__42230\,
            in2 => \N__42595\,
            in3 => \N__26804\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_6_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42231\,
            in1 => \N__39872\,
            in2 => \N__25922\,
            in3 => \N__36815\,
            lcout => \sDAC_data_RNO_7Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_6_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__25919\,
            in1 => \_gnd_net_\,
            in2 => \N__42596\,
            in3 => \N__25910\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_6_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42218\,
            in2 => \N__25901\,
            in3 => \N__25898\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_8Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_6_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011000110010"
        )
    port map (
            in0 => \N__38252\,
            in1 => \N__28859\,
            in2 => \N__25886\,
            in3 => \N__25883\,
            lcout => \sDAC_data_RNO_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_2_0_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46146\,
            lcout => \sDAC_mem_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52297\,
            ce => \N__32851\,
            sr => \N__51713\
        );

    \sDAC_mem_2_1_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50938\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52297\,
            ce => \N__32851\,
            sr => \N__51713\
        );

    \sDAC_mem_2_2_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47245\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52297\,
            ce => \N__32851\,
            sr => \N__51713\
        );

    \sDAC_mem_2_3_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46709\,
            lcout => \sDAC_mem_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52297\,
            ce => \N__32851\,
            sr => \N__51713\
        );

    \sDAC_mem_2_4_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45372\,
            lcout => \sDAC_mem_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52297\,
            ce => \N__32851\,
            sr => \N__51713\
        );

    \sDAC_mem_2_5_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44840\,
            lcout => \sDAC_mem_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52297\,
            ce => \N__32851\,
            sr => \N__51713\
        );

    \sDAC_mem_2_6_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50334\,
            lcout => \sDAC_mem_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52297\,
            ce => \N__32851\,
            sr => \N__51713\
        );

    \sDAC_data_RNO_5_4_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__26249\,
            in1 => \N__25970\,
            in2 => \N__42266\,
            in3 => \N__32564\,
            lcout => \sDAC_data_RNO_5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_7_1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50816\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_7Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52285\,
            ce => \N__44278\,
            sr => \N__51702\
        );

    \sPointer_RNO_2_0_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__44833\,
            in1 => \N__50815\,
            in2 => \N__49994\,
            in3 => \N__46051\,
            lcout => un1_spointer11_2_0_0_a2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_7_0_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46053\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52285\,
            ce => \N__44278\,
            sr => \N__51702\
        );

    \sDAC_mem_7_5_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__44834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_7Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52285\,
            ce => \N__44278\,
            sr => \N__51702\
        );

    \sDAC_mem_7_7_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49892\,
            lcout => \sDAC_mem_7Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52285\,
            ce => \N__44278\,
            sr => \N__51702\
        );

    \sPointer_RNIV9N7_1_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46052\,
            in2 => \_gnd_net_\,
            in3 => \N__26194\,
            lcout => \N_183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPointerReset_RNO_1_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__26195\,
            in1 => \N__26099\,
            in2 => \N__49362\,
            in3 => \N__26048\,
            lcout => \N_1624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_34_0_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46141\,
            lcout => \sDAC_mem_34Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52273\,
            ce => \N__25982\,
            sr => \N__51694\
        );

    \sDAC_mem_34_1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50929\,
            lcout => \sDAC_mem_34Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52273\,
            ce => \N__25982\,
            sr => \N__51694\
        );

    \sDAC_mem_34_2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47246\,
            lcout => \sDAC_mem_34Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52273\,
            ce => \N__25982\,
            sr => \N__51694\
        );

    \sDAC_mem_34_3_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46774\,
            lcout => \sDAC_mem_34Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52273\,
            ce => \N__25982\,
            sr => \N__51694\
        );

    \sDAC_mem_34_4_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45373\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_34Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52273\,
            ce => \N__25982\,
            sr => \N__51694\
        );

    \sDAC_mem_34_5_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44841\,
            lcout => \sDAC_mem_34Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52273\,
            ce => \N__25982\,
            sr => \N__51694\
        );

    \sDAC_mem_34_6_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50481\,
            lcout => \sDAC_mem_34Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52273\,
            ce => \N__25982\,
            sr => \N__51694\
        );

    \sDAC_mem_34_7_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49910\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_34Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52273\,
            ce => \N__25982\,
            sr => \N__51694\
        );

    \sDAC_mem_39_0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46142\,
            lcout => \sDAC_mem_39Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52264\,
            ce => \N__26240\,
            sr => \N__51688\
        );

    \sDAC_mem_39_1_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50930\,
            lcout => \sDAC_mem_39Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52264\,
            ce => \N__26240\,
            sr => \N__51688\
        );

    \sDAC_mem_39_2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47247\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_39Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52264\,
            ce => \N__26240\,
            sr => \N__51688\
        );

    \sDAC_mem_39_3_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46775\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_39Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52264\,
            ce => \N__26240\,
            sr => \N__51688\
        );

    \sDAC_mem_39_4_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45374\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_39Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52264\,
            ce => \N__26240\,
            sr => \N__51688\
        );

    \sDAC_mem_39_5_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45078\,
            lcout => \sDAC_mem_39Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52264\,
            ce => \N__26240\,
            sr => \N__51688\
        );

    \sDAC_mem_39_6_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50482\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_39Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52264\,
            ce => \N__26240\,
            sr => \N__51688\
        );

    \sDAC_mem_39_7_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49911\,
            lcout => \sDAC_mem_39Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52264\,
            ce => \N__26240\,
            sr => \N__51688\
        );

    \un1_spoff_cry_0_c_inv_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27892\,
            in2 => \N__26225\,
            in3 => \N__30188\,
            lcout => \sCounter_i_0\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => un1_spoff_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_1_c_inv_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26210\,
            in2 => \N__27877\,
            in3 => \N__30070\,
            lcout => \sCounter_i_1\,
            ltout => OPEN,
            carryin => un1_spoff_cry_0,
            carryout => un1_spoff_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_2_c_inv_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26339\,
            in2 => \N__27856\,
            in3 => \N__29945\,
            lcout => \sCounter_i_2\,
            ltout => OPEN,
            carryin => un1_spoff_cry_1,
            carryout => un1_spoff_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_3_c_inv_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26327\,
            in2 => \N__28234\,
            in3 => \N__29818\,
            lcout => \sCounter_i_3\,
            ltout => OPEN,
            carryin => un1_spoff_cry_2,
            carryout => un1_spoff_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_4_c_inv_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26315\,
            in2 => \N__28213\,
            in3 => \N__30955\,
            lcout => \sCounter_i_4\,
            ltout => OPEN,
            carryin => un1_spoff_cry_3,
            carryout => un1_spoff_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_5_c_inv_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28189\,
            in2 => \N__26303\,
            in3 => \N__30838\,
            lcout => \sCounter_i_5\,
            ltout => OPEN,
            carryin => un1_spoff_cry_4,
            carryout => un1_spoff_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_6_c_inv_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26288\,
            in2 => \N__28174\,
            in3 => \N__30727\,
            lcout => \sCounter_i_6\,
            ltout => OPEN,
            carryin => un1_spoff_cry_5,
            carryout => un1_spoff_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_7_c_inv_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28150\,
            in2 => \N__26276\,
            in3 => \N__30627\,
            lcout => \sCounter_i_7\,
            ltout => OPEN,
            carryin => un1_spoff_cry_6,
            carryout => un1_spoff_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_8_c_inv_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26780\,
            in2 => \N__28135\,
            in3 => \N__30517\,
            lcout => \sCounter_i_8\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => un1_spoff_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_9_c_inv_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28111\,
            in2 => \N__26768\,
            in3 => \N__30407\,
            lcout => \sCounter_i_9\,
            ltout => OPEN,
            carryin => un1_spoff_cry_8,
            carryout => un1_spoff_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_10_c_inv_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26261\,
            in2 => \N__28096\,
            in3 => \N__30290\,
            lcout => \sCounter_i_10\,
            ltout => OPEN,
            carryin => un1_spoff_cry_9,
            carryout => un1_spoff_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_11_c_inv_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26516\,
            in2 => \N__28357\,
            in3 => \N__32990\,
            lcout => \sCounter_i_11\,
            ltout => OPEN,
            carryin => un1_spoff_cry_10,
            carryout => un1_spoff_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_12_c_inv_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28336\,
            in2 => \N__26504\,
            in3 => \N__31700\,
            lcout => \sCounter_i_12\,
            ltout => OPEN,
            carryin => un1_spoff_cry_11,
            carryout => un1_spoff_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_13_c_inv_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26492\,
            in2 => \N__28318\,
            in3 => \N__31610\,
            lcout => \sCounter_i_13\,
            ltout => OPEN,
            carryin => un1_spoff_cry_12,
            carryout => un1_spoff_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_14_c_inv_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31517\,
            in1 => \N__26480\,
            in2 => \N__28297\,
            in3 => \_gnd_net_\,
            lcout => \sCounter_i_14\,
            ltout => OPEN,
            carryin => un1_spoff_cry_13,
            carryout => un1_spoff_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_15_c_inv_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28273\,
            in2 => \N__26795\,
            in3 => \N__31430\,
            lcout => \sCounter_i_15\,
            ltout => OPEN,
            carryin => un1_spoff_cry_14,
            carryout => un1_spoff_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_16_c_inv_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26357\,
            in2 => \_gnd_net_\,
            in3 => \N__31338\,
            lcout => \sCounter_i_16\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => un1_spoff_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_17_c_inv_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31262\,
            in1 => \N__26351\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sCounter_i_17\,
            ltout => OPEN,
            carryin => un1_spoff_cry_16,
            carryout => un1_spoff_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_18_c_inv_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26345\,
            in2 => \_gnd_net_\,
            in3 => \N__31148\,
            lcout => \sCounter_i_18\,
            ltout => OPEN,
            carryin => un1_spoff_cry_17,
            carryout => un1_spoff_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_19_c_inv_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33225\,
            in1 => \N__26456\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sCounter_i_19\,
            ltout => OPEN,
            carryin => un1_spoff_cry_18,
            carryout => un1_spoff_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_20_c_inv_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26450\,
            in2 => \_gnd_net_\,
            in3 => \N__33332\,
            lcout => \sCounter_i_20\,
            ltout => OPEN,
            carryin => un1_spoff_cry_19,
            carryout => un1_spoff_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_21_c_inv_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33116\,
            in1 => \N__26444\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sCounter_i_21\,
            ltout => OPEN,
            carryin => un1_spoff_cry_20,
            carryout => un1_spoff_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_22_c_inv_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32018\,
            in1 => \N__26438\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sCounter_i_22\,
            ltout => OPEN,
            carryin => un1_spoff_cry_21,
            carryout => un1_spoff_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_23_c_inv_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26432\,
            in2 => \_gnd_net_\,
            in3 => \N__31883\,
            lcout => \sCounter_i_23\,
            ltout => OPEN,
            carryin => un1_spoff_cry_22,
            carryout => un1_spoff_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \poff_obuf_RNO_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__31817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26426\,
            lcout => \N_1683_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__32921\,
            in1 => \N__26363\,
            in2 => \N__26389\,
            in3 => \N__33803\,
            lcout => \sbuttonModeStatusZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_1_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__45752\,
            in1 => \N__45776\,
            in2 => \N__35108\,
            in3 => \N__26372\,
            lcout => \sbuttonModeStatus_0_sqmuxa_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEACQ_0_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46381\,
            lcout => \sEEACQZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52274\,
            ce => \N__26471\,
            sr => \N__51654\
        );

    \sEEACQ_1_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50877\,
            lcout => \sEEACQZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52274\,
            ce => \N__26471\,
            sr => \N__51654\
        );

    \sEEACQ_2_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47458\,
            lcout => \sEEACQZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52274\,
            ce => \N__26471\,
            sr => \N__51654\
        );

    \sEEACQ_3_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46915\,
            lcout => \sEEACQZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52274\,
            ce => \N__26471\,
            sr => \N__51654\
        );

    \sEEACQ_4_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45568\,
            lcout => \sEEACQZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52274\,
            ce => \N__26471\,
            sr => \N__51654\
        );

    \sEEACQ_5_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45080\,
            lcout => \sEEACQZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52274\,
            ce => \N__26471\,
            sr => \N__51654\
        );

    \sEEACQ_6_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50531\,
            lcout => \sEEACQZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52274\,
            ce => \N__26471\,
            sr => \N__51654\
        );

    \sEEACQ_7_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50050\,
            lcout => \sEEACQZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52274\,
            ce => \N__26471\,
            sr => \N__51654\
        );

    \sEEACQ_10_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47460\,
            lcout => \sEEACQZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52286\,
            ce => \N__26525\,
            sr => \N__51651\
        );

    \sEEACQ_11_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46925\,
            lcout => \sEEACQZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52286\,
            ce => \N__26525\,
            sr => \N__51651\
        );

    \sEEACQ_12_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEACQZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52286\,
            ce => \N__26525\,
            sr => \N__51651\
        );

    \sEEACQ_13_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45057\,
            lcout => \sEEACQZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52286\,
            ce => \N__26525\,
            sr => \N__51651\
        );

    \sEEACQ_14_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50544\,
            lcout => \sEEACQZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52286\,
            ce => \N__26525\,
            sr => \N__51651\
        );

    \sEEACQ_15_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50016\,
            lcout => \sEEACQZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52286\,
            ce => \N__26525\,
            sr => \N__51651\
        );

    \sEEACQ_8_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46380\,
            lcout => \sEEACQZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52286\,
            ce => \N__26525\,
            sr => \N__51651\
        );

    \sEEACQ_9_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51018\,
            lcout => \sEEACQZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52286\,
            ce => \N__26525\,
            sr => \N__51651\
        );

    \sEEPoff_11_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46763\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPoffZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52298\,
            ce => \N__26756\,
            sr => \N__51648\
        );

    \sEEPoff_12_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45570\,
            lcout => \sEEPoffZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52298\,
            ce => \N__26756\,
            sr => \N__51648\
        );

    \sEEPoff_13_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45056\,
            lcout => \sEEPoffZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52298\,
            ce => \N__26756\,
            sr => \N__51648\
        );

    \sEEPoff_14_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50545\,
            lcout => \sEEPoffZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52298\,
            ce => \N__26756\,
            sr => \N__51648\
        );

    \sEEPoff_15_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50058\,
            lcout => \sEEPoffZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52298\,
            ce => \N__26756\,
            sr => \N__51648\
        );

    \sEEPoff_8_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46379\,
            lcout => \sEEPoffZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52298\,
            ce => \N__26756\,
            sr => \N__51648\
        );

    \sEEPoff_9_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51062\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPoffZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52298\,
            ce => \N__26756\,
            sr => \N__51648\
        );

    \un4_sacqtime_cry_23_c_RNI2CQM_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__49462\,
            in1 => \N__43315\,
            in2 => \N__39387\,
            in3 => \N__43438\,
            lcout => \un4_sacqtime_cry_23_c_RNI2CQMZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_1_5_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26720\,
            lcout => \RAM_DATA_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52321\,
            ce => \N__51872\,
            sr => \N__51644\
        );

    \RAM_DATA_1_1_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26678\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RAM_DATA_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52321\,
            ce => \N__51872\,
            sr => \N__51644\
        );

    \RAM_DATA_1_10_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26645\,
            lcout => \RAM_DATA_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52321\,
            ce => \N__51872\,
            sr => \N__51644\
        );

    \RAM_DATA_1_11_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26609\,
            lcout => \RAM_DATA_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52321\,
            ce => \N__51872\,
            sr => \N__51644\
        );

    \RAM_DATA_1_13_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26573\,
            lcout => \RAM_DATA_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52321\,
            ce => \N__51872\,
            sr => \N__51644\
        );

    \RAM_DATA_1_14_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26960\,
            lcout => \RAM_DATA_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52321\,
            ce => \N__51872\,
            sr => \N__51644\
        );

    \RAM_DATA_1_2_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26912\,
            lcout => \RAM_DATA_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52321\,
            ce => \N__51872\,
            sr => \N__51644\
        );

    \RAM_DATA_1_6_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26879\,
            lcout => \RAM_DATA_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52339\,
            ce => \N__51889\,
            sr => \N__51642\
        );

    \RAM_DATA_1_0_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26840\,
            lcout => \RAM_DATA_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52339\,
            ce => \N__51889\,
            sr => \N__51642\
        );

    \sDAC_mem_40_0_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46144\,
            lcout => \sDAC_mem_40Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52323\,
            ce => \N__27125\,
            sr => \N__51768\
        );

    \sDAC_mem_40_1_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51075\,
            lcout => \sDAC_mem_40Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52323\,
            ce => \N__27125\,
            sr => \N__51768\
        );

    \sDAC_mem_40_2_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47346\,
            lcout => \sDAC_mem_40Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52323\,
            ce => \N__27125\,
            sr => \N__51768\
        );

    \sDAC_mem_40_3_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46793\,
            lcout => \sDAC_mem_40Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52323\,
            ce => \N__27125\,
            sr => \N__51768\
        );

    \sDAC_mem_40_4_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45529\,
            lcout => \sDAC_mem_40Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52323\,
            ce => \N__27125\,
            sr => \N__51768\
        );

    \sDAC_mem_40_5_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45053\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_40Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52323\,
            ce => \N__27125\,
            sr => \N__51768\
        );

    \sDAC_mem_40_6_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50420\,
            lcout => \sDAC_mem_40Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52323\,
            ce => \N__27125\,
            sr => \N__51768\
        );

    \sDAC_mem_40_7_LC_13_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49995\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_40Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52323\,
            ce => \N__27125\,
            sr => \N__51768\
        );

    \sAddress_RNI9IH12_0_2_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40673\,
            in1 => \N__27020\,
            in2 => \N__41010\,
            in3 => \N__40809\,
            lcout => \sDAC_mem_40_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_3_2_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__40674\,
            in1 => \N__27022\,
            in2 => \N__41011\,
            in3 => \N__40810\,
            lcout => \sDAC_mem_36_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_4_2_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27021\,
            in1 => \N__40811\,
            in2 => \N__41012\,
            in3 => \N__40675\,
            lcout => \sDAC_mem_8_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_rpi_ibuf_RNIRGF52_0_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27110\,
            in1 => \N__27062\,
            in2 => \N__49260\,
            in3 => \N__33769\,
            lcout => \sEEDAC_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_2_2_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__40025\,
            in1 => \_gnd_net_\,
            in2 => \N__40676\,
            in3 => \N__27019\,
            lcout => \sDAC_mem_20_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_1_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26984\,
            in2 => \_gnd_net_\,
            in3 => \N__40024\,
            lcout => \sDAC_mem_21_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_6_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38556\,
            in1 => \N__28478\,
            in2 => \N__38207\,
            in3 => \N__28679\,
            lcout => OPEN,
            ltout => \sDAC_data_2_32_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_6_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__38301\,
            in1 => \N__32354\,
            in2 => \N__27206\,
            in3 => \N__34406\,
            lcout => \sDAC_data_RNO_10Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_6_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38557\,
            in1 => \N__27203\,
            in2 => \N__38208\,
            in3 => \N__36674\,
            lcout => OPEN,
            ltout => \sDAC_data_2_14_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_6_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__38302\,
            in1 => \N__28718\,
            in2 => \N__27197\,
            in3 => \N__39641\,
            lcout => \sDAC_data_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_6_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010101110101"
        )
    port map (
            in0 => \N__37355\,
            in1 => \N__37829\,
            in2 => \N__37472\,
            in3 => \N__27194\,
            lcout => OPEN,
            ltout => \sDAC_data_2_41_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_6_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111000001110"
        )
    port map (
            in0 => \N__37461\,
            in1 => \N__27188\,
            in2 => \N__27182\,
            in3 => \N__27179\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_6_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32099\,
            in1 => \_gnd_net_\,
            in2 => \N__27173\,
            in3 => \N__37636\,
            lcout => \sDAC_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48445\,
            ce => \N__43956\,
            sr => \N__51743\
        );

    \sDAC_mem_3_5_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45001\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52287\,
            ce => \N__44243\,
            sr => \N__51728\
        );

    \sDAC_data_RNO_27_8_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42570\,
            in1 => \N__27161\,
            in2 => \N__42204\,
            in3 => \N__27149\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_8_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42242\,
            in1 => \N__27143\,
            in2 => \N__27134\,
            in3 => \N__27131\,
            lcout => \sDAC_data_RNO_15Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_8_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42569\,
            in1 => \N__27290\,
            in2 => \_gnd_net_\,
            in3 => \N__27278\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_8_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42072\,
            in2 => \N__27266\,
            in3 => \N__27263\,
            lcout => \sDAC_data_RNO_8Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_8_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__27254\,
            in1 => \N__42243\,
            in2 => \N__42580\,
            in3 => \N__27245\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_8_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__36788\,
            in1 => \N__42073\,
            in2 => \N__27236\,
            in3 => \N__39857\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_7Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_8_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010101100100"
        )
    port map (
            in0 => \N__28655\,
            in1 => \N__38303\,
            in2 => \N__27233\,
            in3 => \N__27230\,
            lcout => \sDAC_data_RNO_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_8_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__38476\,
            in1 => \N__27224\,
            in2 => \N__36860\,
            in3 => \N__38288\,
            lcout => OPEN,
            ltout => \sDAC_data_2_14_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_8_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__38289\,
            in1 => \N__32498\,
            in2 => \N__27218\,
            in3 => \N__32549\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_1Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_8_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__37457\,
            in1 => \N__27215\,
            in2 => \N__27209\,
            in3 => \N__27377\,
            lcout => OPEN,
            ltout => \sDAC_data_2_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_8_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__37627\,
            in1 => \N__32087\,
            in2 => \N__27386\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_dataZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48450\,
            ce => \N__43953\,
            sr => \N__51716\
        );

    \sDAC_data_RNO_22_8_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__28565\,
            in1 => \N__38286\,
            in2 => \N__38510\,
            in3 => \N__28814\,
            lcout => OPEN,
            ltout => \sDAC_data_2_32_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_8_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__38287\,
            in1 => \N__32231\,
            in2 => \N__27383\,
            in3 => \N__33581\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_10Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_8_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__37456\,
            in1 => \N__37351\,
            in2 => \N__27380\,
            in3 => \N__27521\,
            lcout => \sDAC_data_2_41_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_3_1_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50928\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52265\,
            ce => \N__44224\,
            sr => \N__51705\
        );

    \sDAC_data_RNO_27_4_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42545\,
            in1 => \N__27371\,
            in2 => \N__42246\,
            in3 => \N__27365\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_4_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__27356\,
            in1 => \N__27350\,
            in2 => \N__27335\,
            in3 => \N__42197\,
            lcout => \sDAC_data_RNO_15Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_4_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27332\,
            in1 => \_gnd_net_\,
            in2 => \N__42574\,
            in3 => \N__27320\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_4_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42198\,
            in2 => \N__27308\,
            in3 => \N__27305\,
            lcout => \sDAC_data_RNO_8Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_4_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42549\,
            in1 => \N__27485\,
            in2 => \N__42247\,
            in3 => \N__27476\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_4_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__36833\,
            in1 => \N__39896\,
            in2 => \N__27464\,
            in3 => \N__42202\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_7Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_4_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010101100100"
        )
    port map (
            in0 => \N__27419\,
            in1 => \N__38111\,
            in2 => \N__27461\,
            in3 => \N__27458\,
            lcout => \sDAC_data_RNO_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_19_3_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27452\,
            in1 => \N__42075\,
            in2 => \_gnd_net_\,
            in3 => \N__27443\,
            lcout => \sDAC_data_RNO_19Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_3_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42076\,
            in1 => \N__45668\,
            in2 => \_gnd_net_\,
            in3 => \N__27584\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_3_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110011101"
        )
    port map (
            in0 => \N__38489\,
            in1 => \N__38290\,
            in2 => \N__27431\,
            in3 => \N__27428\,
            lcout => \sDAC_data_2_24_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_4_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42080\,
            in1 => \N__45653\,
            in2 => \_gnd_net_\,
            in3 => \N__27578\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_4_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110011101"
        )
    port map (
            in0 => \N__38490\,
            in1 => \N__38291\,
            in2 => \N__27422\,
            in3 => \N__27392\,
            lcout => \sDAC_data_2_24_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_19_4_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27413\,
            in1 => \_gnd_net_\,
            in2 => \N__42205\,
            in3 => \N__27404\,
            lcout => \sDAC_data_RNO_19Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_12_0_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46143\,
            lcout => \sDAC_mem_12Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52252\,
            ce => \N__36952\,
            sr => \N__51698\
        );

    \sDAC_mem_12_1_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50931\,
            lcout => \sDAC_mem_12Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52252\,
            ce => \N__36952\,
            sr => \N__51698\
        );

    \sDAC_data_RNO_24_8_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41990\,
            in1 => \N__27572\,
            in2 => \_gnd_net_\,
            in3 => \N__27560\,
            lcout => \sDAC_data_RNO_24Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_8_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42014\,
            in1 => \N__27545\,
            in2 => \_gnd_net_\,
            in3 => \N__27512\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_23Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_8_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__38300\,
            in1 => \N__27530\,
            in2 => \N__27524\,
            in3 => \N__27590\,
            lcout => \sDAC_data_RNO_11Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_28_5_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45077\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_28Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52242\,
            ce => \N__37796\,
            sr => \N__51690\
        );

    \sDAC_data_RNO_30_9_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41989\,
            in1 => \N__41312\,
            in2 => \_gnd_net_\,
            in3 => \N__27506\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_30Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_25_9_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__38249\,
            in1 => \N__38477\,
            in2 => \N__27491\,
            in3 => \N__27695\,
            lcout => OPEN,
            ltout => \sDAC_data_2_39_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_9_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__29423\,
            in1 => \N__38250\,
            in2 => \N__27488\,
            in3 => \N__29636\,
            lcout => \sDAC_data_RNO_11Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_31_9_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42013\,
            in1 => \N__29747\,
            in2 => \_gnd_net_\,
            in3 => \N__27710\,
            lcout => \sDAC_data_RNO_31Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_30_7_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42018\,
            in1 => \N__41339\,
            in2 => \_gnd_net_\,
            in3 => \N__27596\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_30Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_25_7_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__38262\,
            in1 => \N__38425\,
            in2 => \N__27689\,
            in3 => \N__27671\,
            lcout => OPEN,
            ltout => \sDAC_data_2_39_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_7_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__38202\,
            in1 => \N__27602\,
            in2 => \N__27686\,
            in3 => \N__27635\,
            lcout => \sDAC_data_RNO_11Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_31_7_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29768\,
            in1 => \N__42015\,
            in2 => \_gnd_net_\,
            in3 => \N__27683\,
            lcout => \sDAC_data_RNO_31Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_7_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42017\,
            in1 => \N__27665\,
            in2 => \_gnd_net_\,
            in3 => \N__27650\,
            lcout => \sDAC_data_RNO_23Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_7_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27629\,
            in1 => \N__42016\,
            in2 => \_gnd_net_\,
            in3 => \N__27617\,
            lcout => \sDAC_data_RNO_24Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_24_4_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45585\,
            lcout => \sDAC_mem_24Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52233\,
            ce => \N__27741\,
            sr => \N__51683\
        );

    \sDAC_data_RNO_25_8_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38414\,
            in1 => \N__28064\,
            in2 => \N__38285\,
            in3 => \N__29450\,
            lcout => \sDAC_data_2_39_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_31_4_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41607\,
            in1 => \N__29570\,
            in2 => \_gnd_net_\,
            in3 => \N__27836\,
            lcout => \sDAC_data_RNO_31Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_30_4_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42012\,
            in1 => \N__50609\,
            in2 => \_gnd_net_\,
            in3 => \N__27752\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_30Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_25_4_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__38426\,
            in1 => \N__38216\,
            in2 => \N__27824\,
            in3 => \N__27821\,
            lcout => OPEN,
            ltout => \sDAC_data_2_39_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_4_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__38217\,
            in1 => \N__27758\,
            in2 => \N__27815\,
            in3 => \N__27788\,
            lcout => \sDAC_data_RNO_11Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_4_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27812\,
            in1 => \N__42011\,
            in2 => \_gnd_net_\,
            in3 => \N__27800\,
            lcout => \sDAC_data_RNO_23Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_4_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42010\,
            in1 => \N__27782\,
            in2 => \_gnd_net_\,
            in3 => \N__27770\,
            lcout => \sDAC_data_RNO_24Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_24_1_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51017\,
            lcout => \sDAC_mem_24Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52243\,
            ce => \N__27746\,
            sr => \N__51677\
        );

    \sDAC_data_RNO_25_5_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38387\,
            in1 => \N__28076\,
            in2 => \N__38254\,
            in3 => \N__29468\,
            lcout => \sDAC_data_2_39_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_31_5_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41536\,
            in1 => \N__29777\,
            in2 => \_gnd_net_\,
            in3 => \N__28070\,
            lcout => \sDAC_data_RNO_31Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_26_2_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47506\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_26Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52253\,
            ce => \N__28049\,
            sr => \N__51669\
        );

    \sDAC_data_RNO_31_8_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41537\,
            in1 => \N__29756\,
            in2 => \_gnd_net_\,
            in3 => \N__28055\,
            lcout => \sDAC_data_RNO_31Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_26_5_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45079\,
            lcout => \sDAC_mem_26Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52253\,
            ce => \N__28049\,
            sr => \N__51669\
        );

    \spi_master_inst.sclk_gen_u0.delay_clk_i_RNISHDJ_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__27959\,
            in1 => \N__28025\,
            in2 => \_gnd_net_\,
            in3 => \N__28007\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNIK09A_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27958\,
            lcout => \spi_master_inst.sclk_gen_u0.falling_count_start_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_0_c_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27896\,
            in2 => \N__29119\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_14_0_\,
            carryout => un1_sacqtime_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_1_c_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27878\,
            in2 => \N__29086\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_0,
            carryout => un1_sacqtime_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_2_c_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27857\,
            in2 => \N__29050\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_1,
            carryout => un1_sacqtime_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_3_c_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28235\,
            in2 => \N__29023\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_2,
            carryout => un1_sacqtime_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_4_c_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28214\,
            in2 => \N__28996\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_3,
            carryout => un1_sacqtime_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_5_c_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28193\,
            in2 => \N__28960\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_4,
            carryout => un1_sacqtime_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_6_c_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28175\,
            in2 => \N__28930\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_5,
            carryout => un1_sacqtime_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_7_c_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28154\,
            in2 => \N__29377\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_6,
            carryout => un1_sacqtime_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_8_c_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28136\,
            in2 => \N__29341\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => un1_sacqtime_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_9_c_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28115\,
            in2 => \N__29308\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_8,
            carryout => un1_sacqtime_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_10_c_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28097\,
            in2 => \N__29278\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_9,
            carryout => un1_sacqtime_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_11_c_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28358\,
            in2 => \N__29248\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_10,
            carryout => un1_sacqtime_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_12_c_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28337\,
            in2 => \N__29212\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_11,
            carryout => un1_sacqtime_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_13_c_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28319\,
            in2 => \N__29182\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_12,
            carryout => un1_sacqtime_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_14_c_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28298\,
            in2 => \N__29155\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_13,
            carryout => un1_sacqtime_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_15_c_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28277\,
            in2 => \N__29407\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_14,
            carryout => un1_sacqtime_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_16_c_inv_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28259\,
            in2 => \_gnd_net_\,
            in3 => \N__31365\,
            lcout => un1_sacqtime_cry_16_sf,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => un1_sacqtime_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_17_c_inv_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28253\,
            in2 => \_gnd_net_\,
            in3 => \N__31269\,
            lcout => un1_sacqtime_cry_17_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_16,
            carryout => un1_sacqtime_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_18_c_inv_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28247\,
            in2 => \_gnd_net_\,
            in3 => \N__31150\,
            lcout => un1_sacqtime_cry_18_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_17,
            carryout => un1_sacqtime_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_19_c_inv_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33253\,
            in1 => \N__28241\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un1_sacqtime_cry_19_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_18,
            carryout => un1_sacqtime_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_20_c_inv_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28403\,
            in2 => \_gnd_net_\,
            in3 => \N__33373\,
            lcout => un1_sacqtime_cry_20_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_19,
            carryout => un1_sacqtime_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_21_c_inv_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28397\,
            in2 => \_gnd_net_\,
            in3 => \N__33154\,
            lcout => un1_sacqtime_cry_21_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_20,
            carryout => un1_sacqtime_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_22_c_inv_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32027\,
            in1 => \N__28391\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un1_sacqtime_cry_22_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_21,
            carryout => un1_sacqtime_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_23_c_inv_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28385\,
            in2 => \_gnd_net_\,
            in3 => \N__31913\,
            lcout => un1_sacqtime_cry_23_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_22,
            carryout => un1_sacqtime_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_23_THRU_LUT4_0_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28379\,
            lcout => \un1_sacqtime_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sADC_clk_prev_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__34014\,
            in1 => \N__49381\,
            in2 => \N__28376\,
            in3 => \N__48962\,
            lcout => \sADC_clk_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sADC_clk_prev_RNI4BVG_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28372\,
            in2 => \_gnd_net_\,
            in3 => \N__34013\,
            lcout => \N_71\,
            ltout => \N_71_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_23_c_RNIJ7QO_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__49382\,
            in1 => \N__43439\,
            in2 => \N__28364\,
            in3 => \N__43316\,
            lcout => \N_31_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sRAM_pointer_read_0_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39344\,
            in1 => \N__35902\,
            in2 => \_gnd_net_\,
            in3 => \N__28361\,
            lcout => \sRAM_pointer_readZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \sRAM_pointer_read_cry_0\,
            clk => \N__52309\,
            ce => \N__28445\,
            sr => \N__51646\
        );

    \sRAM_pointer_read_1_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39340\,
            in1 => \N__36040\,
            in2 => \_gnd_net_\,
            in3 => \N__28430\,
            lcout => \sRAM_pointer_readZ0Z_1\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_0\,
            carryout => \sRAM_pointer_read_cry_1\,
            clk => \N__52309\,
            ce => \N__28445\,
            sr => \N__51646\
        );

    \sRAM_pointer_read_2_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39345\,
            in1 => \N__36130\,
            in2 => \_gnd_net_\,
            in3 => \N__28427\,
            lcout => \sRAM_pointer_readZ0Z_2\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_1\,
            carryout => \sRAM_pointer_read_cry_2\,
            clk => \N__52309\,
            ce => \N__28445\,
            sr => \N__51646\
        );

    \sRAM_pointer_read_3_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39341\,
            in1 => \N__43366\,
            in2 => \_gnd_net_\,
            in3 => \N__28424\,
            lcout => \sRAM_pointer_readZ0Z_3\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_2\,
            carryout => \sRAM_pointer_read_cry_3\,
            clk => \N__52309\,
            ce => \N__28445\,
            sr => \N__51646\
        );

    \sRAM_pointer_read_4_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39346\,
            in1 => \N__43549\,
            in2 => \_gnd_net_\,
            in3 => \N__28421\,
            lcout => \sRAM_pointer_readZ0Z_4\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_3\,
            carryout => \sRAM_pointer_read_cry_4\,
            clk => \N__52309\,
            ce => \N__28445\,
            sr => \N__51646\
        );

    \sRAM_pointer_read_5_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39342\,
            in1 => \N__35248\,
            in2 => \_gnd_net_\,
            in3 => \N__28418\,
            lcout => \sRAM_pointer_readZ0Z_5\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_4\,
            carryout => \sRAM_pointer_read_cry_5\,
            clk => \N__52309\,
            ce => \N__28445\,
            sr => \N__51646\
        );

    \sRAM_pointer_read_6_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39347\,
            in1 => \N__35983\,
            in2 => \_gnd_net_\,
            in3 => \N__28415\,
            lcout => \sRAM_pointer_readZ0Z_6\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_5\,
            carryout => \sRAM_pointer_read_cry_6\,
            clk => \N__52309\,
            ce => \N__28445\,
            sr => \N__51646\
        );

    \sRAM_pointer_read_7_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39343\,
            in1 => \N__36163\,
            in2 => \_gnd_net_\,
            in3 => \N__28412\,
            lcout => \sRAM_pointer_readZ0Z_7\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_6\,
            carryout => \sRAM_pointer_read_cry_7\,
            clk => \N__52309\,
            ce => \N__28445\,
            sr => \N__51646\
        );

    \sRAM_pointer_read_8_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39395\,
            in1 => \N__43621\,
            in2 => \_gnd_net_\,
            in3 => \N__28409\,
            lcout => \sRAM_pointer_readZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \sRAM_pointer_read_cry_8\,
            clk => \N__52322\,
            ce => \N__28444\,
            sr => \N__51645\
        );

    \sRAM_pointer_read_9_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39391\,
            in1 => \N__36229\,
            in2 => \_gnd_net_\,
            in3 => \N__28406\,
            lcout => \sRAM_pointer_readZ0Z_9\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_8\,
            carryout => \sRAM_pointer_read_cry_9\,
            clk => \N__52322\,
            ce => \N__28444\,
            sr => \N__51645\
        );

    \sRAM_pointer_read_10_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39392\,
            in1 => \N__35839\,
            in2 => \_gnd_net_\,
            in3 => \N__28472\,
            lcout => \sRAM_pointer_readZ0Z_10\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_9\,
            carryout => \sRAM_pointer_read_cry_10\,
            clk => \N__52322\,
            ce => \N__28444\,
            sr => \N__51645\
        );

    \sRAM_pointer_read_11_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39388\,
            in1 => \N__35767\,
            in2 => \_gnd_net_\,
            in3 => \N__28469\,
            lcout => \sRAM_pointer_readZ0Z_11\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_10\,
            carryout => \sRAM_pointer_read_cry_11\,
            clk => \N__52322\,
            ce => \N__28444\,
            sr => \N__51645\
        );

    \sRAM_pointer_read_12_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39393\,
            in1 => \N__35671\,
            in2 => \_gnd_net_\,
            in3 => \N__28466\,
            lcout => \sRAM_pointer_readZ0Z_12\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_11\,
            carryout => \sRAM_pointer_read_cry_12\,
            clk => \N__52322\,
            ce => \N__28444\,
            sr => \N__51645\
        );

    \sRAM_pointer_read_13_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39389\,
            in1 => \N__35632\,
            in2 => \_gnd_net_\,
            in3 => \N__28463\,
            lcout => \sRAM_pointer_readZ0Z_13\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_12\,
            carryout => \sRAM_pointer_read_cry_13\,
            clk => \N__52322\,
            ce => \N__28444\,
            sr => \N__51645\
        );

    \sRAM_pointer_read_14_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39394\,
            in1 => \N__35539\,
            in2 => \_gnd_net_\,
            in3 => \N__28460\,
            lcout => \sRAM_pointer_readZ0Z_14\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_13\,
            carryout => \sRAM_pointer_read_cry_14\,
            clk => \N__52322\,
            ce => \N__28444\,
            sr => \N__51645\
        );

    \sRAM_pointer_read_15_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39390\,
            in1 => \N__35497\,
            in2 => \_gnd_net_\,
            in3 => \N__28457\,
            lcout => \sRAM_pointer_readZ0Z_15\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_14\,
            carryout => \sRAM_pointer_read_cry_15\,
            clk => \N__52322\,
            ce => \N__28444\,
            sr => \N__51645\
        );

    \sRAM_pointer_read_16_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39296\,
            in1 => \N__35425\,
            in2 => \_gnd_net_\,
            in3 => \N__28454\,
            lcout => \sRAM_pointer_readZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \sRAM_pointer_read_cry_16\,
            clk => \N__52330\,
            ce => \N__28443\,
            sr => \N__51643\
        );

    \sRAM_pointer_read_17_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39295\,
            in1 => \N__36367\,
            in2 => \_gnd_net_\,
            in3 => \N__28451\,
            lcout => \sRAM_pointer_readZ0Z_17\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_16\,
            carryout => \sRAM_pointer_read_cry_17\,
            clk => \N__52330\,
            ce => \N__28443\,
            sr => \N__51643\
        );

    \sRAM_pointer_read_18_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39297\,
            in1 => \N__36301\,
            in2 => \_gnd_net_\,
            in3 => \N__28448\,
            lcout => \sRAM_pointer_readZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52330\,
            ce => \N__28443\,
            sr => \N__51643\
        );

    \sDAC_mem_36_0_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46145\,
            lcout => \sDAC_mem_36Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52310\,
            ce => \N__28484\,
            sr => \N__51782\
        );

    \sDAC_mem_36_1_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51074\,
            lcout => \sDAC_mem_36Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52310\,
            ce => \N__28484\,
            sr => \N__51782\
        );

    \sDAC_mem_36_2_LC_14_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47328\,
            lcout => \sDAC_mem_36Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52310\,
            ce => \N__28484\,
            sr => \N__51782\
        );

    \sDAC_mem_36_3_LC_14_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46901\,
            lcout => \sDAC_mem_36Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52310\,
            ce => \N__28484\,
            sr => \N__51782\
        );

    \sDAC_mem_36_4_LC_14_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45530\,
            lcout => \sDAC_mem_36Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52310\,
            ce => \N__28484\,
            sr => \N__51782\
        );

    \sDAC_mem_36_5_LC_14_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45055\,
            lcout => \sDAC_mem_36Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52310\,
            ce => \N__28484\,
            sr => \N__51782\
        );

    \sDAC_mem_36_6_LC_14_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50408\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_36Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52310\,
            ce => \N__28484\,
            sr => \N__51782\
        );

    \sDAC_mem_36_7_LC_14_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49996\,
            lcout => \sDAC_mem_36Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52310\,
            ce => \N__28484\,
            sr => \N__51782\
        );

    \sDAC_data_RNO_29_6_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41813\,
            in1 => \N__35012\,
            in2 => \_gnd_net_\,
            in3 => \N__28577\,
            lcout => \sDAC_data_RNO_29Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_18_3_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46746\,
            lcout => \sDAC_mem_18Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52300\,
            ce => \N__28544\,
            sr => \N__51769\
        );

    \sDAC_data_RNO_29_7_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41810\,
            in1 => \N__33923\,
            in2 => \_gnd_net_\,
            in3 => \N__28571\,
            lcout => \sDAC_data_RNO_29Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_18_4_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45528\,
            lcout => \sDAC_mem_18Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52300\,
            ce => \N__28544\,
            sr => \N__51769\
        );

    \sDAC_data_RNO_29_8_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41811\,
            in1 => \N__33911\,
            in2 => \_gnd_net_\,
            in3 => \N__28556\,
            lcout => \sDAC_data_RNO_29Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_18_5_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45054\,
            lcout => \sDAC_mem_18Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52300\,
            ce => \N__28544\,
            sr => \N__51769\
        );

    \sDAC_data_RNO_29_9_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41812\,
            in1 => \N__34091\,
            in2 => \_gnd_net_\,
            in3 => \N__28550\,
            lcout => \sDAC_data_RNO_29Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_18_6_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50407\,
            lcout => \sDAC_mem_18Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52300\,
            ce => \N__28544\,
            sr => \N__51769\
        );

    \sDAC_data_RNO_19_7_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42093\,
            in1 => \N__28517\,
            in2 => \_gnd_net_\,
            in3 => \N__28505\,
            lcout => \sDAC_data_RNO_19Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_7_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42233\,
            in1 => \N__45134\,
            in2 => \_gnd_net_\,
            in3 => \N__28619\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_7_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__38129\,
            in1 => \N__38553\,
            in2 => \N__28493\,
            in3 => \N__28490\,
            lcout => \sDAC_data_2_24_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_8_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42234\,
            in1 => \N__44624\,
            in2 => \_gnd_net_\,
            in3 => \N__28613\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_8_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__38130\,
            in1 => \N__38554\,
            in2 => \N__28658\,
            in3 => \N__28625\,
            lcout => \sDAC_data_2_24_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_19_8_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42232\,
            in1 => \N__28649\,
            in2 => \_gnd_net_\,
            in3 => \N__28637\,
            lcout => \sDAC_data_RNO_19Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_12_4_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45348\,
            lcout => \sDAC_mem_12Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52288\,
            ce => \N__36960\,
            sr => \N__51756\
        );

    \sDAC_mem_12_5_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__44867\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_12Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52288\,
            ce => \N__36960\,
            sr => \N__51756\
        );

    \sDAC_data_RNO_13_5_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110111"
        )
    port map (
            in0 => \N__28607\,
            in1 => \N__42567\,
            in2 => \N__42192\,
            in3 => \N__28583\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_5_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42067\,
            in1 => \N__28598\,
            in2 => \N__28586\,
            in3 => \N__43835\,
            lcout => \sDAC_data_RNO_5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_6_2_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47364\,
            lcout => \sDAC_mem_6Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52275\,
            ce => \N__36549\,
            sr => \N__51744\
        );

    \sDAC_data_RNO_13_6_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42568\,
            in1 => \N__28745\,
            in2 => \N__42203\,
            in3 => \N__28712\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_6_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42052\,
            in1 => \N__28733\,
            in2 => \N__28721\,
            in3 => \N__43820\,
            lcout => \sDAC_data_RNO_5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_6_3_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46794\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_6Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52275\,
            ce => \N__36549\,
            sr => \N__51744\
        );

    \sDAC_data_RNO_13_7_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42559\,
            in1 => \N__28706\,
            in2 => \N__42193\,
            in3 => \N__36581\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_7_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42068\,
            in1 => \N__28697\,
            in2 => \N__28682\,
            in3 => \N__44312\,
            lcout => \sDAC_data_RNO_5Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_28_6_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41873\,
            in1 => \N__38612\,
            in2 => \_gnd_net_\,
            in3 => \N__28670\,
            lcout => \sDAC_data_RNO_28Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_16_3_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46891\,
            lcout => \sDAC_mem_16Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52266\,
            ce => \N__33508\,
            sr => \N__51729\
        );

    \sDAC_data_RNO_28_7_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41872\,
            in1 => \N__39008\,
            in2 => \_gnd_net_\,
            in3 => \N__28664\,
            lcout => \sDAC_data_RNO_28Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_16_4_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45531\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_16Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52266\,
            ce => \N__33508\,
            sr => \N__51729\
        );

    \sDAC_data_RNO_28_8_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41874\,
            in1 => \N__38993\,
            in2 => \_gnd_net_\,
            in3 => \N__28808\,
            lcout => \sDAC_data_RNO_28Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_16_5_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45081\,
            lcout => \sDAC_mem_16Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52266\,
            ce => \N__33508\,
            sr => \N__51729\
        );

    \sDAC_data_RNO_28_9_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41875\,
            in1 => \N__38978\,
            in2 => \_gnd_net_\,
            in3 => \N__28802\,
            lcout => \sDAC_data_RNO_28Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_16_6_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50468\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_16Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52266\,
            ce => \N__33508\,
            sr => \N__51729\
        );

    \sDAC_data_RNO_10_4_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__34436\,
            in1 => \N__32384\,
            in2 => \N__38210\,
            in3 => \N__28898\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_10Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_4_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__37439\,
            in1 => \N__37344\,
            in2 => \N__28796\,
            in3 => \N__28793\,
            lcout => \sDAC_data_2_41_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_4_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__41144\,
            in1 => \N__28781\,
            in2 => \N__38211\,
            in3 => \N__28904\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_4_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__37440\,
            in1 => \N__28769\,
            in2 => \N__28763\,
            in3 => \N__28760\,
            lcout => OPEN,
            ltout => \sDAC_data_2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_4_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__37628\,
            in1 => \N__32111\,
            in2 => \N__28754\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48457\,
            ce => \N__43950\,
            sr => \N__51717\
        );

    \sDAC_data_RNO_6_4_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38558\,
            in1 => \N__28751\,
            in2 => \N__38212\,
            in3 => \N__41045\,
            lcout => \sDAC_data_2_14_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_4_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38555\,
            in1 => \N__34787\,
            in2 => \N__38209\,
            in3 => \N__29594\,
            lcout => \sDAC_data_2_32_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_19_5_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42082\,
            in1 => \N__28892\,
            in2 => \_gnd_net_\,
            in3 => \N__28883\,
            lcout => \sDAC_data_RNO_19Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_5_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41809\,
            in1 => \N__45638\,
            in2 => \_gnd_net_\,
            in3 => \N__28820\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_5_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__38168\,
            in1 => \N__38551\,
            in2 => \N__28871\,
            in3 => \N__28868\,
            lcout => \sDAC_data_2_24_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_6_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41808\,
            in1 => \N__45623\,
            in2 => \_gnd_net_\,
            in3 => \N__29126\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_6_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__38169\,
            in1 => \N__38550\,
            in2 => \N__28862\,
            in3 => \N__28826\,
            lcout => \sDAC_data_2_24_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_19_6_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28847\,
            in1 => \N__42081\,
            in2 => \_gnd_net_\,
            in3 => \N__28838\,
            lcout => \sDAC_data_RNO_19Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_12_2_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47345\,
            lcout => \sDAC_mem_12Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52244\,
            ce => \N__36965\,
            sr => \N__51706\
        );

    \sDAC_mem_12_3_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46853\,
            lcout => \sDAC_mem_12Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52244\,
            ce => \N__36965\,
            sr => \N__51706\
        );

    \un5_sdacdyn_cry_0_c_inv_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30216\,
            in2 => \N__29096\,
            in3 => \N__29120\,
            lcout => \sEEACQ_i_0\,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => un5_sdacdyn_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_1_c_inv_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30096\,
            in2 => \N__29063\,
            in3 => \N__29087\,
            lcout => \sEEACQ_i_1\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_0,
            carryout => un5_sdacdyn_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_2_c_inv_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29033\,
            in2 => \N__29997\,
            in3 => \N__29054\,
            lcout => \sEEACQ_i_2\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_1,
            carryout => un5_sdacdyn_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_3_c_inv_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29871\,
            in2 => \N__29006\,
            in3 => \N__29027\,
            lcout => \sEEACQ_i_3\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_2,
            carryout => un5_sdacdyn_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_4_c_inv_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31001\,
            in2 => \N__28973\,
            in3 => \N__28997\,
            lcout => \sEEACQ_i_4\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_3,
            carryout => un5_sdacdyn_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_5_c_inv_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30881\,
            in2 => \N__28943\,
            in3 => \N__28964\,
            lcout => \sEEACQ_i_5\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_4,
            carryout => un5_sdacdyn_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_6_c_inv_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28934\,
            in1 => \N__30762\,
            in2 => \N__28913\,
            in3 => \_gnd_net_\,
            lcout => \sEEACQ_i_6\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_5,
            carryout => un5_sdacdyn_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_7_c_inv_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29378\,
            in1 => \N__30652\,
            in2 => \N__29354\,
            in3 => \_gnd_net_\,
            lcout => \sEEACQ_i_7\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_6,
            carryout => un5_sdacdyn_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_8_c_inv_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30551\,
            in2 => \N__29324\,
            in3 => \N__29345\,
            lcout => \sEEACQ_i_8\,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => un5_sdacdyn_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_9_c_inv_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30445\,
            in2 => \N__29291\,
            in3 => \N__29315\,
            lcout => \sEEACQ_i_9\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_8,
            carryout => un5_sdacdyn_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_10_c_inv_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30337\,
            in2 => \N__29258\,
            in3 => \N__29282\,
            lcout => \sEEACQ_i_10\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_9,
            carryout => un5_sdacdyn_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_11_c_inv_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33052\,
            in2 => \N__29225\,
            in3 => \N__29249\,
            lcout => \sEEACQ_i_11\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_10,
            carryout => un5_sdacdyn_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_12_c_inv_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31732\,
            in2 => \N__29195\,
            in3 => \N__29216\,
            lcout => \sEEACQ_i_12\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_11,
            carryout => un5_sdacdyn_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_13_c_inv_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31644\,
            in2 => \N__29165\,
            in3 => \N__29186\,
            lcout => \sEEACQ_i_13\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_12,
            carryout => un5_sdacdyn_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_14_c_inv_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29132\,
            in2 => \N__31579\,
            in3 => \N__29156\,
            lcout => \sEEACQ_i_14\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_13,
            carryout => un5_sdacdyn_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_15_c_inv_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31454\,
            in2 => \N__29390\,
            in3 => \N__29411\,
            lcout => \sEEACQ_i_15\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_14,
            carryout => un5_sdacdyn_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_16_c_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31389\,
            in2 => \N__52570\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => un5_sdacdyn_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_17_c_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52491\,
            in2 => \N__31284\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_16,
            carryout => un5_sdacdyn_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_18_c_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31162\,
            in2 => \N__52571\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_17,
            carryout => un5_sdacdyn_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_19_c_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52495\,
            in2 => \N__33274\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_18,
            carryout => un5_sdacdyn_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_20_c_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33375\,
            in2 => \N__52572\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_19,
            carryout => un5_sdacdyn_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_21_c_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52499\,
            in2 => \N__33169\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_20,
            carryout => un5_sdacdyn_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_22_c_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32037\,
            in2 => \N__52573\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_21,
            carryout => un5_sdacdyn_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_23_c_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52503\,
            in2 => \N__31936\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_22,
            carryout => un5_sdacdyn_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_23_c_RNIELG28_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__29557\,
            in1 => \N__36899\,
            in2 => \N__31052\,
            in3 => \N__29528\,
            lcout => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_pointer_0_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41566\,
            in2 => \_gnd_net_\,
            in3 => \N__37584\,
            lcout => \sDAC_mem_pointerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48469\,
            ce => \N__43951\,
            sr => \N__51678\
        );

    \sDAC_data_RNO_30_10_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41565\,
            in1 => \N__42803\,
            in2 => \_gnd_net_\,
            in3 => \N__29525\,
            lcout => \sDAC_data_RNO_30Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_31_10_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29735\,
            in1 => \N__41564\,
            in2 => \_gnd_net_\,
            in3 => \N__29513\,
            lcout => \sDAC_data_RNO_31Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_pointer_1_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__37582\,
            in1 => \N__38403\,
            in2 => \_gnd_net_\,
            in3 => \N__41658\,
            lcout => \sDAC_mem_pointerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48469\,
            ce => \N__43951\,
            sr => \N__51678\
        );

    \sDAC_data_10_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32072\,
            in1 => \N__37583\,
            in2 => \_gnd_net_\,
            in3 => \N__32927\,
            lcout => \sDAC_dataZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48469\,
            ce => \N__43951\,
            sr => \N__51678\
        );

    \sDAC_data_RNO_30_5_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41563\,
            in1 => \N__41357\,
            in2 => \_gnd_net_\,
            in3 => \N__29480\,
            lcout => \sDAC_data_RNO_30Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_30_8_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41657\,
            in1 => \N__41369\,
            in2 => \_gnd_net_\,
            in3 => \N__29462\,
            lcout => \sDAC_data_RNO_30Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_9_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41861\,
            in1 => \N__29438\,
            in2 => \_gnd_net_\,
            in3 => \N__29714\,
            lcout => \sDAC_data_RNO_23Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_28_6_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50546\,
            lcout => \sDAC_mem_28Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52254\,
            ce => \N__37807\,
            sr => \N__51670\
        );

    \sDAC_data_RNO_24_3_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41864\,
            in1 => \N__29708\,
            in2 => \_gnd_net_\,
            in3 => \N__29699\,
            lcout => \sDAC_data_RNO_24Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_6_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41720\,
            in1 => \N__29684\,
            in2 => \_gnd_net_\,
            in3 => \N__29675\,
            lcout => \sDAC_data_RNO_24Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_9_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41862\,
            in1 => \N__29663\,
            in2 => \_gnd_net_\,
            in3 => \N__29651\,
            lcout => \sDAC_data_RNO_24Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_28_3_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41721\,
            in1 => \N__38639\,
            in2 => \_gnd_net_\,
            in3 => \N__29624\,
            lcout => \sDAC_data_RNO_28Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_28_4_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41863\,
            in1 => \N__38630\,
            in2 => \_gnd_net_\,
            in3 => \N__29609\,
            lcout => \sDAC_data_RNO_28Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_28_5_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41722\,
            in1 => \N__38621\,
            in2 => \_gnd_net_\,
            in3 => \N__29582\,
            lcout => \sDAC_data_RNO_28Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_27_0_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46235\,
            lcout => \sDAC_mem_27Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52267\,
            ce => \N__29726\,
            sr => \N__51663\
        );

    \sDAC_mem_27_1_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51041\,
            lcout => \sDAC_mem_27Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52267\,
            ce => \N__29726\,
            sr => \N__51663\
        );

    \sDAC_mem_27_2_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47343\,
            lcout => \sDAC_mem_27Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52267\,
            ce => \N__29726\,
            sr => \N__51663\
        );

    \sDAC_mem_27_3_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46905\,
            lcout => \sDAC_mem_27Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52267\,
            ce => \N__29726\,
            sr => \N__51663\
        );

    \sDAC_mem_27_4_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45605\,
            lcout => \sDAC_mem_27Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52267\,
            ce => \N__29726\,
            sr => \N__51663\
        );

    \sDAC_mem_27_5_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45119\,
            lcout => \sDAC_mem_27Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52267\,
            ce => \N__29726\,
            sr => \N__51663\
        );

    \sDAC_mem_27_6_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50541\,
            lcout => \sDAC_mem_27Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52267\,
            ce => \N__29726\,
            sr => \N__51663\
        );

    \sDAC_mem_27_7_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50059\,
            lcout => \sDAC_mem_27Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52267\,
            ce => \N__29726\,
            sr => \N__51663\
        );

    \sEEPonPoff_0_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46234\,
            lcout => \sEEPonPoffZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52276\,
            ce => \N__33677\,
            sr => \N__51657\
        );

    \sEEPonPoff_1_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51040\,
            lcout => \sEEPonPoffZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52276\,
            ce => \N__33677\,
            sr => \N__51657\
        );

    \sEEPonPoff_2_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47344\,
            lcout => \sEEPonPoffZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52276\,
            ce => \N__33677\,
            sr => \N__51657\
        );

    \sEEPonPoff_3_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46764\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoffZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52276\,
            ce => \N__33677\,
            sr => \N__51657\
        );

    \sEEPonPoff_4_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45606\,
            lcout => \sEEPonPoffZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52276\,
            ce => \N__33677\,
            sr => \N__51657\
        );

    \sEEPonPoff_5_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45114\,
            lcout => \sEEPonPoffZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52276\,
            ce => \N__33677\,
            sr => \N__51657\
        );

    \sEEPonPoff_6_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50543\,
            lcout => \sEEPonPoffZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52276\,
            ce => \N__33677\,
            sr => \N__51657\
        );

    \sEEPonPoff_7_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50047\,
            lcout => \sEEPonPoffZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52276\,
            ce => \N__33677\,
            sr => \N__51657\
        );

    \un4_spoff_cry_0_c_inv_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30248\,
            in1 => \N__30143\,
            in2 => \N__30242\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoff_i_0\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => un4_spoff_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_1_c_inv_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30026\,
            in2 => \N__30137\,
            in3 => \N__30032\,
            lcout => \sEEPonPoff_i_1\,
            ltout => OPEN,
            carryin => un4_spoff_cry_0,
            carryout => un4_spoff_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_2_c_inv_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30020\,
            in1 => \N__29897\,
            in2 => \N__30014\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoff_i_2\,
            ltout => OPEN,
            carryin => un4_spoff_cry_1,
            carryout => un4_spoff_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_3_c_inv_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29891\,
            in1 => \N__29783\,
            in2 => \N__29884\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoff_i_3\,
            ltout => OPEN,
            carryin => un4_spoff_cry_2,
            carryout => un4_spoff_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_4_c_inv_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31067\,
            in1 => \N__30920\,
            in2 => \N__31060\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoff_i_4\,
            ltout => OPEN,
            carryin => un4_spoff_cry_3,
            carryout => un4_spoff_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_5_c_inv_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30914\,
            in1 => \N__30803\,
            in2 => \N__30908\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoff_i_5\,
            ltout => OPEN,
            carryin => un4_spoff_cry_4,
            carryout => un4_spoff_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_6_c_inv_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30797\,
            in1 => \N__30692\,
            in2 => \N__30791\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoff_i_6\,
            ltout => OPEN,
            carryin => un4_spoff_cry_5,
            carryout => un4_spoff_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_7_c_inv_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30581\,
            in2 => \N__30686\,
            in3 => \N__30587\,
            lcout => \sEEPonPoff_i_7\,
            ltout => OPEN,
            carryin => un4_spoff_cry_6,
            carryout => un4_spoff_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_8_c_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30571\,
            in2 => \N__52671\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => un4_spoff_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_9_c_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52602\,
            in2 => \N__30470\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_8,
            carryout => un4_spoff_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_10_c_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30360\,
            in2 => \N__52668\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_9,
            carryout => un4_spoff_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_11_c_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52590\,
            in2 => \N__33062\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_10,
            carryout => un4_spoff_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_12_c_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31747\,
            in2 => \N__52669\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_11,
            carryout => un4_spoff_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_13_c_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52594\,
            in2 => \N__31664\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_12,
            carryout => un4_spoff_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_14_c_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31578\,
            in2 => \N__52670\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_13,
            carryout => un4_spoff_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_15_c_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52598\,
            in2 => \N__31484\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_14,
            carryout => un4_spoff_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_16_c_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52536\,
            in2 => \N__31397\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => un4_spoff_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_17_c_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31283\,
            in2 => \N__52623\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_16,
            carryout => un4_spoff_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_18_c_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52540\,
            in2 => \N__31176\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_17,
            carryout => un4_spoff_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_19_c_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33273\,
            in2 => \N__52624\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_18,
            carryout => un4_spoff_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_20_c_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52544\,
            in2 => \N__33388\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_19,
            carryout => un4_spoff_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_21_c_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33167\,
            in2 => \N__52625\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_20,
            carryout => un4_spoff_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_22_c_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52548\,
            in2 => \N__32048\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_21,
            carryout => un4_spoff_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_23_c_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31929\,
            in2 => \N__52626\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_22,
            carryout => un4_spoff_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_23_THRU_LUT4_0_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31820\,
            lcout => \un4_spoff_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.data_in_3_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37526\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48446\,
            ce => \N__43903\,
            sr => \N__51796\
        );

    \spi_master_inst.spi_data_path_u1.data_in_4_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31793\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48446\,
            ce => \N__43903\,
            sr => \N__51796\
        );

    \spi_master_inst.spi_data_path_u1.data_in_7_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32132\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48446\,
            ce => \N__43903\,
            sr => \N__51796\
        );

    \spi_master_inst.spi_data_path_u1.data_in_8_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31760\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48446\,
            ce => \N__43903\,
            sr => \N__51796\
        );

    \spi_master_inst.spi_data_path_u1.data_in_9_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32288\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48446\,
            ce => \N__43903\,
            sr => \N__51796\
        );

    \sEEDAC_0_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46233\,
            lcout => \sEEDACZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52289\,
            ce => \N__32057\,
            sr => \_gnd_net_\
        );

    \sEEDAC_1_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50982\,
            lcout => \sEEDACZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52289\,
            ce => \N__32057\,
            sr => \_gnd_net_\
        );

    \sEEDAC_2_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47347\,
            lcout => \sEEDACZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52289\,
            ce => \N__32057\,
            sr => \_gnd_net_\
        );

    \sEEDAC_3_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46750\,
            lcout => \sEEDACZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52289\,
            ce => \N__32057\,
            sr => \_gnd_net_\
        );

    \sEEDAC_4_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45506\,
            lcout => \sEEDACZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52289\,
            ce => \N__32057\,
            sr => \_gnd_net_\
        );

    \sEEDAC_5_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44980\,
            lcout => \sEEDACZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52289\,
            ce => \N__32057\,
            sr => \_gnd_net_\
        );

    \sEEDAC_6_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50409\,
            lcout => \sEEDACZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52289\,
            ce => \N__32057\,
            sr => \_gnd_net_\
        );

    \sEEDAC_7_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50052\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEDACZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52289\,
            ce => \N__32057\,
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_7_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__34385\,
            in1 => \N__33602\,
            in2 => \N__38258\,
            in3 => \N__32189\,
            lcout => \sDAC_data_RNO_10Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_7_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38508\,
            in1 => \N__32204\,
            in2 => \N__38200\,
            in3 => \N__32198\,
            lcout => \sDAC_data_2_32_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_7_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38509\,
            in1 => \N__34187\,
            in2 => \N__38257\,
            in3 => \N__36881\,
            lcout => OPEN,
            ltout => \sDAC_data_2_14_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_7_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__32327\,
            in1 => \N__38230\,
            in2 => \N__32183\,
            in3 => \N__32180\,
            lcout => \sDAC_data_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_7_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010101110101"
        )
    port map (
            in0 => \N__37342\,
            in1 => \N__32174\,
            in2 => \N__37487\,
            in3 => \N__32159\,
            lcout => OPEN,
            ltout => \sDAC_data_2_41_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_7_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111000001110"
        )
    port map (
            in0 => \N__34142\,
            in1 => \N__37485\,
            in2 => \N__32153\,
            in3 => \N__32150\,
            lcout => OPEN,
            ltout => \sDAC_data_2_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_7_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32144\,
            in1 => \_gnd_net_\,
            in2 => \N__32135\,
            in3 => \N__37637\,
            lcout => \sDAC_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48453\,
            ce => \N__43954\,
            sr => \N__51770\
        );

    \sDAC_data_RNO_1_9_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__32453\,
            in1 => \N__32684\,
            in2 => \N__38256\,
            in3 => \N__32279\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_9_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__37486\,
            in1 => \N__34253\,
            in2 => \N__32123\,
            in3 => \N__32237\,
            lcout => OPEN,
            ltout => \sDAC_data_2_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_9_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32300\,
            in1 => \_gnd_net_\,
            in2 => \N__32291\,
            in3 => \N__37630\,
            lcout => \sDAC_dataZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48456\,
            ce => \N__43952\,
            sr => \N__51757\
        );

    \sDAC_data_RNO_6_9_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110111"
        )
    port map (
            in0 => \N__34337\,
            in1 => \N__38533\,
            in2 => \N__38201\,
            in3 => \N__34460\,
            lcout => \sDAC_data_2_14_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_9_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38532\,
            in1 => \N__32273\,
            in2 => \N__38255\,
            in3 => \N__32264\,
            lcout => OPEN,
            ltout => \sDAC_data_2_32_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_9_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__38104\,
            in1 => \N__33560\,
            in2 => \N__32258\,
            in3 => \N__32216\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_10Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_9_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__37462\,
            in1 => \N__37341\,
            in2 => \N__32255\,
            in3 => \N__32252\,
            lcout => \sDAC_data_2_41_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_20_8_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34067\,
            in1 => \N__42146\,
            in2 => \_gnd_net_\,
            in3 => \N__32222\,
            lcout => \sDAC_data_RNO_20Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_20_5_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45068\,
            lcout => \sDAC_mem_20Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52255\,
            ce => \N__36637\,
            sr => \N__51745\
        );

    \sDAC_data_RNO_20_9_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42114\,
            in1 => \N__34058\,
            in2 => \_gnd_net_\,
            in3 => \N__32210\,
            lcout => \sDAC_data_RNO_20Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_20_6_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_20Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52255\,
            ce => \N__36637\,
            sr => \N__51745\
        );

    \sDAC_data_RNO_21_3_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42112\,
            in1 => \N__36515\,
            in2 => \_gnd_net_\,
            in3 => \N__32408\,
            lcout => \sDAC_data_RNO_21Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_21_4_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42147\,
            in1 => \N__36503\,
            in2 => \_gnd_net_\,
            in3 => \N__32396\,
            lcout => \sDAC_data_RNO_21Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_21_5_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42113\,
            in1 => \N__36491\,
            in2 => \_gnd_net_\,
            in3 => \N__32378\,
            lcout => \sDAC_data_RNO_21Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_21_6_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42145\,
            in1 => \N__36776\,
            in2 => \_gnd_net_\,
            in3 => \N__32366\,
            lcout => \sDAC_data_RNO_21Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_4_3_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46779\,
            lcout => \sDAC_mem_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52245\,
            ce => \N__42640\,
            sr => \N__51730\
        );

    \sDAC_data_RNO_12_7_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42426\,
            in1 => \N__32342\,
            in2 => \N__42248\,
            in3 => \N__32318\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_7_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42211\,
            in1 => \N__41123\,
            in2 => \N__32330\,
            in3 => \N__44483\,
            lcout => \sDAC_data_RNO_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_4_4_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45509\,
            lcout => \sDAC_mem_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52245\,
            ce => \N__42640\,
            sr => \N__51730\
        );

    \sDAC_data_RNO_12_8_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__42432\,
            in1 => \N__32312\,
            in2 => \N__36479\,
            in3 => \N__42209\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_8_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42210\,
            in1 => \N__41111\,
            in2 => \N__32552\,
            in3 => \N__44471\,
            lcout => \sDAC_data_RNO_4Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_13_8_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42425\,
            in1 => \N__32537\,
            in2 => \N__42213\,
            in3 => \N__32486\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_8_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42149\,
            in1 => \N__32522\,
            in2 => \N__32513\,
            in3 => \N__32510\,
            lcout => \sDAC_data_RNO_5Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_6_5_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45067\,
            lcout => \sDAC_mem_6Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52234\,
            ce => \N__36553\,
            sr => \N__51718\
        );

    \sDAC_data_RNO_13_9_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42525\,
            in1 => \N__32480\,
            in2 => \N__42238\,
            in3 => \N__32444\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_9_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__44297\,
            in1 => \N__42153\,
            in2 => \N__32465\,
            in3 => \N__32462\,
            lcout => \sDAC_data_RNO_5Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_6_6_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50463\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_6Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52234\,
            ce => \N__36553\,
            sr => \N__51718\
        );

    \sDAC_data_RNO_16_10_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42424\,
            in1 => \N__32438\,
            in2 => \N__42212\,
            in3 => \N__32423\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_10_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42148\,
            in1 => \N__39830\,
            in2 => \N__32702\,
            in3 => \N__37028\,
            lcout => \sDAC_data_RNO_7Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_12_9_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__42576\,
            in1 => \N__32699\,
            in2 => \N__32672\,
            in3 => \N__42000\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_9_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__44459\,
            in1 => \N__41988\,
            in2 => \N__32687\,
            in3 => \N__41099\,
            lcout => \sDAC_data_RNO_4Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_4_6_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50516\,
            lcout => \sDAC_mem_4Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52224\,
            ce => \N__42636\,
            sr => \N__51707\
        );

    \sDAC_data_RNO_13_10_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42511\,
            in1 => \N__32663\,
            in2 => \N__42172\,
            in3 => \N__36569\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_10_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__41986\,
            in1 => \N__32648\,
            in2 => \N__32636\,
            in3 => \N__32633\,
            lcout => \sDAC_data_RNO_5Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_13_3_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42512\,
            in1 => \N__32621\,
            in2 => \N__42173\,
            in3 => \N__36611\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_3_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__41987\,
            in1 => \N__32606\,
            in2 => \N__32594\,
            in3 => \N__32591\,
            lcout => \sDAC_data_RNO_5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_13_4_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42510\,
            in1 => \N__32579\,
            in2 => \N__42171\,
            in3 => \N__36596\,
            lcout => \sDAC_data_2_13_bm_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_27_10_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42515\,
            in1 => \N__32873\,
            in2 => \N__42097\,
            in3 => \N__32861\,
            lcout => \sDAC_data_2_6_bm_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_2_7_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50009\,
            lcout => \sDAC_mem_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52218\,
            ce => \N__32855\,
            sr => \N__51699\
        );

    \sDAC_data_RNO_18_10_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41891\,
            in1 => \N__44597\,
            in2 => \_gnd_net_\,
            in3 => \N__32828\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_10_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__38166\,
            in1 => \N__38500\,
            in2 => \N__32813\,
            in3 => \N__32780\,
            lcout => \sDAC_data_2_24_ns_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_19_10_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41887\,
            in1 => \N__32810\,
            in2 => \_gnd_net_\,
            in3 => \N__32795\,
            lcout => \sDAC_data_RNO_19Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_10_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42521\,
            in1 => \N__32774\,
            in2 => \_gnd_net_\,
            in3 => \N__32759\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_10_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__41892\,
            in1 => \_gnd_net_\,
            in2 => \N__32741\,
            in3 => \N__32738\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_8Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_10_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011000110010"
        )
    port map (
            in0 => \N__38167\,
            in1 => \N__32720\,
            in2 => \N__32714\,
            in3 => \N__32711\,
            lcout => \sDAC_data_RNO_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \button_debounce_counter_esr_RNO_0_23_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__45722\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49427\,
            lcout => \LED3_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNITC6L_19_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33374\,
            in1 => \N__33257\,
            in2 => \N__33168\,
            in3 => \N__33047\,
            lcout => g0_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.spi_cs_i_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__47903\,
            in1 => \N__48041\,
            in2 => \_gnd_net_\,
            in3 => \N__47947\,
            lcout => \spi_slave_inst.spi_cs_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_10_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110110101"
        )
    port map (
            in0 => \N__37343\,
            in1 => \N__32879\,
            in2 => \N__37481\,
            in3 => \N__33404\,
            lcout => OPEN,
            ltout => \sDAC_data_2_41_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_10_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111000001110"
        )
    port map (
            in0 => \N__32936\,
            in1 => \N__37471\,
            in2 => \N__32930\,
            in3 => \N__34943\,
            lcout => \sDAC_data_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_0_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35072\,
            in1 => \N__35039\,
            in2 => \N__35057\,
            in3 => \N__35087\,
            lcout => \sbuttonModeStatus_0_sqmuxa_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_21_10_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41804\,
            in1 => \N__36716\,
            in2 => \_gnd_net_\,
            in3 => \N__32909\,
            lcout => \sDAC_data_RNO_21Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_28_10_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41807\,
            in1 => \N__38963\,
            in2 => \_gnd_net_\,
            in3 => \N__33518\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_28Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_10_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__38452\,
            in1 => \N__38115\,
            in2 => \N__32891\,
            in3 => \N__33524\,
            lcout => OPEN,
            ltout => \sDAC_data_2_32_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_10_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__38116\,
            in1 => \N__32888\,
            in2 => \N__32882\,
            in3 => \N__33548\,
            lcout => \sDAC_data_RNO_10Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_20_10_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41805\,
            in1 => \N__34046\,
            in2 => \_gnd_net_\,
            in3 => \N__36653\,
            lcout => \sDAC_data_RNO_20Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_29_10_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34079\,
            in2 => \N__33542\,
            in3 => \N__41806\,
            lcout => \sDAC_data_RNO_29Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_16_7_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50056\,
            lcout => \sDAC_mem_16Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52235\,
            ce => \N__33512\,
            sr => \N__51684\
        );

    \sDAC_data_RNO_25_10_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38448\,
            in1 => \N__33470\,
            in2 => \N__38203\,
            in3 => \N__33464\,
            lcout => \sDAC_data_2_39_ns_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_10_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41606\,
            in1 => \N__33458\,
            in2 => \_gnd_net_\,
            in3 => \N__33449\,
            lcout => \sDAC_data_RNO_24Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_10_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41609\,
            in1 => \N__33434\,
            in2 => \_gnd_net_\,
            in3 => \N__33395\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_23Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_10_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__38117\,
            in1 => \N__33419\,
            in2 => \N__33413\,
            in3 => \N__33410\,
            lcout => \sDAC_data_RNO_11Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_28_7_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50057\,
            lcout => \sDAC_mem_28Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52246\,
            ce => \N__37808\,
            sr => \N__51679\
        );

    \sDAC_data_RNO_31_3_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41605\,
            in1 => \N__33650\,
            in2 => \_gnd_net_\,
            in3 => \N__33644\,
            lcout => \sDAC_data_RNO_31Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_30_3_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41608\,
            in1 => \N__41324\,
            in2 => \_gnd_net_\,
            in3 => \N__33635\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_30Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_25_3_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__38402\,
            in1 => \N__38121\,
            in2 => \N__33620\,
            in3 => \N__33617\,
            lcout => OPEN,
            ltout => \sDAC_data_2_39_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_3_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__38122\,
            in1 => \N__33611\,
            in2 => \N__33605\,
            in3 => \N__33845\,
            lcout => \sDAC_data_RNO_11Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_21_7_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41866\,
            in1 => \N__36764\,
            in2 => \_gnd_net_\,
            in3 => \N__33587\,
            lcout => \sDAC_data_RNO_21Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_22_4_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45603\,
            lcout => \sDAC_mem_22Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52256\,
            ce => \N__33893\,
            sr => \N__51671\
        );

    \sDAC_data_RNO_21_8_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41868\,
            in1 => \N__36746\,
            in2 => \_gnd_net_\,
            in3 => \N__33566\,
            lcout => \sDAC_data_RNO_21Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_22_5_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45118\,
            lcout => \sDAC_mem_22Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52256\,
            ce => \N__33893\,
            sr => \N__51671\
        );

    \sDAC_data_RNO_21_9_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41867\,
            in1 => \N__36728\,
            in2 => \_gnd_net_\,
            in3 => \N__33899\,
            lcout => \sDAC_data_RNO_21Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_22_6_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50542\,
            lcout => \sDAC_mem_22Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52256\,
            ce => \N__33893\,
            sr => \N__51671\
        );

    \sDAC_data_RNO_23_3_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41865\,
            in1 => \N__33869\,
            in2 => \_gnd_net_\,
            in3 => \N__33860\,
            lcout => \sDAC_data_RNO_23Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_6_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41985\,
            in1 => \N__33839\,
            in2 => \_gnd_net_\,
            in3 => \N__33827\,
            lcout => \sDAC_data_RNO_23Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_4_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35344\,
            in1 => \N__35122\,
            in2 => \N__35330\,
            in3 => \N__35359\,
            lcout => \sbuttonModeStatus_0_sqmuxa_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_5_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35180\,
            in1 => \N__35141\,
            in2 => \N__35285\,
            in3 => \N__35162\,
            lcout => OPEN,
            ltout => \sbuttonModeStatus_0_sqmuxa_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_2_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38843\,
            in1 => \N__38765\,
            in2 => \N__33812\,
            in3 => \N__33809\,
            lcout => \sbuttonModeStatus_0_sqmuxa_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_6_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__33791\,
            in1 => \N__40072\,
            in2 => \_gnd_net_\,
            in3 => \N__33773\,
            lcout => \sEEPonPoff_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_nWE_obuf_RNO_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__48961\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34015\,
            lcout => \RAM_nWE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sRead_data_RNO_0_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39163\,
            in2 => \_gnd_net_\,
            in3 => \N__39139\,
            lcout => OPEN,
            ltout => \sRead_data_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sRead_data_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001100"
        )
    port map (
            in0 => \N__33983\,
            in1 => \N__43735\,
            in2 => \N__34031\,
            in3 => \N__48952\,
            lcout => \sRead_dataZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52277\,
            ce => 'H',
            sr => \N__51658\
        );

    \sCounterRAM_RNIS8L63_1_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39029\,
            in1 => \N__33965\,
            in2 => \N__39608\,
            in3 => \N__33971\,
            lcout => \N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sSPI_MSB0LSB1_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001001111001100"
        )
    port map (
            in0 => \N__43336\,
            in1 => \N__39164\,
            in2 => \N__43487\,
            in3 => \N__39140\,
            lcout => \sSPI_MSB0LSBZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52277\,
            ce => 'H',
            sr => \N__51658\
        );

    \sADC_clk_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__34006\,
            in1 => \N__43335\,
            in2 => \N__46970\,
            in3 => \N__43446\,
            lcout => \ADC_clk_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52277\,
            ce => 'H',
            sr => \N__51658\
        );

    \sRead_data_RNI74VQ_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__33982\,
            in1 => \N__39548\,
            in2 => \_gnd_net_\,
            in3 => \N__39566\,
            lcout => spi_data_miso_0_sqmuxa_2_i_o2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterRAM_RNISREI1_7_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__39530\,
            in1 => \N__39047\,
            in2 => \N__39479\,
            in3 => \N__39584\,
            lcout => spi_data_miso_0_sqmuxa_2_i_o2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_1_3_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33959\,
            lcout => \RAM_DATA_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52311\,
            ce => \N__51890\,
            sr => \N__51647\
        );

    \sDAC_mem_19_4_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45508\,
            lcout => \sDAC_mem_19Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52290\,
            ce => \N__34997\,
            sr => \N__51806\
        );

    \sDAC_mem_19_5_LC_16_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44982\,
            lcout => \sDAC_mem_19Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52290\,
            ce => \N__34997\,
            sr => \N__51806\
        );

    \sDAC_mem_19_6_LC_16_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50484\,
            lcout => \sDAC_mem_19Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52290\,
            ce => \N__34997\,
            sr => \N__51806\
        );

    \sDAC_mem_19_7_LC_16_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50054\,
            lcout => \sDAC_mem_19Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52290\,
            ce => \N__34997\,
            sr => \N__51806\
        );

    \sDAC_mem_21_0_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46385\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_21Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52278\,
            ce => \N__34247\,
            sr => \N__51797\
        );

    \sDAC_mem_21_1_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51053\,
            lcout => \sDAC_mem_21Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52278\,
            ce => \N__34247\,
            sr => \N__51797\
        );

    \sDAC_mem_21_2_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47348\,
            lcout => \sDAC_mem_21Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52278\,
            ce => \N__34247\,
            sr => \N__51797\
        );

    \sDAC_mem_21_3_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46751\,
            lcout => \sDAC_mem_21Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52278\,
            ce => \N__34247\,
            sr => \N__51797\
        );

    \sDAC_mem_21_4_LC_16_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45507\,
            lcout => \sDAC_mem_21Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52278\,
            ce => \N__34247\,
            sr => \N__51797\
        );

    \sDAC_mem_21_5_LC_16_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__44981\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_21Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52278\,
            ce => \N__34247\,
            sr => \N__51797\
        );

    \sDAC_mem_21_6_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50483\,
            lcout => \sDAC_mem_21Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52278\,
            ce => \N__34247\,
            sr => \N__51797\
        );

    \sDAC_mem_21_7_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50053\,
            lcout => \sDAC_mem_21Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52278\,
            ce => \N__34247\,
            sr => \N__51797\
        );

    \sDAC_mem_3_4_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45349\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52268\,
            ce => \N__44237\,
            sr => \N__51783\
        );

    \sDAC_data_RNO_27_7_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42557\,
            in1 => \N__34235\,
            in2 => \N__42264\,
            in3 => \N__34223\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_7_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42095\,
            in1 => \N__34211\,
            in2 => \N__34196\,
            in3 => \N__34193\,
            lcout => \sDAC_data_RNO_15Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_7_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42558\,
            in1 => \N__34181\,
            in2 => \N__42265\,
            in3 => \N__34169\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_7_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__36800\,
            in1 => \N__42259\,
            in2 => \N__34157\,
            in3 => \N__39680\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_7Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_7_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010101100100"
        )
    port map (
            in0 => \N__34154\,
            in1 => \N__38131\,
            in2 => \N__34145\,
            in3 => \N__34121\,
            lcout => \sDAC_data_RNO_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_7_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42096\,
            in1 => \N__34136\,
            in2 => \_gnd_net_\,
            in3 => \N__34097\,
            lcout => \sDAC_data_RNO_8Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_7_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42556\,
            in1 => \N__34115\,
            in2 => \_gnd_net_\,
            in3 => \N__34106\,
            lcout => \sDAC_data_RNO_17Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_3_6_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52257\,
            ce => \N__44244\,
            sr => \N__51771\
        );

    \sDAC_data_RNO_27_9_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42551\,
            in1 => \N__34376\,
            in2 => \N__42239\,
            in3 => \N__34364\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_9_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42165\,
            in1 => \N__34355\,
            in2 => \N__34346\,
            in3 => \N__34343\,
            lcout => \sDAC_data_RNO_15Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_9_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42552\,
            in1 => \N__34331\,
            in2 => \_gnd_net_\,
            in3 => \N__34316\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_9_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42157\,
            in2 => \N__34301\,
            in3 => \N__34298\,
            lcout => \sDAC_data_RNO_8Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_9_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__34289\,
            in1 => \N__42166\,
            in2 => \N__42575\,
            in3 => \N__34277\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_9_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42167\,
            in1 => \N__39842\,
            in2 => \N__34265\,
            in3 => \N__37040\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_7Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_9_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101100010"
        )
    port map (
            in0 => \N__38031\,
            in1 => \N__36983\,
            in2 => \N__34262\,
            in3 => \N__34259\,
            lcout => \sDAC_data_RNO_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_32_6_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50486\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_32Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52247\,
            ce => \N__41265\,
            sr => \N__51758\
        );

    \sDAC_data_RNO_26_9_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42430\,
            in1 => \N__44324\,
            in2 => \_gnd_net_\,
            in3 => \N__44423\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_9_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__42111\,
            in1 => \_gnd_net_\,
            in2 => \N__34469\,
            in3 => \N__34466\,
            lcout => \sDAC_data_RNO_14Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_20_3_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34454\,
            in1 => \N__42105\,
            in2 => \_gnd_net_\,
            in3 => \N__36449\,
            lcout => \sDAC_data_RNO_20Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_20_4_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42104\,
            in1 => \N__34445\,
            in2 => \_gnd_net_\,
            in3 => \N__36437\,
            lcout => \sDAC_data_RNO_20Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_20_5_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34424\,
            in1 => \N__42109\,
            in2 => \_gnd_net_\,
            in3 => \N__36425\,
            lcout => \sDAC_data_RNO_20Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_20_6_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__36413\,
            in1 => \_gnd_net_\,
            in2 => \N__42214\,
            in3 => \N__34415\,
            lcout => \sDAC_data_RNO_20Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_20_7_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34394\,
            in1 => \N__42110\,
            in2 => \_gnd_net_\,
            in3 => \N__36662\,
            lcout => \sDAC_data_RNO_20Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_pointer_RNI3NFH_1_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42168\,
            in2 => \N__38552\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \sDAC_mem_pointer_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_pointer_2_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__37632\,
            in1 => \N__38001\,
            in2 => \_gnd_net_\,
            in3 => \N__34577\,
            lcout => \sDAC_mem_pointerZ0Z_2\,
            ltout => OPEN,
            carryin => \sDAC_mem_pointer_0_cry_1\,
            carryout => \sDAC_mem_pointer_0_cry_2\,
            clk => \N__48462\,
            ce => \N__43949\,
            sr => \N__51746\
        );

    \sDAC_mem_pointer_3_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__37635\,
            in1 => \N__37327\,
            in2 => \_gnd_net_\,
            in3 => \N__34574\,
            lcout => \sDAC_mem_pointerZ0Z_3\,
            ltout => OPEN,
            carryin => \sDAC_mem_pointer_0_cry_2\,
            carryout => \sDAC_mem_pointer_0_cry_3\,
            clk => \N__48462\,
            ce => \N__43949\,
            sr => \N__51746\
        );

    \sDAC_mem_pointer_4_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__37633\,
            in1 => \N__37419\,
            in2 => \_gnd_net_\,
            in3 => \N__34571\,
            lcout => \sDAC_mem_pointerZ0Z_4\,
            ltout => OPEN,
            carryin => \sDAC_mem_pointer_0_cry_3\,
            carryout => \sDAC_mem_pointer_0_cry_4\,
            clk => \N__48462\,
            ce => \N__43949\,
            sr => \N__51746\
        );

    \sDAC_mem_pointer_5_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__42433\,
            in1 => \N__37634\,
            in2 => \_gnd_net_\,
            in3 => \N__34568\,
            lcout => \sDAC_mem_pointerZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48462\,
            ce => \N__43949\,
            sr => \N__51746\
        );

    \sDAC_mem_3_2_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47447\,
            lcout => \sDAC_mem_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52225\,
            ce => \N__44246\,
            sr => \N__51731\
        );

    \sDAC_data_RNO_27_5_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42427\,
            in1 => \N__34565\,
            in2 => \N__42240\,
            in3 => \N__34553\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_5_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42143\,
            in1 => \N__34541\,
            in2 => \N__34523\,
            in3 => \N__34520\,
            lcout => \sDAC_data_RNO_15Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_5_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42428\,
            in1 => \N__34514\,
            in2 => \_gnd_net_\,
            in3 => \N__34502\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_5_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42161\,
            in2 => \N__34487\,
            in3 => \N__34484\,
            lcout => \sDAC_data_RNO_8Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_5_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42429\,
            in1 => \N__34757\,
            in2 => \N__42241\,
            in3 => \N__34742\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_5_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42144\,
            in1 => \N__39884\,
            in2 => \N__34727\,
            in3 => \N__36821\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_7Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_5_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101100010"
        )
    port map (
            in0 => \N__37997\,
            in1 => \N__34724\,
            in2 => \N__34715\,
            in3 => \N__34712\,
            lcout => \sDAC_data_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_3_0_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46314\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52219\,
            ce => \N__44245\,
            sr => \N__51719\
        );

    \sDAC_data_RNO_27_3_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42522\,
            in1 => \N__34706\,
            in2 => \N__42174\,
            in3 => \N__34694\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_3_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__41983\,
            in1 => \N__34682\,
            in2 => \N__34664\,
            in3 => \N__34661\,
            lcout => \sDAC_data_RNO_15Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_3_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42523\,
            in1 => \N__34655\,
            in2 => \_gnd_net_\,
            in3 => \N__34637\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_3_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42006\,
            in2 => \N__34622\,
            in3 => \N__34619\,
            lcout => \sDAC_data_RNO_8Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_3_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42524\,
            in1 => \N__34607\,
            in2 => \N__42175\,
            in3 => \N__34592\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_3_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__41984\,
            in1 => \N__39908\,
            in2 => \N__34898\,
            in3 => \N__36845\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_7Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_3_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101100010"
        )
    port map (
            in0 => \N__38097\,
            in1 => \N__34895\,
            in2 => \N__34883\,
            in3 => \N__34880\,
            lcout => \sDAC_data_RNO_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_8_3_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__40428\,
            in1 => \N__34874\,
            in2 => \_gnd_net_\,
            in3 => \N__40028\,
            lcout => \sDAC_mem_19_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_19_0_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46315\,
            lcout => \sDAC_mem_19Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52212\,
            ce => \N__34990\,
            sr => \N__51708\
        );

    \sDAC_data_RNO_29_3_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41885\,
            in1 => \N__34829\,
            in2 => \_gnd_net_\,
            in3 => \N__34823\,
            lcout => \sDAC_data_RNO_29Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_19_1_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50985\,
            lcout => \sDAC_mem_19Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52212\,
            ce => \N__34990\,
            sr => \N__51708\
        );

    \sDAC_data_RNO_29_4_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41884\,
            in1 => \N__34808\,
            in2 => \_gnd_net_\,
            in3 => \N__34802\,
            lcout => \sDAC_data_RNO_29Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_19_2_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47496\,
            lcout => \sDAC_mem_19Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52212\,
            ce => \N__34990\,
            sr => \N__51708\
        );

    \sDAC_data_RNO_29_5_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41886\,
            in1 => \N__34775\,
            in2 => \_gnd_net_\,
            in3 => \N__34769\,
            lcout => \sDAC_data_RNO_29Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_19_3_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46854\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_19Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52212\,
            ce => \N__34990\,
            sr => \N__51708\
        );

    \sDAC_data_RNO_15_10_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__34976\,
            in1 => \N__44261\,
            in2 => \N__42170\,
            in3 => \N__34964\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_15Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_10_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__38231\,
            in1 => \N__38526\,
            in2 => \N__34958\,
            in3 => \N__34904\,
            lcout => OPEN,
            ltout => \sDAC_data_2_14_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_10_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__38030\,
            in1 => \N__34955\,
            in2 => \N__34946\,
            in3 => \N__34916\,
            lcout => \sDAC_data_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_26_10_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44414\,
            in1 => \N__42513\,
            in2 => \_gnd_net_\,
            in3 => \N__44543\,
            lcout => \sDAC_data_RNO_26Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_12_10_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42514\,
            in1 => \N__34937\,
            in2 => \N__42169\,
            in3 => \N__36461\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_10_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__41982\,
            in1 => \N__41087\,
            in2 => \N__34919\,
            in3 => \N__44447\,
            lcout => \sDAC_data_RNO_4Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_10_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41975\,
            in1 => \N__39623\,
            in2 => \_gnd_net_\,
            in3 => \N__34910\,
            lcout => \sDAC_data_RNO_14Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_button_debounce_counter_cry_1_c_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45772\,
            in2 => \N__45751\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_13_0_\,
            carryout => un1_button_debounce_counter_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \button_debounce_counter_2_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49428\,
            in1 => \N__35101\,
            in2 => \_gnd_net_\,
            in3 => \N__35090\,
            lcout => \button_debounce_counterZ0Z_2\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_1,
            carryout => un1_button_debounce_counter_cry_2,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__45714\
        );

    \button_debounce_counter_3_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49191\,
            in1 => \N__35086\,
            in2 => \_gnd_net_\,
            in3 => \N__35075\,
            lcout => \button_debounce_counterZ0Z_3\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_2,
            carryout => un1_button_debounce_counter_cry_3,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__45714\
        );

    \button_debounce_counter_4_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49429\,
            in1 => \N__35071\,
            in2 => \_gnd_net_\,
            in3 => \N__35060\,
            lcout => \button_debounce_counterZ0Z_4\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_3,
            carryout => un1_button_debounce_counter_cry_4,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__45714\
        );

    \button_debounce_counter_5_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49192\,
            in1 => \N__35053\,
            in2 => \_gnd_net_\,
            in3 => \N__35042\,
            lcout => \button_debounce_counterZ0Z_5\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_4,
            carryout => un1_button_debounce_counter_cry_5,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__45714\
        );

    \button_debounce_counter_6_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49430\,
            in1 => \N__35035\,
            in2 => \_gnd_net_\,
            in3 => \N__35024\,
            lcout => \button_debounce_counterZ0Z_6\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_5,
            carryout => un1_button_debounce_counter_cry_6,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__45714\
        );

    \button_debounce_counter_7_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49193\,
            in1 => \N__38815\,
            in2 => \_gnd_net_\,
            in3 => \N__35021\,
            lcout => \button_debounce_counterZ0Z_7\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_6,
            carryout => un1_button_debounce_counter_cry_7,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__45714\
        );

    \button_debounce_counter_8_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49431\,
            in1 => \N__38779\,
            in2 => \_gnd_net_\,
            in3 => \N__35018\,
            lcout => \button_debounce_counterZ0Z_8\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_7,
            carryout => un1_button_debounce_counter_cry_8,
            clk => \N__48476\,
            ce => 'H',
            sr => \N__45714\
        );

    \button_debounce_counter_9_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49295\,
            in1 => \N__38830\,
            in2 => \_gnd_net_\,
            in3 => \N__35015\,
            lcout => \button_debounce_counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_16_14_0_\,
            carryout => un1_button_debounce_counter_cry_9,
            clk => \N__48480\,
            ce => 'H',
            sr => \N__45715\
        );

    \button_debounce_counter_10_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49288\,
            in1 => \N__38794\,
            in2 => \_gnd_net_\,
            in3 => \N__35195\,
            lcout => \button_debounce_counterZ0Z_10\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_9,
            carryout => un1_button_debounce_counter_cry_10,
            clk => \N__48480\,
            ce => 'H',
            sr => \N__45715\
        );

    \button_debounce_counter_11_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49292\,
            in1 => \N__38857\,
            in2 => \_gnd_net_\,
            in3 => \N__35192\,
            lcout => \button_debounce_counterZ0Z_11\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_10,
            carryout => un1_button_debounce_counter_cry_11,
            clk => \N__48480\,
            ce => 'H',
            sr => \N__45715\
        );

    \button_debounce_counter_12_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49289\,
            in1 => \N__38890\,
            in2 => \_gnd_net_\,
            in3 => \N__35189\,
            lcout => \button_debounce_counterZ0Z_12\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_11,
            carryout => un1_button_debounce_counter_cry_12,
            clk => \N__48480\,
            ce => 'H',
            sr => \N__45715\
        );

    \button_debounce_counter_13_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49293\,
            in1 => \N__38905\,
            in2 => \_gnd_net_\,
            in3 => \N__35186\,
            lcout => \button_debounce_counterZ0Z_13\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_12,
            carryout => un1_button_debounce_counter_cry_13,
            clk => \N__48480\,
            ce => 'H',
            sr => \N__45715\
        );

    \button_debounce_counter_14_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49290\,
            in1 => \N__38872\,
            in2 => \_gnd_net_\,
            in3 => \N__35183\,
            lcout => \button_debounce_counterZ0Z_14\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_13,
            carryout => un1_button_debounce_counter_cry_14,
            clk => \N__48480\,
            ce => 'H',
            sr => \N__45715\
        );

    \button_debounce_counter_15_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49294\,
            in1 => \N__35179\,
            in2 => \_gnd_net_\,
            in3 => \N__35165\,
            lcout => \button_debounce_counterZ0Z_15\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_14,
            carryout => un1_button_debounce_counter_cry_15,
            clk => \N__48480\,
            ce => 'H',
            sr => \N__45715\
        );

    \button_debounce_counter_16_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49291\,
            in1 => \N__35158\,
            in2 => \_gnd_net_\,
            in3 => \N__35144\,
            lcout => \button_debounce_counterZ0Z_16\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_15,
            carryout => un1_button_debounce_counter_cry_16,
            clk => \N__48480\,
            ce => 'H',
            sr => \N__45715\
        );

    \button_debounce_counter_17_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49302\,
            in1 => \N__35140\,
            in2 => \_gnd_net_\,
            in3 => \N__35126\,
            lcout => \button_debounce_counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => un1_button_debounce_counter_cry_17,
            clk => \N__48483\,
            ce => 'H',
            sr => \N__45716\
        );

    \button_debounce_counter_18_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49305\,
            in1 => \N__35123\,
            in2 => \_gnd_net_\,
            in3 => \N__35111\,
            lcout => \button_debounce_counterZ0Z_18\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_17,
            carryout => un1_button_debounce_counter_cry_18,
            clk => \N__48483\,
            ce => 'H',
            sr => \N__45716\
        );

    \button_debounce_counter_19_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49303\,
            in1 => \N__35360\,
            in2 => \_gnd_net_\,
            in3 => \N__35348\,
            lcout => \button_debounce_counterZ0Z_19\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_18,
            carryout => un1_button_debounce_counter_cry_19,
            clk => \N__48483\,
            ce => 'H',
            sr => \N__45716\
        );

    \button_debounce_counter_20_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49306\,
            in1 => \N__35345\,
            in2 => \_gnd_net_\,
            in3 => \N__35333\,
            lcout => \button_debounce_counterZ0Z_20\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_19,
            carryout => un1_button_debounce_counter_cry_20,
            clk => \N__48483\,
            ce => 'H',
            sr => \N__45716\
        );

    \button_debounce_counter_21_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49304\,
            in1 => \N__35329\,
            in2 => \_gnd_net_\,
            in3 => \N__35315\,
            lcout => \button_debounce_counterZ0Z_21\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_20,
            carryout => un1_button_debounce_counter_cry_21,
            clk => \N__48483\,
            ce => 'H',
            sr => \N__45716\
        );

    \button_debounce_counter_22_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__49307\,
            in1 => \N__35305\,
            in2 => \_gnd_net_\,
            in3 => \N__35291\,
            lcout => \button_debounce_counterZ0Z_22\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_21,
            carryout => un1_button_debounce_counter_cry_22,
            clk => \N__48483\,
            ce => 'H',
            sr => \N__45716\
        );

    \un1_button_debounce_counter_cry_22_c_THRU_CRY_0_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52510\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_22,
            carryout => \un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_button_debounce_counter_cry_22_c_THRU_CRY_1_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__52586\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO\,
            carryout => \un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \button_debounce_counter_esr_23_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35284\,
            in2 => \_gnd_net_\,
            in3 => \N__35288\,
            lcout => \button_debounce_counterZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48486\,
            ce => \N__35270\,
            sr => \N__45717\
        );

    \sRAM_ADD_5_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__43344\,
            in1 => \N__35255\,
            in2 => \N__43491\,
            in3 => \N__35237\,
            lcout => \RAM_ADD_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52269\,
            ce => \N__43218\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_0_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__35909\,
            in1 => \N__43450\,
            in2 => \N__35891\,
            in3 => \N__43337\,
            lcout => \RAM_ADD_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52269\,
            ce => \N__43218\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_10_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__43338\,
            in1 => \N__35846\,
            in2 => \N__43488\,
            in3 => \N__35828\,
            lcout => \RAM_ADD_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52269\,
            ce => \N__43218\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_11_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__35774\,
            in1 => \N__43454\,
            in2 => \N__35756\,
            in3 => \N__43339\,
            lcout => \RAM_ADD_c_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52269\,
            ce => \N__43218\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_12_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__43340\,
            in1 => \N__35705\,
            in2 => \N__43489\,
            in3 => \N__35678\,
            lcout => \RAM_ADD_c_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52269\,
            ce => \N__43218\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_13_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__35639\,
            in1 => \N__43458\,
            in2 => \N__35621\,
            in3 => \N__43341\,
            lcout => \RAM_ADD_c_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52269\,
            ce => \N__43218\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_14_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__43342\,
            in1 => \N__35576\,
            in2 => \N__43490\,
            in3 => \N__35549\,
            lcout => \RAM_ADD_c_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52269\,
            ce => \N__43218\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_15_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__35504\,
            in1 => \N__43462\,
            in2 => \N__35486\,
            in3 => \N__43343\,
            lcout => \RAM_ADD_c_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52269\,
            ce => \N__43218\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_16_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__35432\,
            in1 => \N__43492\,
            in2 => \N__35414\,
            in3 => \N__43348\,
            lcout => \RAM_ADD_c_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52279\,
            ce => \N__43226\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_17_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__43349\,
            in1 => \N__36404\,
            in2 => \N__36377\,
            in3 => \N__43496\,
            lcout => \RAM_ADD_c_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52279\,
            ce => \N__43226\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_18_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__36338\,
            in1 => \N__43493\,
            in2 => \N__36311\,
            in3 => \N__43350\,
            lcout => \RAM_ADD_c_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52279\,
            ce => \N__43226\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_9_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__43355\,
            in1 => \N__36266\,
            in2 => \N__36239\,
            in3 => \N__43499\,
            lcout => \RAM_ADD_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52279\,
            ce => \N__43226\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_7_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__36197\,
            in1 => \N__43495\,
            in2 => \N__36170\,
            in3 => \N__43354\,
            lcout => \RAM_ADD_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52279\,
            ce => \N__43226\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_2_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__43352\,
            in1 => \N__36134\,
            in2 => \N__36119\,
            in3 => \N__43497\,
            lcout => \RAM_ADD_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52279\,
            ce => \N__43226\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_1_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__36074\,
            in1 => \N__43494\,
            in2 => \N__36047\,
            in3 => \N__43351\,
            lcout => \RAM_ADD_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52279\,
            ce => \N__43226\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_6_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__43353\,
            in1 => \N__36017\,
            in2 => \N__35990\,
            in3 => \N__43498\,
            lcout => \RAM_ADD_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52279\,
            ce => \N__43226\,
            sr => \_gnd_net_\
        );

    \RAM_DATA_1_4_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35951\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RAM_DATA_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52301\,
            ce => \N__51895\,
            sr => \N__51650\
        );

    \sDAC_mem_pointer_6_LC_17_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_mem_pointerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48447\,
            ce => \N__43957\,
            sr => \N__51823\
        );

    \sDAC_mem_pointer_7_LC_17_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_mem_pointerZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48447\,
            ce => \N__43957\,
            sr => \N__51823\
        );

    \sDAC_mem_4_2_LC_17_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47438\,
            lcout => \sDAC_mem_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52281\,
            ce => \N__42626\,
            sr => \N__51813\
        );

    \sDAC_mem_4_5_LC_17_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45104\,
            lcout => \sDAC_mem_4Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52281\,
            ce => \N__42626\,
            sr => \N__51813\
        );

    \sDAC_mem_4_7_LC_17_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50055\,
            lcout => \sDAC_mem_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52281\,
            ce => \N__42626\,
            sr => \N__51813\
        );

    \sDAC_mem_20_0_LC_17_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46386\,
            lcout => \sDAC_mem_20Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52270\,
            ce => \N__36638\,
            sr => \N__51807\
        );

    \sDAC_mem_20_1_LC_17_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51054\,
            lcout => \sDAC_mem_20Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52270\,
            ce => \N__36638\,
            sr => \N__51807\
        );

    \sDAC_mem_20_2_LC_17_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47437\,
            lcout => \sDAC_mem_20Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52270\,
            ce => \N__36638\,
            sr => \N__51807\
        );

    \sDAC_mem_20_3_LC_17_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46752\,
            lcout => \sDAC_mem_20Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52270\,
            ce => \N__36638\,
            sr => \N__51807\
        );

    \sDAC_mem_20_4_LC_17_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45558\,
            lcout => \sDAC_mem_20Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52270\,
            ce => \N__36638\,
            sr => \N__51807\
        );

    \sDAC_mem_20_7_LC_17_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49865\,
            lcout => \sDAC_mem_20Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52270\,
            ce => \N__36638\,
            sr => \N__51807\
        );

    \sDAC_mem_6_0_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46388\,
            lcout => \sDAC_mem_6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52258\,
            ce => \N__36554\,
            sr => \N__51798\
        );

    \sDAC_mem_6_1_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51052\,
            lcout => \sDAC_mem_6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52258\,
            ce => \N__36554\,
            sr => \N__51798\
        );

    \sDAC_mem_6_4_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45350\,
            lcout => \sDAC_mem_6Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52258\,
            ce => \N__36554\,
            sr => \N__51798\
        );

    \sDAC_mem_6_7_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49847\,
            lcout => \sDAC_mem_6Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52258\,
            ce => \N__36554\,
            sr => \N__51798\
        );

    \sDAC_mem_23_0_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46387\,
            lcout => \sDAC_mem_23Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52248\,
            ce => \N__36701\,
            sr => \N__51784\
        );

    \sDAC_mem_23_1_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51055\,
            lcout => \sDAC_mem_23Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52248\,
            ce => \N__36701\,
            sr => \N__51784\
        );

    \sDAC_mem_23_2_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47446\,
            lcout => \sDAC_mem_23Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52248\,
            ce => \N__36701\,
            sr => \N__51784\
        );

    \sDAC_mem_23_3_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46858\,
            lcout => \sDAC_mem_23Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52248\,
            ce => \N__36701\,
            sr => \N__51784\
        );

    \sDAC_mem_23_4_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45559\,
            lcout => \sDAC_mem_23Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52248\,
            ce => \N__36701\,
            sr => \N__51784\
        );

    \sDAC_mem_23_5_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45100\,
            lcout => \sDAC_mem_23Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52248\,
            ce => \N__36701\,
            sr => \N__51784\
        );

    \sDAC_mem_23_6_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50485\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_23Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52248\,
            ce => \N__36701\,
            sr => \N__51784\
        );

    \sDAC_mem_23_7_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49866\,
            lcout => \sDAC_mem_23Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52248\,
            ce => \N__36701\,
            sr => \N__51784\
        );

    \sDAC_mem_32_3_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46920\,
            lcout => \sDAC_mem_32Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52236\,
            ce => \N__41258\,
            sr => \N__51772\
        );

    \sDAC_data_RNO_26_6_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42422\,
            in1 => \N__44360\,
            in2 => \_gnd_net_\,
            in3 => \N__44102\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_6_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42189\,
            in2 => \N__36683\,
            in3 => \N__36680\,
            lcout => \sDAC_data_RNO_14Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_26_7_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__42423\,
            in1 => \N__44093\,
            in2 => \_gnd_net_\,
            in3 => \N__44348\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_7_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42190\,
            in2 => \N__36884\,
            in3 => \N__36869\,
            lcout => \sDAC_data_RNO_14Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_32_4_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45592\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_32Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52236\,
            ce => \N__41258\,
            sr => \N__51772\
        );

    \sDAC_data_RNO_26_8_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42431\,
            in1 => \N__44336\,
            in2 => \_gnd_net_\,
            in3 => \N__44084\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_8_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__42191\,
            in1 => \_gnd_net_\,
            in2 => \N__36863\,
            in3 => \N__39632\,
            lcout => \sDAC_data_RNO_14Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_9_0_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46352\,
            lcout => \sDAC_mem_9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52226\,
            ce => \N__39818\,
            sr => \N__51759\
        );

    \sDAC_mem_9_1_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51070\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52226\,
            ce => \N__39818\,
            sr => \N__51759\
        );

    \sDAC_mem_9_2_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47439\,
            lcout => \sDAC_mem_9Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52226\,
            ce => \N__39818\,
            sr => \N__51759\
        );

    \sDAC_mem_9_3_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46859\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_9Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52226\,
            ce => \N__39818\,
            sr => \N__51759\
        );

    \sDAC_mem_9_4_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45560\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_9Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52226\,
            ce => \N__39818\,
            sr => \N__51759\
        );

    \sDAC_mem_9_5_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45103\,
            lcout => \sDAC_mem_9Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52226\,
            ce => \N__39818\,
            sr => \N__51759\
        );

    \sDAC_mem_9_6_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50487\,
            lcout => \sDAC_mem_9Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52226\,
            ce => \N__39818\,
            sr => \N__51759\
        );

    \sDAC_mem_9_7_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49867\,
            lcout => \sDAC_mem_9Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52226\,
            ce => \N__39818\,
            sr => \N__51759\
        );

    \sDAC_data_RNO_19_9_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41841\,
            in1 => \N__37016\,
            in2 => \_gnd_net_\,
            in3 => \N__37007\,
            lcout => \sDAC_data_RNO_19Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_9_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42142\,
            in1 => \N__44609\,
            in2 => \_gnd_net_\,
            in3 => \N__36971\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_9_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__38096\,
            in1 => \N__38460\,
            in2 => \N__36992\,
            in3 => \N__36989\,
            lcout => \sDAC_data_2_24_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_12_6_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50488\,
            lcout => \sDAC_mem_12Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52220\,
            ce => \N__36964\,
            sr => \N__51747\
        );

    \sDAC_mem_pointer_RNIAIV21_3_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__38095\,
            in1 => \N__38459\,
            in2 => \N__42074\,
            in3 => \N__37305\,
            lcout => OPEN,
            ltout => \op_le_op_le_un15_sdacdynlt4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_pointer_RNI4LV52_4_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__37390\,
            in1 => \N__42411\,
            in2 => \N__36902\,
            in3 => \N__37172\,
            lcout => un17_sdacdyn_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_pointer_RNIF3GH_6_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37196\,
            in2 => \_gnd_net_\,
            in3 => \N__37181\,
            lcout => un17_sdacdyn_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_26_3_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42421\,
            in1 => \N__44390\,
            in2 => \_gnd_net_\,
            in3 => \N__44135\,
            lcout => \sDAC_data_RNO_26Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_5_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__37166\,
            in1 => \N__41375\,
            in2 => \N__38196\,
            in3 => \N__37100\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_5_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__37442\,
            in1 => \N__37154\,
            in2 => \N__37148\,
            in3 => \N__37046\,
            lcout => OPEN,
            ltout => \sDAC_data_2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_5_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37145\,
            in2 => \N__37130\,
            in3 => \N__37631\,
            lcout => \sDAC_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48470\,
            ce => \N__43947\,
            sr => \N__51732\
        );

    \sDAC_data_RNO_6_5_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38530\,
            in1 => \N__37106\,
            in2 => \N__38253\,
            in3 => \N__41288\,
            lcout => \sDAC_data_2_14_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_5_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__38506\,
            in1 => \N__37094\,
            in2 => \N__38195\,
            in3 => \N__37088\,
            lcout => OPEN,
            ltout => \sDAC_data_2_32_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_5_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__37073\,
            in1 => \N__38091\,
            in2 => \N__37064\,
            in3 => \N__37061\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_10Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_5_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110011101"
        )
    port map (
            in0 => \N__37334\,
            in1 => \N__37441\,
            in2 => \N__37049\,
            in3 => \N__37205\,
            lcout => \sDAC_data_2_41_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_3_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__37676\,
            in1 => \N__38177\,
            in2 => \N__41189\,
            in3 => \N__37244\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_3_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011101110"
        )
    port map (
            in0 => \N__37664\,
            in1 => \N__37455\,
            in2 => \N__37658\,
            in3 => \N__37256\,
            lcout => OPEN,
            ltout => \sDAC_data_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_3_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__37655\,
            in1 => \_gnd_net_\,
            in2 => \N__37640\,
            in3 => \N__37629\,
            lcout => \sDAC_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48473\,
            ce => \N__43948\,
            sr => \N__51720\
        );

    \sDAC_data_RNO_10_3_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__37511\,
            in1 => \N__37499\,
            in2 => \N__38232\,
            in3 => \N__37220\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_10Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_3_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__37454\,
            in1 => \N__37335\,
            in2 => \N__37271\,
            in3 => \N__37268\,
            lcout => \sDAC_data_2_41_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_3_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__38507\,
            in1 => \N__41054\,
            in2 => \N__38233\,
            in3 => \N__37250\,
            lcout => \sDAC_data_2_14_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_3_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__37238\,
            in1 => \N__38170\,
            in2 => \N__38531\,
            in3 => \N__37226\,
            lcout => \sDAC_data_2_32_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_5_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__37712\,
            in1 => \N__38579\,
            in2 => \N__38251\,
            in3 => \N__37214\,
            lcout => \sDAC_data_RNO_11Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_5_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42036\,
            in1 => \N__38597\,
            in2 => \_gnd_net_\,
            in3 => \N__37814\,
            lcout => \sDAC_data_RNO_23Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_30_6_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38573\,
            in1 => \N__41345\,
            in2 => \_gnd_net_\,
            in3 => \N__42038\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_30Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_25_6_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__38190\,
            in1 => \N__38511\,
            in2 => \N__38306\,
            in3 => \N__37682\,
            lcout => OPEN,
            ltout => \sDAC_data_2_39_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_6_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__38194\,
            in1 => \N__37856\,
            in2 => \N__37844\,
            in3 => \N__37841\,
            lcout => \sDAC_data_RNO_11Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_28_2_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47492\,
            lcout => \sDAC_mem_28Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52213\,
            ce => \N__37806\,
            sr => \N__51709\
        );

    \sDAC_data_RNO_24_5_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37739\,
            in1 => \N__37724\,
            in2 => \_gnd_net_\,
            in3 => \N__42037\,
            lcout => \sDAC_data_RNO_24Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_31_6_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__42035\,
            in1 => \N__37706\,
            in2 => \_gnd_net_\,
            in3 => \N__37694\,
            lcout => \sDAC_data_RNO_31Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_c_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42787\,
            in2 => \N__42772\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_LUT4_0_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42729\,
            in2 => \_gnd_net_\,
            in3 => \N__38672\,
            lcout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0\,
            carryout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_LUT4_0_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42678\,
            in2 => \_gnd_net_\,
            in3 => \N__38669\,
            lcout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1\,
            carryout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_3_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48303\,
            in2 => \_gnd_net_\,
            in3 => \N__38666\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2\,
            carryout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3\,
            clk => \N__48263\,
            ce => 'H',
            sr => \N__51700\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_4_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48324\,
            in2 => \_gnd_net_\,
            in3 => \N__38663\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3\,
            carryout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4\,
            clk => \N__48263\,
            ce => 'H',
            sr => \N__51700\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_5_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38653\,
            in2 => \_gnd_net_\,
            in3 => \N__38660\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48263\,
            ce => 'H',
            sr => \N__51700\
        );

    \sDAC_mem_17_0_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46293\,
            lcout => \sDAC_mem_17Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52227\,
            ce => \N__39920\,
            sr => \N__51691\
        );

    \sDAC_mem_17_1_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50880\,
            lcout => \sDAC_mem_17Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52227\,
            ce => \N__39920\,
            sr => \N__51691\
        );

    \sDAC_mem_17_2_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47511\,
            lcout => \sDAC_mem_17Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52227\,
            ce => \N__39920\,
            sr => \N__51691\
        );

    \sDAC_mem_17_3_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46907\,
            lcout => \sDAC_mem_17Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52227\,
            ce => \N__39920\,
            sr => \N__51691\
        );

    \sDAC_mem_17_4_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45611\,
            lcout => \sDAC_mem_17Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52227\,
            ce => \N__39920\,
            sr => \N__51691\
        );

    \sDAC_mem_17_5_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45107\,
            lcout => \sDAC_mem_17Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52227\,
            ce => \N__39920\,
            sr => \N__51691\
        );

    \sDAC_mem_17_6_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50527\,
            lcout => \sDAC_mem_17Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52227\,
            ce => \N__39920\,
            sr => \N__51691\
        );

    \sDAC_mem_17_7_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49874\,
            lcout => \sDAC_mem_17Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52227\,
            ce => \N__39920\,
            sr => \N__51691\
        );

    \spi_data_miso_6_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__38951\,
            in1 => \N__43767\,
            in2 => \N__38930\,
            in3 => \N__48946\,
            lcout => \spi_data_misoZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52237\,
            ce => \N__43687\,
            sr => \N__51685\
        );

    \sbuttonModeStatus_RNO_6_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38906\,
            in1 => \N__38891\,
            in2 => \N__38876\,
            in3 => \N__38858\,
            lcout => \sbuttonModeStatus_0_sqmuxa_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_7_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38834\,
            in1 => \N__38816\,
            in2 => \N__38801\,
            in3 => \N__38780\,
            lcout => \sbuttonModeStatus_0_sqmuxa_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_data_miso_0_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__38756\,
            in1 => \N__48902\,
            in2 => \N__38738\,
            in3 => \N__43768\,
            lcout => \spi_data_misoZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52249\,
            ce => \N__43686\,
            sr => \N__51680\
        );

    \spi_data_miso_4_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__38714\,
            in1 => \N__48903\,
            in2 => \N__38693\,
            in3 => \N__43769\,
            lcout => \spi_data_misoZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52249\,
            ce => \N__43686\,
            sr => \N__51680\
        );

    \reset_rpi_ibuf_RNI8S8K1_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011100000"
        )
    port map (
            in0 => \N__48899\,
            in1 => \N__39129\,
            in2 => \N__49433\,
            in3 => \N__49479\,
            lcout => \N_67_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_23_c_RNITTS3_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43445\,
            in2 => \_gnd_net_\,
            in3 => \N__43334\,
            lcout => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\,
            ltout => \un4_sacqtime_cry_23_c_RNITTSZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sSPI_MSB0LSB1_RNILL2C1_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__39165\,
            in1 => \N__39248\,
            in2 => \N__39194\,
            in3 => \N__39127\,
            lcout => \N_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sSPI_MSB0LSB1_RNIOT3R1_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001010"
        )
    port map (
            in0 => \N__39128\,
            in1 => \N__49484\,
            in2 => \N__39173\,
            in3 => \N__48897\,
            lcout => \N_70_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sSPI_MSB0LSB1_RNIGRPG4_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__48898\,
            in1 => \N__43736\,
            in2 => \N__39172\,
            in3 => \N__39130\,
            lcout => \sSPI_MSB0LSB1_RNIGRPGZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_11_15_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000010100000"
        )
    port map (
            in0 => \N__48900\,
            in1 => \N__39082\,
            in2 => \N__49432\,
            in3 => \N__49483\,
            lcout => \RAM_DATA_cl_11Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52259\,
            ce => 'H',
            sr => \N__51672\
        );

    \RAM_DATA_cl_12_15_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__39058\,
            in1 => \N__49386\,
            in2 => \N__49495\,
            in3 => \N__48901\,
            lcout => \RAM_DATA_cl_12Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52259\,
            ce => 'H',
            sr => \N__51672\
        );

    \sCounterRAM_0_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39509\,
            in1 => \N__39046\,
            in2 => \_gnd_net_\,
            in3 => \N__39032\,
            lcout => \sCounterRAMZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \sCounterRAM_cry_0\,
            clk => \N__52271\,
            ce => 'H',
            sr => \N__51664\
        );

    \sCounterRAM_1_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39505\,
            in1 => \N__39025\,
            in2 => \_gnd_net_\,
            in3 => \N__39011\,
            lcout => \sCounterRAMZ0Z_1\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_0\,
            carryout => \sCounterRAM_cry_1\,
            clk => \N__52271\,
            ce => 'H',
            sr => \N__51664\
        );

    \sCounterRAM_2_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39510\,
            in1 => \N__39601\,
            in2 => \_gnd_net_\,
            in3 => \N__39587\,
            lcout => \sCounterRAMZ0Z_2\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_1\,
            carryout => \sCounterRAM_cry_2\,
            clk => \N__52271\,
            ce => 'H',
            sr => \N__51664\
        );

    \sCounterRAM_3_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39506\,
            in1 => \N__39583\,
            in2 => \_gnd_net_\,
            in3 => \N__39569\,
            lcout => \sCounterRAMZ0Z_3\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_2\,
            carryout => \sCounterRAM_cry_3\,
            clk => \N__52271\,
            ce => 'H',
            sr => \N__51664\
        );

    \sCounterRAM_4_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39511\,
            in1 => \N__39565\,
            in2 => \_gnd_net_\,
            in3 => \N__39551\,
            lcout => \sCounterRAMZ0Z_4\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_3\,
            carryout => \sCounterRAM_cry_4\,
            clk => \N__52271\,
            ce => 'H',
            sr => \N__51664\
        );

    \sCounterRAM_5_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39507\,
            in1 => \N__39547\,
            in2 => \_gnd_net_\,
            in3 => \N__39533\,
            lcout => \sCounterRAMZ0Z_5\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_4\,
            carryout => \sCounterRAM_cry_5\,
            clk => \N__52271\,
            ce => 'H',
            sr => \N__51664\
        );

    \sCounterRAM_6_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39512\,
            in1 => \N__39529\,
            in2 => \_gnd_net_\,
            in3 => \N__39515\,
            lcout => \sCounterRAMZ0Z_6\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_5\,
            carryout => \sCounterRAM_cry_6\,
            clk => \N__52271\,
            ce => 'H',
            sr => \N__51664\
        );

    \sCounterRAM_7_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39508\,
            in1 => \N__39475\,
            in2 => \_gnd_net_\,
            in3 => \N__39482\,
            lcout => \sCounterRAMZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52271\,
            ce => 'H',
            sr => \N__51664\
        );

    \RAM_DATA_cl_6_15_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__48948\,
            in1 => \N__49413\,
            in2 => \N__39445\,
            in3 => \N__49536\,
            lcout => \RAM_DATA_cl_6Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52280\,
            ce => 'H',
            sr => \N__51659\
        );

    \RAM_DATA_cl_7_15_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__39421\,
            in1 => \N__49531\,
            in2 => \N__49440\,
            in3 => \N__48949\,
            lcout => \RAM_DATA_cl_7Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52280\,
            ce => 'H',
            sr => \N__51659\
        );

    \RAM_DATA_cl_8_15_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__48950\,
            in1 => \N__49417\,
            in2 => \N__39772\,
            in3 => \N__49537\,
            lcout => \RAM_DATA_cl_8Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52280\,
            ce => 'H',
            sr => \N__51659\
        );

    \RAM_DATA_cl_9_15_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__48951\,
            in1 => \N__49418\,
            in2 => \N__39742\,
            in3 => \N__49538\,
            lcout => \RAM_DATA_cl_9Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52280\,
            ce => 'H',
            sr => \N__51659\
        );

    \RAM_DATA_cl_15_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__39712\,
            in1 => \N__49530\,
            in2 => \N__49439\,
            in3 => \N__48947\,
            lcout => \RAM_DATA_clZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52280\,
            ce => 'H',
            sr => \N__51659\
        );

    \RAM_DATA_1_7_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \RAM_DATA_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52291\,
            ce => \N__51896\,
            sr => \N__51653\
        );

    \sDAC_mem_41_4_LC_18_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45600\,
            lcout => \sDAC_mem_41Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52260\,
            ce => \N__39806\,
            sr => \N__51814\
        );

    \sDAC_data_RNO_12_6_LC_18_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42550\,
            in1 => \N__39668\,
            in2 => \N__42263\,
            in3 => \N__39656\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_6_LC_18_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42094\,
            in1 => \N__41132\,
            in2 => \N__39644\,
            in3 => \N__44495\,
            lcout => \sDAC_data_RNO_4Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_32_5_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45101\,
            lcout => \sDAC_mem_32Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52238\,
            ce => \N__41275\,
            sr => \N__51799\
        );

    \sDAC_mem_32_7_LC_18_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_32Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52238\,
            ce => \N__41275\,
            sr => \N__51799\
        );

    \sDAC_mem_41_0_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46389\,
            lcout => \sDAC_mem_41Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52228\,
            ce => \N__39802\,
            sr => \N__51785\
        );

    \sDAC_mem_41_1_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51050\,
            lcout => \sDAC_mem_41Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52228\,
            ce => \N__39802\,
            sr => \N__51785\
        );

    \sDAC_mem_41_2_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47481\,
            lcout => \sDAC_mem_41Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52228\,
            ce => \N__39802\,
            sr => \N__51785\
        );

    \sDAC_mem_41_3_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46921\,
            lcout => \sDAC_mem_41Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52228\,
            ce => \N__39802\,
            sr => \N__51785\
        );

    \sDAC_mem_41_5_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45102\,
            lcout => \sDAC_mem_41Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52228\,
            ce => \N__39802\,
            sr => \N__51785\
        );

    \sDAC_mem_41_6_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50379\,
            lcout => \sDAC_mem_41Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52228\,
            ce => \N__39802\,
            sr => \N__51785\
        );

    \sDAC_mem_41_7_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50034\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_41Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52228\,
            ce => \N__39802\,
            sr => \N__51785\
        );

    \sAddress_RNI9IH12_9_5_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__40799\,
            in1 => \N__41026\,
            in2 => \N__41000\,
            in3 => \N__40418\,
            lcout => \sDAC_mem_9_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_1_5_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40417\,
            in1 => \N__40978\,
            in2 => \N__41027\,
            in3 => \N__40797\,
            lcout => \sDAC_mem_41_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI6VH7_6_1_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__40652\,
            in1 => \N__40546\,
            in2 => \_gnd_net_\,
            in3 => \N__40197\,
            lcout => \sAddress_RNI6VH7_6Z0Z_1\,
            ltout => \sAddress_RNI6VH7_6Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_1_3_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40416\,
            in2 => \N__41015\,
            in3 => \N__40027\,
            lcout => \sDAC_mem_25_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_4_5_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__40798\,
            in1 => \_gnd_net_\,
            in2 => \N__40999\,
            in3 => \N__40053\,
            lcout => \sDAC_mem_1_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_0_5_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__40052\,
            in1 => \N__40985\,
            in2 => \_gnd_net_\,
            in3 => \N__40800\,
            lcout => \sDAC_mem_33_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIAM2A_1_1_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__40651\,
            in1 => \N__40547\,
            in2 => \N__40429\,
            in3 => \N__40196\,
            lcout => \sAddress_RNIAM2A_1Z0Z_1\,
            ltout => \sAddress_RNIAM2A_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_0_1_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__40031\,
            in3 => \N__40026\,
            lcout => \sDAC_mem_17_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_37_0_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46374\,
            lcout => \sDAC_mem_37Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52214\,
            ce => \N__41075\,
            sr => \N__51760\
        );

    \sDAC_mem_37_1_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51042\,
            lcout => \sDAC_mem_37Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52214\,
            ce => \N__41075\,
            sr => \N__51760\
        );

    \sDAC_mem_37_2_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47484\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_37Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52214\,
            ce => \N__41075\,
            sr => \N__51760\
        );

    \sDAC_mem_37_3_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46855\,
            lcout => \sDAC_mem_37Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52214\,
            ce => \N__41075\,
            sr => \N__51760\
        );

    \sDAC_mem_37_4_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45593\,
            lcout => \sDAC_mem_37Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52214\,
            ce => \N__41075\,
            sr => \N__51760\
        );

    \sDAC_mem_37_5_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45106\,
            lcout => \sDAC_mem_37Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52214\,
            ce => \N__41075\,
            sr => \N__51760\
        );

    \sDAC_mem_37_6_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50380\,
            lcout => \sDAC_mem_37Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52214\,
            ce => \N__41075\,
            sr => \N__51760\
        );

    \sDAC_mem_37_7_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50037\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_37Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52214\,
            ce => \N__41075\,
            sr => \N__51760\
        );

    \sDAC_data_RNO_14_3_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__42188\,
            in1 => \N__41033\,
            in2 => \_gnd_net_\,
            in3 => \N__41060\,
            lcout => \sDAC_data_RNO_14Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_26_4_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42526\,
            in1 => \N__44378\,
            in2 => \_gnd_net_\,
            in3 => \N__44123\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_4_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42001\,
            in2 => \N__41048\,
            in3 => \N__41297\,
            lcout => \sDAC_data_RNO_14Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_32_0_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46344\,
            lcout => \sDAC_mem_32Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52208\,
            ce => \N__41276\,
            sr => \N__51748\
        );

    \sDAC_mem_32_1_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51063\,
            lcout => \sDAC_mem_32Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52208\,
            ce => \N__41276\,
            sr => \N__51748\
        );

    \sDAC_data_RNO_26_5_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42527\,
            in1 => \N__44369\,
            in2 => \_gnd_net_\,
            in3 => \N__44111\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_5_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42002\,
            in2 => \N__41291\,
            in3 => \N__41282\,
            lcout => \sDAC_data_RNO_14Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_32_2_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47497\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_32Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52208\,
            ce => \N__41276\,
            sr => \N__51748\
        );

    \sDAC_data_RNO_12_3_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42528\,
            in1 => \N__41213\,
            in2 => \N__42244\,
            in3 => \N__41177\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_3_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42033\,
            in1 => \N__41201\,
            in2 => \N__41192\,
            in3 => \N__44522\,
            lcout => \sDAC_data_RNO_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_4_0_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46384\,
            lcout => \sDAC_mem_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52205\,
            ce => \N__42641\,
            sr => \N__51733\
        );

    \sDAC_data_RNO_12_4_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__42566\,
            in1 => \N__41171\,
            in2 => \N__42650\,
            in3 => \N__42181\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_4_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__44513\,
            in1 => \N__42032\,
            in2 => \N__41156\,
            in3 => \N__41153\,
            lcout => \sDAC_data_RNO_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_4_1_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51077\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52205\,
            ce => \N__42641\,
            sr => \N__51733\
        );

    \sDAC_data_RNO_12_5_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__42529\,
            in1 => \N__42293\,
            in2 => \N__42245\,
            in3 => \N__42278\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_5_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__42034\,
            in1 => \N__41387\,
            in2 => \N__41378\,
            in3 => \N__44504\,
            lcout => \sDAC_data_RNO_4Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_25_5_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45115\,
            lcout => \sDAC_mem_25Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52209\,
            ce => \N__50593\,
            sr => \N__51721\
        );

    \sDAC_mem_25_2_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47507\,
            lcout => \sDAC_mem_25Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52209\,
            ce => \N__50593\,
            sr => \N__51721\
        );

    \sDAC_mem_25_3_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46923\,
            lcout => \sDAC_mem_25Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52209\,
            ce => \N__50593\,
            sr => \N__51721\
        );

    \sDAC_mem_25_4_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45607\,
            lcout => \sDAC_mem_25Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52209\,
            ce => \N__50593\,
            sr => \N__51721\
        );

    \sDAC_mem_25_0_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46317\,
            lcout => \sDAC_mem_25Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52209\,
            ce => \N__50593\,
            sr => \N__51721\
        );

    \sDAC_mem_25_6_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50381\,
            lcout => \sDAC_mem_25Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52209\,
            ce => \N__50593\,
            sr => \N__51721\
        );

    \sDAC_mem_25_7_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50063\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_25Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52209\,
            ce => \N__50593\,
            sr => \N__51721\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_0_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101110110000"
        )
    port map (
            in0 => \N__51213\,
            in1 => \N__42706\,
            in2 => \N__42791\,
            in3 => \N__42768\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48264\,
            ce => 'H',
            sr => \N__51710\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_1_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000010100"
        )
    port map (
            in0 => \N__42705\,
            in1 => \N__42746\,
            in2 => \N__42736\,
            in3 => \N__51214\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48264\,
            ce => 'H',
            sr => \N__51710\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_2_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001110001100"
        )
    port map (
            in0 => \N__51215\,
            in1 => \N__42679\,
            in2 => \N__42710\,
            in3 => \N__42689\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48264\,
            ce => 'H',
            sr => \N__51710\
        );

    \spi_slave_inst.txdata_reg_i_RNI3KQC_1_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47519\,
            in1 => \N__45782\,
            in2 => \_gnd_net_\,
            in3 => \N__48729\,
            lcout => \spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.txdata_reg_i_RNI5MQC_2_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48730\,
            in1 => \N__45674\,
            in2 => \_gnd_net_\,
            in3 => \N__45797\,
            lcout => \spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.txdata_reg_i_RNI7OQC_3_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45686\,
            in1 => \N__50558\,
            in2 => \_gnd_net_\,
            in3 => \N__48731\,
            lcout => \spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.data_in_reg_i_0_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__42659\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52221\,
            ce => \N__42830\,
            sr => \N__51701\
        );

    \spi_slave_inst.data_in_reg_i_1_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43700\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52221\,
            ce => \N__42830\,
            sr => \N__51701\
        );

    \spi_slave_inst.data_in_reg_i_2_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42854\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52221\,
            ce => \N__42830\,
            sr => \N__51701\
        );

    \spi_slave_inst.data_in_reg_i_3_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42896\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52221\,
            ce => \N__42830\,
            sr => \N__51701\
        );

    \spi_slave_inst.data_in_reg_i_4_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42845\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52221\,
            ce => \N__42830\,
            sr => \N__51701\
        );

    \spi_slave_inst.data_in_reg_i_5_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42989\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52221\,
            ce => \N__42830\,
            sr => \N__51701\
        );

    \spi_slave_inst.data_in_reg_i_6_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42836\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52221\,
            ce => \N__42830\,
            sr => \N__51701\
        );

    \spi_slave_inst.data_in_reg_i_7_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42944\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52221\,
            ce => \N__42830\,
            sr => \N__51701\
        );

    \sCounterADC_0_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46960\,
            in1 => \N__46409\,
            in2 => \_gnd_net_\,
            in3 => \N__42812\,
            lcout => \sCounterADCZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \sCounterADC_cry_0\,
            clk => \N__52229\,
            ce => \N__48960\,
            sr => \N__51692\
        );

    \sCounterADC_1_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46956\,
            in1 => \N__46421\,
            in2 => \_gnd_net_\,
            in3 => \N__42809\,
            lcout => \sCounterADCZ0Z_1\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_0\,
            carryout => \sCounterADC_cry_1\,
            clk => \N__52229\,
            ce => \N__48960\,
            sr => \N__51692\
        );

    \sCounterADC_2_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46961\,
            in1 => \N__47018\,
            in2 => \_gnd_net_\,
            in3 => \N__42806\,
            lcout => \sCounterADCZ0Z_2\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_1\,
            carryout => \sCounterADC_cry_2\,
            clk => \N__52229\,
            ce => \N__48960\,
            sr => \N__51692\
        );

    \sCounterADC_3_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46957\,
            in1 => \N__47000\,
            in2 => \_gnd_net_\,
            in3 => \N__43082\,
            lcout => \sCounterADCZ0Z_3\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_2\,
            carryout => \sCounterADC_cry_3\,
            clk => \N__52229\,
            ce => \N__48960\,
            sr => \N__51692\
        );

    \sCounterADC_4_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46962\,
            in1 => \N__43069\,
            in2 => \_gnd_net_\,
            in3 => \N__43055\,
            lcout => \sCounterADCZ0Z_4\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_3\,
            carryout => \sCounterADC_cry_4\,
            clk => \N__52229\,
            ce => \N__48960\,
            sr => \N__51692\
        );

    \sCounterADC_5_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46958\,
            in1 => \N__43042\,
            in2 => \_gnd_net_\,
            in3 => \N__43028\,
            lcout => \sCounterADCZ0Z_5\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_4\,
            carryout => \sCounterADC_cry_5\,
            clk => \N__52229\,
            ce => \N__48960\,
            sr => \N__51692\
        );

    \sCounterADC_6_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46963\,
            in1 => \N__45844\,
            in2 => \_gnd_net_\,
            in3 => \N__43025\,
            lcout => \sCounterADCZ0Z_6\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_5\,
            carryout => \sCounterADC_cry_6\,
            clk => \N__52229\,
            ce => \N__48960\,
            sr => \N__51692\
        );

    \sCounterADC_7_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__46959\,
            in1 => \N__45857\,
            in2 => \_gnd_net_\,
            in3 => \N__43022\,
            lcout => \sCounterADCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52229\,
            ce => \N__48960\,
            sr => \N__51692\
        );

    \spi_data_miso_5_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__43019\,
            in1 => \N__43001\,
            in2 => \N__43772\,
            in3 => \N__48910\,
            lcout => \spi_data_misoZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52239\,
            ce => \N__43691\,
            sr => \N__51686\
        );

    \spi_data_miso_7_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__48911\,
            in1 => \N__42980\,
            in2 => \N__42968\,
            in3 => \N__43766\,
            lcout => \spi_data_misoZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52239\,
            ce => \N__43691\,
            sr => \N__51686\
        );

    \spi_data_miso_3_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__48909\,
            in1 => \N__42935\,
            in2 => \N__42917\,
            in3 => \N__43765\,
            lcout => \spi_data_misoZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52239\,
            ce => \N__43691\,
            sr => \N__51686\
        );

    \spi_data_miso_2_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__42887\,
            in1 => \N__42872\,
            in2 => \N__43771\,
            in3 => \N__48908\,
            lcout => \spi_data_misoZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52239\,
            ce => \N__43691\,
            sr => \N__51686\
        );

    \spi_data_miso_1_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__43808\,
            in1 => \N__43787\,
            in2 => \N__43770\,
            in3 => \N__48907\,
            lcout => \spi_data_misoZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52239\,
            ce => \N__43691\,
            sr => \N__51686\
        );

    \sRAM_ADD_8_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__43347\,
            in1 => \N__43661\,
            in2 => \N__43634\,
            in3 => \N__43468\,
            lcout => \RAM_ADD_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52250\,
            ce => \N__43225\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_4_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__43346\,
            in1 => \N__43589\,
            in2 => \N__43562\,
            in3 => \N__43467\,
            lcout => \RAM_ADD_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52250\,
            ce => \N__43225\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_3_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__43520\,
            in1 => \N__43466\,
            in2 => \N__43376\,
            in3 => \N__43345\,
            lcout => \RAM_ADD_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52250\,
            ce => \N__43225\,
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_13_15_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__43183\,
            in1 => \N__49527\,
            in2 => \N__49436\,
            in3 => \N__48930\,
            lcout => \RAM_DATA_cl_13Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52261\,
            ce => 'H',
            sr => \N__51673\
        );

    \RAM_DATA_cl_14_15_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__48931\,
            in1 => \N__49400\,
            in2 => \N__43159\,
            in3 => \N__49532\,
            lcout => \RAM_DATA_cl_14Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52261\,
            ce => 'H',
            sr => \N__51673\
        );

    \RAM_DATA_cl_15_15_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__43126\,
            in1 => \N__49528\,
            in2 => \N__49437\,
            in3 => \N__48932\,
            lcout => \RAM_DATA_cl_15Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52261\,
            ce => 'H',
            sr => \N__51673\
        );

    \RAM_DATA_cl_1_15_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__48933\,
            in1 => \N__49404\,
            in2 => \N__43099\,
            in3 => \N__49533\,
            lcout => \RAM_DATA_cl_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52261\,
            ce => 'H',
            sr => \N__51673\
        );

    \RAM_DATA_cl_10_15_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__44056\,
            in1 => \N__49526\,
            in2 => \N__49435\,
            in3 => \N__48929\,
            lcout => \RAM_DATA_cl_10Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52261\,
            ce => 'H',
            sr => \N__51673\
        );

    \RAM_DATA_cl_3_15_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__48935\,
            in1 => \N__49406\,
            in2 => \N__44032\,
            in3 => \N__49535\,
            lcout => \RAM_DATA_cl_3Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52261\,
            ce => 'H',
            sr => \N__51673\
        );

    \RAM_DATA_cl_4_15_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__43999\,
            in1 => \N__49529\,
            in2 => \N__49438\,
            in3 => \N__48936\,
            lcout => \RAM_DATA_cl_4Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52261\,
            ce => 'H',
            sr => \N__51673\
        );

    \RAM_DATA_cl_2_15_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000010001000"
        )
    port map (
            in0 => \N__48934\,
            in1 => \N__49405\,
            in2 => \N__43975\,
            in3 => \N__49534\,
            lcout => \RAM_DATA_cl_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52261\,
            ce => 'H',
            sr => \N__51673\
        );

    \sDAC_data_2_LC_19_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48454\,
            ce => \N__43955\,
            sr => \N__51826\
        );

    \spi_master_inst.spi_data_path_u1.data_in_2_LC_19_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43916\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48458\,
            ce => \N__43907\,
            sr => \N__51824\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_2_LC_19_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43853\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48460\,
            ce => 'H',
            sr => \N__51820\
        );

    \sDAC_mem_7_2_LC_19_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47329\,
            lcout => \sDAC_mem_7Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52240\,
            ce => \N__44285\,
            sr => \N__51815\
        );

    \sDAC_mem_7_3_LC_19_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46789\,
            lcout => \sDAC_mem_7Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52240\,
            ce => \N__44285\,
            sr => \N__51815\
        );

    \sDAC_mem_7_4_LC_19_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45359\,
            lcout => \sDAC_mem_7Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52240\,
            ce => \N__44285\,
            sr => \N__51815\
        );

    \sDAC_mem_7_6_LC_19_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50374\,
            lcout => \sDAC_mem_7Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52240\,
            ce => \N__44285\,
            sr => \N__51815\
        );

    \sDAC_mem_3_7_LC_19_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50033\,
            lcout => \sDAC_mem_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52230\,
            ce => \N__44239\,
            sr => \N__51808\
        );

    \sDAC_mem_1_0_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46390\,
            lcout => \sDAC_mem_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52222\,
            ce => \N__44402\,
            sr => \N__51800\
        );

    \sDAC_mem_1_1_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51051\,
            lcout => \sDAC_mem_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52222\,
            ce => \N__44402\,
            sr => \N__51800\
        );

    \sDAC_mem_1_2_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47482\,
            lcout => \sDAC_mem_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52222\,
            ce => \N__44402\,
            sr => \N__51800\
        );

    \sDAC_mem_1_3_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46922\,
            lcout => \sDAC_mem_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52222\,
            ce => \N__44402\,
            sr => \N__51800\
        );

    \sDAC_mem_1_4_LC_19_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45561\,
            lcout => \sDAC_mem_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52222\,
            ce => \N__44402\,
            sr => \N__51800\
        );

    \sDAC_mem_1_5_LC_19_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45064\,
            lcout => \sDAC_mem_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52222\,
            ce => \N__44402\,
            sr => \N__51800\
        );

    \sDAC_mem_1_6_LC_19_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50464\,
            lcout => \sDAC_mem_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52222\,
            ce => \N__44402\,
            sr => \N__51800\
        );

    \sDAC_mem_1_7_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50035\,
            lcout => \sDAC_mem_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52222\,
            ce => \N__44402\,
            sr => \N__51800\
        );

    \sDAC_mem_33_0_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46382\,
            lcout => \sDAC_mem_33Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52215\,
            ce => \N__44531\,
            sr => \N__51786\
        );

    \sDAC_mem_33_1_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51076\,
            lcout => \sDAC_mem_33Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52215\,
            ce => \N__44531\,
            sr => \N__51786\
        );

    \sDAC_mem_33_2_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47483\,
            lcout => \sDAC_mem_33Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52215\,
            ce => \N__44531\,
            sr => \N__51786\
        );

    \sDAC_mem_33_3_LC_19_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46857\,
            lcout => \sDAC_mem_33Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52215\,
            ce => \N__44531\,
            sr => \N__51786\
        );

    \sDAC_mem_33_4_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45562\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_33Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52215\,
            ce => \N__44531\,
            sr => \N__51786\
        );

    \sDAC_mem_33_5_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45065\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_33Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52215\,
            ce => \N__44531\,
            sr => \N__51786\
        );

    \sDAC_mem_33_6_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50465\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_33Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52215\,
            ce => \N__44531\,
            sr => \N__51786\
        );

    \sDAC_mem_33_7_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50036\,
            lcout => \sDAC_mem_33Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52215\,
            ce => \N__44531\,
            sr => \N__51786\
        );

    \sDAC_mem_5_0_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46383\,
            lcout => \sDAC_mem_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52210\,
            ce => \N__44435\,
            sr => \N__51773\
        );

    \sDAC_mem_5_1_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51043\,
            lcout => \sDAC_mem_5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52210\,
            ce => \N__44435\,
            sr => \N__51773\
        );

    \sDAC_mem_5_2_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47485\,
            lcout => \sDAC_mem_5Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52210\,
            ce => \N__44435\,
            sr => \N__51773\
        );

    \sDAC_mem_5_3_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46856\,
            lcout => \sDAC_mem_5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52210\,
            ce => \N__44435\,
            sr => \N__51773\
        );

    \sDAC_mem_5_4_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__45563\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52210\,
            ce => \N__44435\,
            sr => \N__51773\
        );

    \sDAC_mem_5_5_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45066\,
            lcout => \sDAC_mem_5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52210\,
            ce => \N__44435\,
            sr => \N__51773\
        );

    \sDAC_mem_5_6_LC_19_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50466\,
            lcout => \sDAC_mem_5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52210\,
            ce => \N__44435\,
            sr => \N__51773\
        );

    \sDAC_mem_5_7_LC_19_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50061\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_5Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52210\,
            ce => \N__44435\,
            sr => \N__51773\
        );

    \sDAC_mem_13_0_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46345\,
            lcout => \sDAC_mem_13Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52206\,
            ce => \N__44585\,
            sr => \N__51761\
        );

    \sDAC_mem_13_1_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51064\,
            lcout => \sDAC_mem_13Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52206\,
            ce => \N__44585\,
            sr => \N__51761\
        );

    \sDAC_mem_13_2_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47498\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_13Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52206\,
            ce => \N__44585\,
            sr => \N__51761\
        );

    \sDAC_mem_13_3_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46906\,
            lcout => \sDAC_mem_13Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52206\,
            ce => \N__44585\,
            sr => \N__51761\
        );

    \sDAC_mem_13_4_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45602\,
            lcout => \sDAC_mem_13Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52206\,
            ce => \N__44585\,
            sr => \N__51761\
        );

    \sDAC_mem_13_5_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45105\,
            lcout => \sDAC_mem_13Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52206\,
            ce => \N__44585\,
            sr => \N__51761\
        );

    \sDAC_mem_13_6_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50526\,
            lcout => \sDAC_mem_13Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52206\,
            ce => \N__44585\,
            sr => \N__51761\
        );

    \sDAC_mem_13_7_LC_19_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50062\,
            lcout => \sDAC_mem_13Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52206\,
            ce => \N__44585\,
            sr => \N__51761\
        );

    \spi_slave_inst.tx_ready_i_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__51191\,
            in1 => \N__44557\,
            in2 => \N__49390\,
            in3 => \N__51089\,
            lcout => \spi_slave_inst.tx_ready_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52203\,
            ce => 'H',
            sr => \N__51749\
        );

    \spi_slave_inst.txdata_reg_i_4_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45824\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52207\,
            ce => 'H',
            sr => \N__51734\
        );

    \spi_slave_inst.txdata_reg_i_0_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45815\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52207\,
            ce => 'H',
            sr => \N__51734\
        );

    \spi_slave_inst.txdata_reg_i_2_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45806\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52207\,
            ce => 'H',
            sr => \N__51734\
        );

    \spi_slave_inst.txdata_reg_i_1_LC_19_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45791\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52207\,
            ce => 'H',
            sr => \N__51734\
        );

    \button_debounce_counter_1_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__45744\,
            in1 => \N__49240\,
            in2 => \_gnd_net_\,
            in3 => \N__45771\,
            lcout => \button_debounce_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48487\,
            ce => 'H',
            sr => \N__45718\
        );

    \button_debounce_counter_0_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49145\,
            in2 => \_gnd_net_\,
            in3 => \N__45743\,
            lcout => \button_debounce_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48487\,
            ce => 'H',
            sr => \N__45718\
        );

    \spi_slave_inst.txdata_reg_i_3_LC_19_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45692\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52216\,
            ce => 'H',
            sr => \N__51711\
        );

    \spi_slave_inst.txdata_reg_i_6_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45680\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52216\,
            ce => 'H',
            sr => \N__51711\
        );

    \spi_slave_inst.txdata_reg_i_5_LC_19_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47525\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52216\,
            ce => 'H',
            sr => \N__51711\
        );

    \sEEADC_freq_2_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47513\,
            lcout => \sEEADC_freqZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52231\,
            ce => \N__49576\,
            sr => \_gnd_net_\
        );

    \sEEADC_freq_RNI4KIA1_2_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__47017\,
            in1 => \N__47006\,
            in2 => \N__46430\,
            in3 => \N__46999\,
            lcout => OPEN,
            ltout => \un11_sacqtime_NE_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEADC_freq_RNI01BA5_0_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46988\,
            in1 => \N__45830\,
            in2 => \N__46973\,
            in3 => \N__46397\,
            lcout => \un11_sacqtime_NE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEADC_freq_3_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46765\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEADC_freqZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52231\,
            ce => \N__49576\,
            sr => \_gnd_net_\
        );

    \sEEADC_freq_RNISBIA1_0_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__45872\,
            in1 => \N__46420\,
            in2 => \N__45866\,
            in3 => \N__46408\,
            lcout => \un11_sacqtime_NE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEADC_freq_0_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46316\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEADC_freqZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52231\,
            ce => \N__49576\,
            sr => \_gnd_net_\
        );

    \sEEADC_freq_1_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51019\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEADC_freqZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52231\,
            ce => \N__49576\,
            sr => \_gnd_net_\
        );

    \sEEADC_freq_RNIK4JA1_6_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__50072\,
            in1 => \N__45856\,
            in2 => \N__45845\,
            in3 => \N__49586\,
            lcout => \un11_sacqtime_NE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_1_8_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47717\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RAM_DATA_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52241\,
            ce => \N__51882\,
            sr => \N__51687\
        );

    \RAM_DATA_1_9_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47678\,
            lcout => \RAM_DATA_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52241\,
            ce => \N__51882\,
            sr => \N__51687\
        );

    \RAM_DATA_1_12_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47636\,
            lcout => \RAM_DATA_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52241\,
            ce => \N__51882\,
            sr => \N__51687\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ00Q2_0_LC_20_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48052\,
            in2 => \_gnd_net_\,
            in3 => \N__47782\,
            lcout => spi_miso_ft_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_8_LC_20_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47582\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48463\,
            ce => 'H',
            sr => \N__51825\
        );

    \sCounterDAC_0_LC_20_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48126\,
            lcout => \sCounterDACZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48463\,
            ce => 'H',
            sr => \N__51825\
        );

    \spi_slave_inst.spi_cs_LC_20_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__47928\,
            in1 => \N__48051\,
            in2 => \_gnd_net_\,
            in3 => \N__47887\,
            lcout => \spi_slave_inst.spi_csZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_spi_start_LC_20_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__48554\,
            in1 => \N__48539\,
            in2 => \N__47545\,
            in3 => \N__48140\,
            lcout => \sDAC_spi_startZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48466\,
            ce => 'H',
            sr => \N__51816\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNIOASC_5_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__51263\,
            in1 => \N__51242\,
            in2 => \N__48689\,
            in3 => \N__48772\,
            lcout => OPEN,
            ltout => \spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNI1DAJ_1_LC_20_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48717\,
            in2 => \N__48059\,
            in3 => \N__48753\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_i6\,
            ltout => \spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1_1_LC_20_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__48056\,
            in1 => \N__47929\,
            in2 => \N__47906\,
            in3 => \N__47888\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNIUCSS_1_LC_20_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47831\,
            in1 => \N__47816\,
            in2 => \_gnd_net_\,
            in3 => \N__48755\,
            lcout => OPEN,
            ltout => \spi_slave_inst.N_1393_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNIA0LM2_0_LC_20_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__47723\,
            in1 => \N__51178\,
            in2 => \N__47801\,
            in3 => \N__48773\,
            lcout => spi_miso,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.txdata_reg_i_RNI1IQC_0_LC_20_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47765\,
            in1 => \N__47753\,
            in2 => \_gnd_net_\,
            in3 => \N__48718\,
            lcout => OPEN,
            ltout => \spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ8SS_1_LC_20_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__48754\,
            in1 => \_gnd_net_\,
            in2 => \N__47741\,
            in3 => \N__47738\,
            lcout => \spi_slave_inst.N_1396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_RNI9VC2_3_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48668\,
            in2 => \_gnd_net_\,
            in3 => \N__48127\,
            lcout => m15_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_1_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__48131\,
            in1 => \_gnd_net_\,
            in2 => \N__48097\,
            in3 => \_gnd_net_\,
            lcout => \sCounterDACZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48477\,
            ce => 'H',
            sr => \N__51787\
        );

    \sCounterDAC_RNIHIJ3_1_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__48637\,
            in1 => \N__48090\,
            in2 => \_gnd_net_\,
            in3 => \N__48665\,
            lcout => m8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_RNI4HQ4_9_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__48568\,
            in1 => \N__48073\,
            in2 => \N__48509\,
            in3 => \N__48591\,
            lcout => \N_23_mux\,
            ltout => \N_23_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_RNIFI77_1_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010000"
        )
    port map (
            in0 => \N__48636\,
            in1 => \N__48089\,
            in2 => \N__48191\,
            in3 => \_gnd_net_\,
            lcout => \N_25_mux\,
            ltout => \N_25_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_RNIBR1C_5_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48533\,
            in1 => \N__48611\,
            in2 => \N__48188\,
            in3 => \N__48185\,
            lcout => op_eq_scounterdac10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_RNI05RA_5_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__48161\,
            in1 => \N__48155\,
            in2 => \N__48619\,
            in3 => \N__48129\,
            lcout => \N_30_mux\,
            ltout => \N_30_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_6_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__48534\,
            in1 => \N__48578\,
            in2 => \N__48149\,
            in3 => \N__48592\,
            lcout => \sCounterDACZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48477\,
            ce => 'H',
            sr => \N__51787\
        );

    \sDAC_spi_start_RNO_0_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__48667\,
            in1 => \N__48130\,
            in2 => \N__48620\,
            in3 => \N__48146\,
            lcout => \N_32_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_scounterdac_cry_1_c_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48128\,
            in2 => \N__48098\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_20_10_0_\,
            carryout => un2_scounterdac_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_2_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48074\,
            in2 => \_gnd_net_\,
            in3 => \N__48062\,
            lcout => \sCounterDACZ0Z_2\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_1,
            carryout => un2_scounterdac_cry_2,
            clk => \N__48481\,
            ce => 'H',
            sr => \N__51774\
        );

    \sCounterDAC_3_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48666\,
            in2 => \_gnd_net_\,
            in3 => \N__48641\,
            lcout => \sCounterDACZ0Z_3\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_2,
            carryout => un2_scounterdac_cry_3,
            clk => \N__48481\,
            ce => 'H',
            sr => \N__51774\
        );

    \sCounterDAC_4_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48638\,
            in2 => \_gnd_net_\,
            in3 => \N__48623\,
            lcout => \sCounterDACZ0Z_4\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_3,
            carryout => un2_scounterdac_cry_4,
            clk => \N__48481\,
            ce => 'H',
            sr => \N__51774\
        );

    \sCounterDAC_5_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48618\,
            in2 => \_gnd_net_\,
            in3 => \N__48596\,
            lcout => \sCounterDACZ0Z_5\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_4,
            carryout => un2_scounterdac_cry_5,
            clk => \N__48481\,
            ce => 'H',
            sr => \N__51774\
        );

    \un2_scounterdac_cry_5_THRU_LUT4_0_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48593\,
            in2 => \_gnd_net_\,
            in3 => \N__48572\,
            lcout => \un2_scounterdac_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_5,
            carryout => un2_scounterdac_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_7_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48569\,
            in2 => \_gnd_net_\,
            in3 => \N__48557\,
            lcout => \sCounterDACZ0Z_7\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_6,
            carryout => un2_scounterdac_cry_7,
            clk => \N__48481\,
            ce => 'H',
            sr => \N__51774\
        );

    \sCounterDAC_8_LC_20_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001101000100"
        )
    port map (
            in0 => \N__48553\,
            in1 => \N__48535\,
            in2 => \_gnd_net_\,
            in3 => \N__48515\,
            lcout => \sCounterDACZ0Z_8\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_7,
            carryout => un2_scounterdac_cry_8,
            clk => \N__48481\,
            ce => 'H',
            sr => \N__51774\
        );

    \sCounterDAC_9_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48505\,
            in2 => \_gnd_net_\,
            in3 => \N__48512\,
            lcout => \sCounterDACZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48484\,
            ce => 'H',
            sr => \N__51762\
        );

    \spi_slave_inst.rx_done_pos_sclk_i_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__48341\,
            in1 => \N__48328\,
            in2 => \_gnd_net_\,
            in3 => \N__48305\,
            lcout => \spi_slave_inst.rx_done_pos_sclk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48266\,
            ce => \N__48232\,
            sr => \N__51735\
        );

    \spi_slave_inst.txdata_reg_i_7_LC_20_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50570\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52217\,
            ce => 'H',
            sr => \N__51712\
        );

    \sEEADC_freq_6_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50480\,
            lcout => \sEEADC_freqZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52223\,
            ce => \N__49580\,
            sr => \_gnd_net_\
        );

    \sEEADC_freq_7_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50048\,
            lcout => \sEEADC_freqZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52223\,
            ce => \N__49580\,
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_5_15_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__48802\,
            in1 => \N__49494\,
            in2 => \N__49434\,
            in3 => \N__48956\,
            lcout => \RAM_DATA_cl_5Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52232\,
            ce => 'H',
            sr => \N__51693\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_0_LC_22_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__51143\,
            in1 => \N__48771\,
            in2 => \N__48791\,
            in3 => \N__48790\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_22_7_0_\,
            carryout => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0\,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51821\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_1_LC_22_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__51145\,
            in1 => \N__48752\,
            in2 => \_gnd_net_\,
            in3 => \N__48734\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0\,
            carryout => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1\,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51821\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_2_LC_22_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__51144\,
            in1 => \N__48713\,
            in2 => \_gnd_net_\,
            in3 => \N__48692\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1\,
            carryout => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2\,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51821\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_3_LC_22_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48685\,
            in2 => \_gnd_net_\,
            in3 => \N__48671\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2\,
            carryout => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3\,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51821\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_4_LC_22_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51262\,
            in2 => \_gnd_net_\,
            in3 => \N__51248\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3\,
            carryout => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4\,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51821\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_5_LC_22_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51241\,
            in2 => \_gnd_net_\,
            in3 => \N__51245\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51821\
        );

    \spi_slave_inst.tx_done_neg_sclk_i_LC_22_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__51197\,
            in1 => \N__51124\,
            in2 => \_gnd_net_\,
            in3 => \N__51146\,
            lcout => \spi_slave_inst.tx_done_neg_sclk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__51821\
        );

    \spi_slave_inst.tx_done_reg1_i_LC_22_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51125\,
            lcout => \spi_slave_inst.tx_done_reg1_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52204\,
            ce => 'H',
            sr => \N__51817\
        );

    \spi_slave_inst.tx_done_reg2_i_LC_22_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51113\,
            lcout => \spi_slave_inst.tx_done_reg2_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52202\,
            ce => 'H',
            sr => \N__51809\
        );

    \spi_slave_inst.tx_done_reg3_i_LC_22_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51101\,
            lcout => \spi_slave_inst.tx_done_reg3_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52202\,
            ce => 'H',
            sr => \N__51809\
        );

    \CONSTANT_ONE_LUT4_LC_22_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_ready_i_RNO_0_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51107\,
            in2 => \_gnd_net_\,
            in3 => \N__51100\,
            lcout => \spi_slave_inst.un4_tx_done_reg2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_25_1_LC_22_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51029\,
            lcout => \sDAC_mem_25Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52201\,
            ce => \N__50594\,
            sr => \N__51775\
        );

    \RAM_DATA_1_15_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52408\,
            lcout => \RAM_DATA_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52211\,
            ce => \N__51894\,
            sr => \N__51722\
        );
end \INTERFACE\;
