-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 13 2018 07:24:19

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MATTY_MAIN_VHDL" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MATTY_MAIN_VHDL
entity MATTY_MAIN_VHDL is
port (
    RAM_DATA : inout std_logic_vector(15 downto 0);
    RAM_ADD : out std_logic_vector(18 downto 0);
    spi_sclk_ft : in std_logic;
    button_trig : in std_logic;
    ADC9 : in std_logic;
    spi_cs_ft : in std_logic;
    poff : out std_logic;
    RAM_nOE : out std_logic;
    ADC0 : in std_logic;
    spi_mosi_flash : out std_logic;
    spi_miso_flash : in std_logic;
    trig_ft : in std_logic;
    spi_miso_rpi : out std_logic;
    RAM_nWE : out std_logic;
    DAC_cs : out std_logic;
    ADC6 : in std_logic;
    spi_select : in std_logic;
    clk : in std_logic;
    ADC4 : in std_logic;
    trig_rpi : in std_logic;
    top_tour2 : in std_logic;
    spi_cs_rpi : in std_logic;
    DAC_sclk : out std_logic;
    ADC_clk : out std_logic;
    ADC3 : in std_logic;
    trig_ext : in std_logic;
    spi_mosi_rpi : in std_logic;
    spi_mosi_ft : in std_logic;
    cs_rpi2flash : in std_logic;
    spi_cs_flash : out std_logic;
    pon : out std_logic;
    RAM_nCE : out std_logic;
    LED3 : out std_logic;
    ADC1 : in std_logic;
    reset_rpi : in std_logic;
    RAM_nLB : out std_logic;
    LED_MODE : out std_logic;
    ADC8 : in std_logic;
    spi_sclk_rpi : in std_logic;
    ADC7 : in std_logic;
    top_tour1 : in std_logic;
    spi_miso_ft : out std_logic;
    button_mode : in std_logic;
    DAC_mosi : out std_logic;
    ADC5 : in std_logic;
    reset_ft : in std_logic;
    LED_ACQ : out std_logic;
    spi_sclk_flash : out std_logic;
    reset_alim : in std_logic;
    RAM_nUB : out std_logic;
    ADC2 : in std_logic);
end MATTY_MAIN_VHDL;

-- Architecture of MATTY_MAIN_VHDL
-- View name is \INTERFACE\
architecture \INTERFACE\ of MATTY_MAIN_VHDL is

signal \N__54196\ : std_logic;
signal \N__54195\ : std_logic;
signal \N__54194\ : std_logic;
signal \N__54187\ : std_logic;
signal \N__54186\ : std_logic;
signal \N__54185\ : std_logic;
signal \N__54178\ : std_logic;
signal \N__54177\ : std_logic;
signal \N__54176\ : std_logic;
signal \N__54169\ : std_logic;
signal \N__54168\ : std_logic;
signal \N__54167\ : std_logic;
signal \N__54160\ : std_logic;
signal \N__54159\ : std_logic;
signal \N__54158\ : std_logic;
signal \N__54151\ : std_logic;
signal \N__54150\ : std_logic;
signal \N__54149\ : std_logic;
signal \N__54142\ : std_logic;
signal \N__54141\ : std_logic;
signal \N__54140\ : std_logic;
signal \N__54133\ : std_logic;
signal \N__54132\ : std_logic;
signal \N__54131\ : std_logic;
signal \N__54124\ : std_logic;
signal \N__54123\ : std_logic;
signal \N__54122\ : std_logic;
signal \N__54115\ : std_logic;
signal \N__54114\ : std_logic;
signal \N__54113\ : std_logic;
signal \N__54106\ : std_logic;
signal \N__54105\ : std_logic;
signal \N__54104\ : std_logic;
signal \N__54097\ : std_logic;
signal \N__54096\ : std_logic;
signal \N__54095\ : std_logic;
signal \N__54088\ : std_logic;
signal \N__54087\ : std_logic;
signal \N__54086\ : std_logic;
signal \N__54079\ : std_logic;
signal \N__54078\ : std_logic;
signal \N__54077\ : std_logic;
signal \N__54070\ : std_logic;
signal \N__54069\ : std_logic;
signal \N__54068\ : std_logic;
signal \N__54061\ : std_logic;
signal \N__54060\ : std_logic;
signal \N__54059\ : std_logic;
signal \N__54052\ : std_logic;
signal \N__54051\ : std_logic;
signal \N__54050\ : std_logic;
signal \N__54043\ : std_logic;
signal \N__54042\ : std_logic;
signal \N__54041\ : std_logic;
signal \N__54034\ : std_logic;
signal \N__54033\ : std_logic;
signal \N__54032\ : std_logic;
signal \N__54025\ : std_logic;
signal \N__54024\ : std_logic;
signal \N__54023\ : std_logic;
signal \N__54016\ : std_logic;
signal \N__54015\ : std_logic;
signal \N__54014\ : std_logic;
signal \N__54007\ : std_logic;
signal \N__54006\ : std_logic;
signal \N__54005\ : std_logic;
signal \N__53998\ : std_logic;
signal \N__53997\ : std_logic;
signal \N__53996\ : std_logic;
signal \N__53989\ : std_logic;
signal \N__53988\ : std_logic;
signal \N__53987\ : std_logic;
signal \N__53980\ : std_logic;
signal \N__53979\ : std_logic;
signal \N__53978\ : std_logic;
signal \N__53971\ : std_logic;
signal \N__53970\ : std_logic;
signal \N__53969\ : std_logic;
signal \N__53962\ : std_logic;
signal \N__53961\ : std_logic;
signal \N__53960\ : std_logic;
signal \N__53953\ : std_logic;
signal \N__53952\ : std_logic;
signal \N__53951\ : std_logic;
signal \N__53944\ : std_logic;
signal \N__53943\ : std_logic;
signal \N__53942\ : std_logic;
signal \N__53935\ : std_logic;
signal \N__53934\ : std_logic;
signal \N__53933\ : std_logic;
signal \N__53926\ : std_logic;
signal \N__53925\ : std_logic;
signal \N__53924\ : std_logic;
signal \N__53917\ : std_logic;
signal \N__53916\ : std_logic;
signal \N__53915\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53907\ : std_logic;
signal \N__53906\ : std_logic;
signal \N__53899\ : std_logic;
signal \N__53898\ : std_logic;
signal \N__53897\ : std_logic;
signal \N__53890\ : std_logic;
signal \N__53889\ : std_logic;
signal \N__53888\ : std_logic;
signal \N__53881\ : std_logic;
signal \N__53880\ : std_logic;
signal \N__53879\ : std_logic;
signal \N__53872\ : std_logic;
signal \N__53871\ : std_logic;
signal \N__53870\ : std_logic;
signal \N__53863\ : std_logic;
signal \N__53862\ : std_logic;
signal \N__53861\ : std_logic;
signal \N__53854\ : std_logic;
signal \N__53853\ : std_logic;
signal \N__53852\ : std_logic;
signal \N__53845\ : std_logic;
signal \N__53844\ : std_logic;
signal \N__53843\ : std_logic;
signal \N__53836\ : std_logic;
signal \N__53835\ : std_logic;
signal \N__53834\ : std_logic;
signal \N__53827\ : std_logic;
signal \N__53826\ : std_logic;
signal \N__53825\ : std_logic;
signal \N__53818\ : std_logic;
signal \N__53817\ : std_logic;
signal \N__53816\ : std_logic;
signal \N__53809\ : std_logic;
signal \N__53808\ : std_logic;
signal \N__53807\ : std_logic;
signal \N__53800\ : std_logic;
signal \N__53799\ : std_logic;
signal \N__53798\ : std_logic;
signal \N__53791\ : std_logic;
signal \N__53790\ : std_logic;
signal \N__53789\ : std_logic;
signal \N__53782\ : std_logic;
signal \N__53781\ : std_logic;
signal \N__53780\ : std_logic;
signal \N__53773\ : std_logic;
signal \N__53772\ : std_logic;
signal \N__53771\ : std_logic;
signal \N__53764\ : std_logic;
signal \N__53763\ : std_logic;
signal \N__53762\ : std_logic;
signal \N__53755\ : std_logic;
signal \N__53754\ : std_logic;
signal \N__53753\ : std_logic;
signal \N__53746\ : std_logic;
signal \N__53745\ : std_logic;
signal \N__53744\ : std_logic;
signal \N__53737\ : std_logic;
signal \N__53736\ : std_logic;
signal \N__53735\ : std_logic;
signal \N__53728\ : std_logic;
signal \N__53727\ : std_logic;
signal \N__53726\ : std_logic;
signal \N__53719\ : std_logic;
signal \N__53718\ : std_logic;
signal \N__53717\ : std_logic;
signal \N__53710\ : std_logic;
signal \N__53709\ : std_logic;
signal \N__53708\ : std_logic;
signal \N__53701\ : std_logic;
signal \N__53700\ : std_logic;
signal \N__53699\ : std_logic;
signal \N__53692\ : std_logic;
signal \N__53691\ : std_logic;
signal \N__53690\ : std_logic;
signal \N__53683\ : std_logic;
signal \N__53682\ : std_logic;
signal \N__53681\ : std_logic;
signal \N__53674\ : std_logic;
signal \N__53673\ : std_logic;
signal \N__53672\ : std_logic;
signal \N__53665\ : std_logic;
signal \N__53664\ : std_logic;
signal \N__53663\ : std_logic;
signal \N__53656\ : std_logic;
signal \N__53655\ : std_logic;
signal \N__53654\ : std_logic;
signal \N__53647\ : std_logic;
signal \N__53646\ : std_logic;
signal \N__53645\ : std_logic;
signal \N__53638\ : std_logic;
signal \N__53637\ : std_logic;
signal \N__53636\ : std_logic;
signal \N__53629\ : std_logic;
signal \N__53628\ : std_logic;
signal \N__53627\ : std_logic;
signal \N__53620\ : std_logic;
signal \N__53619\ : std_logic;
signal \N__53618\ : std_logic;
signal \N__53611\ : std_logic;
signal \N__53610\ : std_logic;
signal \N__53609\ : std_logic;
signal \N__53602\ : std_logic;
signal \N__53601\ : std_logic;
signal \N__53600\ : std_logic;
signal \N__53593\ : std_logic;
signal \N__53592\ : std_logic;
signal \N__53591\ : std_logic;
signal \N__53584\ : std_logic;
signal \N__53583\ : std_logic;
signal \N__53582\ : std_logic;
signal \N__53575\ : std_logic;
signal \N__53574\ : std_logic;
signal \N__53573\ : std_logic;
signal \N__53566\ : std_logic;
signal \N__53565\ : std_logic;
signal \N__53564\ : std_logic;
signal \N__53557\ : std_logic;
signal \N__53556\ : std_logic;
signal \N__53555\ : std_logic;
signal \N__53548\ : std_logic;
signal \N__53547\ : std_logic;
signal \N__53546\ : std_logic;
signal \N__53539\ : std_logic;
signal \N__53538\ : std_logic;
signal \N__53537\ : std_logic;
signal \N__53530\ : std_logic;
signal \N__53529\ : std_logic;
signal \N__53528\ : std_logic;
signal \N__53521\ : std_logic;
signal \N__53520\ : std_logic;
signal \N__53519\ : std_logic;
signal \N__53512\ : std_logic;
signal \N__53511\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53503\ : std_logic;
signal \N__53502\ : std_logic;
signal \N__53501\ : std_logic;
signal \N__53494\ : std_logic;
signal \N__53493\ : std_logic;
signal \N__53492\ : std_logic;
signal \N__53485\ : std_logic;
signal \N__53484\ : std_logic;
signal \N__53483\ : std_logic;
signal \N__53476\ : std_logic;
signal \N__53475\ : std_logic;
signal \N__53474\ : std_logic;
signal \N__53457\ : std_logic;
signal \N__53454\ : std_logic;
signal \N__53451\ : std_logic;
signal \N__53450\ : std_logic;
signal \N__53449\ : std_logic;
signal \N__53446\ : std_logic;
signal \N__53443\ : std_logic;
signal \N__53440\ : std_logic;
signal \N__53437\ : std_logic;
signal \N__53436\ : std_logic;
signal \N__53433\ : std_logic;
signal \N__53430\ : std_logic;
signal \N__53427\ : std_logic;
signal \N__53424\ : std_logic;
signal \N__53415\ : std_logic;
signal \N__53414\ : std_logic;
signal \N__53411\ : std_logic;
signal \N__53410\ : std_logic;
signal \N__53407\ : std_logic;
signal \N__53406\ : std_logic;
signal \N__53405\ : std_logic;
signal \N__53402\ : std_logic;
signal \N__53399\ : std_logic;
signal \N__53396\ : std_logic;
signal \N__53395\ : std_logic;
signal \N__53390\ : std_logic;
signal \N__53387\ : std_logic;
signal \N__53382\ : std_logic;
signal \N__53379\ : std_logic;
signal \N__53372\ : std_logic;
signal \N__53369\ : std_logic;
signal \N__53364\ : std_logic;
signal \N__53361\ : std_logic;
signal \N__53358\ : std_logic;
signal \N__53357\ : std_logic;
signal \N__53354\ : std_logic;
signal \N__53351\ : std_logic;
signal \N__53346\ : std_logic;
signal \N__53343\ : std_logic;
signal \N__53340\ : std_logic;
signal \N__53337\ : std_logic;
signal \N__53336\ : std_logic;
signal \N__53335\ : std_logic;
signal \N__53332\ : std_logic;
signal \N__53331\ : std_logic;
signal \N__53326\ : std_logic;
signal \N__53323\ : std_logic;
signal \N__53322\ : std_logic;
signal \N__53319\ : std_logic;
signal \N__53316\ : std_logic;
signal \N__53313\ : std_logic;
signal \N__53310\ : std_logic;
signal \N__53305\ : std_logic;
signal \N__53298\ : std_logic;
signal \N__53295\ : std_logic;
signal \N__53292\ : std_logic;
signal \N__53289\ : std_logic;
signal \N__53286\ : std_logic;
signal \N__53283\ : std_logic;
signal \N__53282\ : std_logic;
signal \N__53281\ : std_logic;
signal \N__53280\ : std_logic;
signal \N__53279\ : std_logic;
signal \N__53278\ : std_logic;
signal \N__53277\ : std_logic;
signal \N__53276\ : std_logic;
signal \N__53275\ : std_logic;
signal \N__53274\ : std_logic;
signal \N__53273\ : std_logic;
signal \N__53272\ : std_logic;
signal \N__53271\ : std_logic;
signal \N__53270\ : std_logic;
signal \N__53269\ : std_logic;
signal \N__53268\ : std_logic;
signal \N__53267\ : std_logic;
signal \N__53266\ : std_logic;
signal \N__53265\ : std_logic;
signal \N__53264\ : std_logic;
signal \N__53263\ : std_logic;
signal \N__53262\ : std_logic;
signal \N__53261\ : std_logic;
signal \N__53260\ : std_logic;
signal \N__53259\ : std_logic;
signal \N__53258\ : std_logic;
signal \N__53257\ : std_logic;
signal \N__53256\ : std_logic;
signal \N__53255\ : std_logic;
signal \N__53254\ : std_logic;
signal \N__53253\ : std_logic;
signal \N__53252\ : std_logic;
signal \N__53251\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53249\ : std_logic;
signal \N__53248\ : std_logic;
signal \N__53247\ : std_logic;
signal \N__53246\ : std_logic;
signal \N__53245\ : std_logic;
signal \N__53244\ : std_logic;
signal \N__53243\ : std_logic;
signal \N__53242\ : std_logic;
signal \N__53241\ : std_logic;
signal \N__53154\ : std_logic;
signal \N__53151\ : std_logic;
signal \N__53148\ : std_logic;
signal \N__53147\ : std_logic;
signal \N__53146\ : std_logic;
signal \N__53145\ : std_logic;
signal \N__53144\ : std_logic;
signal \N__53143\ : std_logic;
signal \N__53142\ : std_logic;
signal \N__53141\ : std_logic;
signal \N__53140\ : std_logic;
signal \N__53139\ : std_logic;
signal \N__53138\ : std_logic;
signal \N__53137\ : std_logic;
signal \N__53136\ : std_logic;
signal \N__53135\ : std_logic;
signal \N__53134\ : std_logic;
signal \N__53133\ : std_logic;
signal \N__53132\ : std_logic;
signal \N__53131\ : std_logic;
signal \N__53130\ : std_logic;
signal \N__53129\ : std_logic;
signal \N__53128\ : std_logic;
signal \N__53127\ : std_logic;
signal \N__53126\ : std_logic;
signal \N__53125\ : std_logic;
signal \N__53124\ : std_logic;
signal \N__53123\ : std_logic;
signal \N__53122\ : std_logic;
signal \N__53121\ : std_logic;
signal \N__53120\ : std_logic;
signal \N__53119\ : std_logic;
signal \N__53118\ : std_logic;
signal \N__53117\ : std_logic;
signal \N__53116\ : std_logic;
signal \N__53115\ : std_logic;
signal \N__53114\ : std_logic;
signal \N__53113\ : std_logic;
signal \N__53112\ : std_logic;
signal \N__53111\ : std_logic;
signal \N__53110\ : std_logic;
signal \N__53109\ : std_logic;
signal \N__53108\ : std_logic;
signal \N__53107\ : std_logic;
signal \N__53106\ : std_logic;
signal \N__53105\ : std_logic;
signal \N__53104\ : std_logic;
signal \N__53103\ : std_logic;
signal \N__53102\ : std_logic;
signal \N__53101\ : std_logic;
signal \N__53100\ : std_logic;
signal \N__53099\ : std_logic;
signal \N__53098\ : std_logic;
signal \N__53097\ : std_logic;
signal \N__53096\ : std_logic;
signal \N__53095\ : std_logic;
signal \N__53094\ : std_logic;
signal \N__53093\ : std_logic;
signal \N__53092\ : std_logic;
signal \N__53091\ : std_logic;
signal \N__53090\ : std_logic;
signal \N__53089\ : std_logic;
signal \N__53088\ : std_logic;
signal \N__53087\ : std_logic;
signal \N__53086\ : std_logic;
signal \N__53085\ : std_logic;
signal \N__53084\ : std_logic;
signal \N__53083\ : std_logic;
signal \N__53082\ : std_logic;
signal \N__53081\ : std_logic;
signal \N__53080\ : std_logic;
signal \N__53079\ : std_logic;
signal \N__53078\ : std_logic;
signal \N__53077\ : std_logic;
signal \N__53076\ : std_logic;
signal \N__53075\ : std_logic;
signal \N__53074\ : std_logic;
signal \N__53073\ : std_logic;
signal \N__53072\ : std_logic;
signal \N__53071\ : std_logic;
signal \N__53070\ : std_logic;
signal \N__53069\ : std_logic;
signal \N__53068\ : std_logic;
signal \N__53067\ : std_logic;
signal \N__53066\ : std_logic;
signal \N__53065\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53063\ : std_logic;
signal \N__53062\ : std_logic;
signal \N__53061\ : std_logic;
signal \N__53060\ : std_logic;
signal \N__53059\ : std_logic;
signal \N__53058\ : std_logic;
signal \N__53057\ : std_logic;
signal \N__53056\ : std_logic;
signal \N__53055\ : std_logic;
signal \N__53054\ : std_logic;
signal \N__53053\ : std_logic;
signal \N__53052\ : std_logic;
signal \N__53051\ : std_logic;
signal \N__53050\ : std_logic;
signal \N__53049\ : std_logic;
signal \N__53048\ : std_logic;
signal \N__53047\ : std_logic;
signal \N__53046\ : std_logic;
signal \N__53045\ : std_logic;
signal \N__53044\ : std_logic;
signal \N__53043\ : std_logic;
signal \N__53042\ : std_logic;
signal \N__53041\ : std_logic;
signal \N__53040\ : std_logic;
signal \N__53039\ : std_logic;
signal \N__53038\ : std_logic;
signal \N__53037\ : std_logic;
signal \N__53036\ : std_logic;
signal \N__53035\ : std_logic;
signal \N__53034\ : std_logic;
signal \N__53033\ : std_logic;
signal \N__53032\ : std_logic;
signal \N__53031\ : std_logic;
signal \N__53030\ : std_logic;
signal \N__53029\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53027\ : std_logic;
signal \N__53026\ : std_logic;
signal \N__53025\ : std_logic;
signal \N__53024\ : std_logic;
signal \N__53023\ : std_logic;
signal \N__53022\ : std_logic;
signal \N__53021\ : std_logic;
signal \N__53020\ : std_logic;
signal \N__53019\ : std_logic;
signal \N__53018\ : std_logic;
signal \N__53017\ : std_logic;
signal \N__53016\ : std_logic;
signal \N__53015\ : std_logic;
signal \N__53014\ : std_logic;
signal \N__53013\ : std_logic;
signal \N__53012\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53010\ : std_logic;
signal \N__53009\ : std_logic;
signal \N__53008\ : std_logic;
signal \N__53007\ : std_logic;
signal \N__53006\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__53004\ : std_logic;
signal \N__53003\ : std_logic;
signal \N__53002\ : std_logic;
signal \N__53001\ : std_logic;
signal \N__53000\ : std_logic;
signal \N__52999\ : std_logic;
signal \N__52998\ : std_logic;
signal \N__52997\ : std_logic;
signal \N__52996\ : std_logic;
signal \N__52995\ : std_logic;
signal \N__52994\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52992\ : std_logic;
signal \N__52991\ : std_logic;
signal \N__52990\ : std_logic;
signal \N__52989\ : std_logic;
signal \N__52988\ : std_logic;
signal \N__52987\ : std_logic;
signal \N__52986\ : std_logic;
signal \N__52985\ : std_logic;
signal \N__52984\ : std_logic;
signal \N__52983\ : std_logic;
signal \N__52982\ : std_logic;
signal \N__52981\ : std_logic;
signal \N__52980\ : std_logic;
signal \N__52979\ : std_logic;
signal \N__52978\ : std_logic;
signal \N__52977\ : std_logic;
signal \N__52976\ : std_logic;
signal \N__52975\ : std_logic;
signal \N__52974\ : std_logic;
signal \N__52973\ : std_logic;
signal \N__52972\ : std_logic;
signal \N__52971\ : std_logic;
signal \N__52970\ : std_logic;
signal \N__52969\ : std_logic;
signal \N__52968\ : std_logic;
signal \N__52967\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52599\ : std_logic;
signal \N__52596\ : std_logic;
signal \N__52593\ : std_logic;
signal \N__52592\ : std_logic;
signal \N__52589\ : std_logic;
signal \N__52586\ : std_logic;
signal \N__52583\ : std_logic;
signal \N__52580\ : std_logic;
signal \N__52577\ : std_logic;
signal \N__52574\ : std_logic;
signal \N__52569\ : std_logic;
signal \N__52566\ : std_logic;
signal \N__52563\ : std_logic;
signal \N__52560\ : std_logic;
signal \N__52557\ : std_logic;
signal \N__52554\ : std_logic;
signal \N__52551\ : std_logic;
signal \N__52548\ : std_logic;
signal \N__52547\ : std_logic;
signal \N__52542\ : std_logic;
signal \N__52541\ : std_logic;
signal \N__52540\ : std_logic;
signal \N__52537\ : std_logic;
signal \N__52534\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52524\ : std_logic;
signal \N__52521\ : std_logic;
signal \N__52520\ : std_logic;
signal \N__52519\ : std_logic;
signal \N__52516\ : std_logic;
signal \N__52513\ : std_logic;
signal \N__52512\ : std_logic;
signal \N__52511\ : std_logic;
signal \N__52508\ : std_logic;
signal \N__52503\ : std_logic;
signal \N__52500\ : std_logic;
signal \N__52497\ : std_logic;
signal \N__52488\ : std_logic;
signal \N__52487\ : std_logic;
signal \N__52484\ : std_logic;
signal \N__52481\ : std_logic;
signal \N__52476\ : std_logic;
signal \N__52475\ : std_logic;
signal \N__52472\ : std_logic;
signal \N__52469\ : std_logic;
signal \N__52464\ : std_logic;
signal \N__52463\ : std_logic;
signal \N__52460\ : std_logic;
signal \N__52457\ : std_logic;
signal \N__52454\ : std_logic;
signal \N__52449\ : std_logic;
signal \N__52446\ : std_logic;
signal \N__52445\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52441\ : std_logic;
signal \N__52438\ : std_logic;
signal \N__52435\ : std_logic;
signal \N__52430\ : std_logic;
signal \N__52425\ : std_logic;
signal \N__52422\ : std_logic;
signal \N__52421\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52419\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52415\ : std_logic;
signal \N__52414\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52404\ : std_logic;
signal \N__52401\ : std_logic;
signal \N__52398\ : std_logic;
signal \N__52395\ : std_logic;
signal \N__52390\ : std_logic;
signal \N__52387\ : std_logic;
signal \N__52384\ : std_logic;
signal \N__52381\ : std_logic;
signal \N__52378\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52372\ : std_logic;
signal \N__52369\ : std_logic;
signal \N__52362\ : std_logic;
signal \N__52359\ : std_logic;
signal \N__52356\ : std_logic;
signal \N__52353\ : std_logic;
signal \N__52350\ : std_logic;
signal \N__52347\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52343\ : std_logic;
signal \N__52340\ : std_logic;
signal \N__52337\ : std_logic;
signal \N__52334\ : std_logic;
signal \N__52331\ : std_logic;
signal \N__52328\ : std_logic;
signal \N__52325\ : std_logic;
signal \N__52320\ : std_logic;
signal \N__52317\ : std_logic;
signal \N__52314\ : std_logic;
signal \N__52311\ : std_logic;
signal \N__52308\ : std_logic;
signal \N__52305\ : std_logic;
signal \N__52304\ : std_logic;
signal \N__52301\ : std_logic;
signal \N__52298\ : std_logic;
signal \N__52297\ : std_logic;
signal \N__52296\ : std_logic;
signal \N__52291\ : std_logic;
signal \N__52288\ : std_logic;
signal \N__52285\ : std_logic;
signal \N__52278\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52272\ : std_logic;
signal \N__52269\ : std_logic;
signal \N__52266\ : std_logic;
signal \N__52263\ : std_logic;
signal \N__52260\ : std_logic;
signal \N__52257\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52253\ : std_logic;
signal \N__52250\ : std_logic;
signal \N__52247\ : std_logic;
signal \N__52244\ : std_logic;
signal \N__52241\ : std_logic;
signal \N__52236\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52232\ : std_logic;
signal \N__52229\ : std_logic;
signal \N__52226\ : std_logic;
signal \N__52225\ : std_logic;
signal \N__52222\ : std_logic;
signal \N__52219\ : std_logic;
signal \N__52216\ : std_logic;
signal \N__52213\ : std_logic;
signal \N__52206\ : std_logic;
signal \N__52203\ : std_logic;
signal \N__52200\ : std_logic;
signal \N__52199\ : std_logic;
signal \N__52194\ : std_logic;
signal \N__52193\ : std_logic;
signal \N__52190\ : std_logic;
signal \N__52187\ : std_logic;
signal \N__52184\ : std_logic;
signal \N__52179\ : std_logic;
signal \N__52176\ : std_logic;
signal \N__52173\ : std_logic;
signal \N__52170\ : std_logic;
signal \N__52167\ : std_logic;
signal \N__52164\ : std_logic;
signal \N__52161\ : std_logic;
signal \N__52160\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52158\ : std_logic;
signal \N__52157\ : std_logic;
signal \N__52156\ : std_logic;
signal \N__52155\ : std_logic;
signal \N__52154\ : std_logic;
signal \N__52153\ : std_logic;
signal \N__52152\ : std_logic;
signal \N__52151\ : std_logic;
signal \N__52150\ : std_logic;
signal \N__52149\ : std_logic;
signal \N__52148\ : std_logic;
signal \N__52147\ : std_logic;
signal \N__52146\ : std_logic;
signal \N__52145\ : std_logic;
signal \N__52144\ : std_logic;
signal \N__52143\ : std_logic;
signal \N__52142\ : std_logic;
signal \N__52141\ : std_logic;
signal \N__52140\ : std_logic;
signal \N__52139\ : std_logic;
signal \N__52138\ : std_logic;
signal \N__52137\ : std_logic;
signal \N__52132\ : std_logic;
signal \N__52123\ : std_logic;
signal \N__52122\ : std_logic;
signal \N__52121\ : std_logic;
signal \N__52120\ : std_logic;
signal \N__52119\ : std_logic;
signal \N__52118\ : std_logic;
signal \N__52117\ : std_logic;
signal \N__52116\ : std_logic;
signal \N__52115\ : std_logic;
signal \N__52114\ : std_logic;
signal \N__52113\ : std_logic;
signal \N__52112\ : std_logic;
signal \N__52111\ : std_logic;
signal \N__52110\ : std_logic;
signal \N__52109\ : std_logic;
signal \N__52108\ : std_logic;
signal \N__52107\ : std_logic;
signal \N__52106\ : std_logic;
signal \N__52105\ : std_logic;
signal \N__52104\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52096\ : std_logic;
signal \N__52095\ : std_logic;
signal \N__52094\ : std_logic;
signal \N__52093\ : std_logic;
signal \N__52092\ : std_logic;
signal \N__52091\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52083\ : std_logic;
signal \N__52082\ : std_logic;
signal \N__52081\ : std_logic;
signal \N__52080\ : std_logic;
signal \N__52079\ : std_logic;
signal \N__52078\ : std_logic;
signal \N__52077\ : std_logic;
signal \N__52076\ : std_logic;
signal \N__52075\ : std_logic;
signal \N__52074\ : std_logic;
signal \N__52073\ : std_logic;
signal \N__52068\ : std_logic;
signal \N__52067\ : std_logic;
signal \N__52066\ : std_logic;
signal \N__52065\ : std_logic;
signal \N__52064\ : std_logic;
signal \N__52059\ : std_logic;
signal \N__52054\ : std_logic;
signal \N__52047\ : std_logic;
signal \N__52042\ : std_logic;
signal \N__52041\ : std_logic;
signal \N__52036\ : std_logic;
signal \N__52031\ : std_logic;
signal \N__52028\ : std_logic;
signal \N__52023\ : std_logic;
signal \N__52020\ : std_logic;
signal \N__52019\ : std_logic;
signal \N__52018\ : std_logic;
signal \N__52017\ : std_logic;
signal \N__52016\ : std_logic;
signal \N__52015\ : std_logic;
signal \N__52014\ : std_logic;
signal \N__52013\ : std_logic;
signal \N__52012\ : std_logic;
signal \N__52009\ : std_logic;
signal \N__52008\ : std_logic;
signal \N__52007\ : std_logic;
signal \N__52006\ : std_logic;
signal \N__52005\ : std_logic;
signal \N__52004\ : std_logic;
signal \N__52003\ : std_logic;
signal \N__52002\ : std_logic;
signal \N__52001\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51999\ : std_logic;
signal \N__51998\ : std_logic;
signal \N__51997\ : std_logic;
signal \N__51996\ : std_logic;
signal \N__51995\ : std_logic;
signal \N__51994\ : std_logic;
signal \N__51993\ : std_logic;
signal \N__51986\ : std_logic;
signal \N__51985\ : std_logic;
signal \N__51984\ : std_logic;
signal \N__51983\ : std_logic;
signal \N__51980\ : std_logic;
signal \N__51975\ : std_logic;
signal \N__51974\ : std_logic;
signal \N__51973\ : std_logic;
signal \N__51972\ : std_logic;
signal \N__51971\ : std_logic;
signal \N__51970\ : std_logic;
signal \N__51963\ : std_logic;
signal \N__51958\ : std_logic;
signal \N__51951\ : std_logic;
signal \N__51948\ : std_logic;
signal \N__51945\ : std_logic;
signal \N__51934\ : std_logic;
signal \N__51931\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51917\ : std_logic;
signal \N__51914\ : std_logic;
signal \N__51911\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51909\ : std_logic;
signal \N__51908\ : std_logic;
signal \N__51907\ : std_logic;
signal \N__51906\ : std_logic;
signal \N__51905\ : std_logic;
signal \N__51904\ : std_logic;
signal \N__51903\ : std_logic;
signal \N__51902\ : std_logic;
signal \N__51897\ : std_logic;
signal \N__51896\ : std_logic;
signal \N__51895\ : std_logic;
signal \N__51894\ : std_logic;
signal \N__51893\ : std_logic;
signal \N__51892\ : std_logic;
signal \N__51891\ : std_logic;
signal \N__51890\ : std_logic;
signal \N__51889\ : std_logic;
signal \N__51888\ : std_logic;
signal \N__51887\ : std_logic;
signal \N__51886\ : std_logic;
signal \N__51885\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51881\ : std_logic;
signal \N__51880\ : std_logic;
signal \N__51879\ : std_logic;
signal \N__51878\ : std_logic;
signal \N__51875\ : std_logic;
signal \N__51868\ : std_logic;
signal \N__51867\ : std_logic;
signal \N__51866\ : std_logic;
signal \N__51865\ : std_logic;
signal \N__51864\ : std_logic;
signal \N__51861\ : std_logic;
signal \N__51858\ : std_logic;
signal \N__51851\ : std_logic;
signal \N__51848\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51836\ : std_logic;
signal \N__51831\ : std_logic;
signal \N__51826\ : std_logic;
signal \N__51819\ : std_logic;
signal \N__51818\ : std_logic;
signal \N__51817\ : std_logic;
signal \N__51816\ : std_logic;
signal \N__51815\ : std_logic;
signal \N__51814\ : std_logic;
signal \N__51813\ : std_logic;
signal \N__51812\ : std_logic;
signal \N__51811\ : std_logic;
signal \N__51810\ : std_logic;
signal \N__51809\ : std_logic;
signal \N__51808\ : std_logic;
signal \N__51805\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51803\ : std_logic;
signal \N__51802\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51785\ : std_logic;
signal \N__51778\ : std_logic;
signal \N__51773\ : std_logic;
signal \N__51772\ : std_logic;
signal \N__51771\ : std_logic;
signal \N__51770\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51758\ : std_logic;
signal \N__51755\ : std_logic;
signal \N__51752\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51742\ : std_logic;
signal \N__51737\ : std_logic;
signal \N__51730\ : std_logic;
signal \N__51727\ : std_logic;
signal \N__51722\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51704\ : std_logic;
signal \N__51695\ : std_logic;
signal \N__51684\ : std_logic;
signal \N__51681\ : std_logic;
signal \N__51678\ : std_logic;
signal \N__51671\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51663\ : std_logic;
signal \N__51656\ : std_logic;
signal \N__51651\ : std_logic;
signal \N__51648\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51638\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51624\ : std_logic;
signal \N__51617\ : std_logic;
signal \N__51610\ : std_logic;
signal \N__51603\ : std_logic;
signal \N__51602\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51600\ : std_logic;
signal \N__51599\ : std_logic;
signal \N__51598\ : std_logic;
signal \N__51597\ : std_logic;
signal \N__51596\ : std_logic;
signal \N__51595\ : std_logic;
signal \N__51594\ : std_logic;
signal \N__51589\ : std_logic;
signal \N__51582\ : std_logic;
signal \N__51577\ : std_logic;
signal \N__51570\ : std_logic;
signal \N__51565\ : std_logic;
signal \N__51556\ : std_logic;
signal \N__51555\ : std_logic;
signal \N__51554\ : std_logic;
signal \N__51553\ : std_logic;
signal \N__51552\ : std_logic;
signal \N__51551\ : std_logic;
signal \N__51542\ : std_logic;
signal \N__51541\ : std_logic;
signal \N__51540\ : std_logic;
signal \N__51539\ : std_logic;
signal \N__51538\ : std_logic;
signal \N__51537\ : std_logic;
signal \N__51530\ : std_logic;
signal \N__51521\ : std_logic;
signal \N__51514\ : std_logic;
signal \N__51503\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51501\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51495\ : std_logic;
signal \N__51494\ : std_logic;
signal \N__51493\ : std_logic;
signal \N__51490\ : std_logic;
signal \N__51481\ : std_logic;
signal \N__51480\ : std_logic;
signal \N__51479\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51477\ : std_logic;
signal \N__51472\ : std_logic;
signal \N__51461\ : std_logic;
signal \N__51454\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51434\ : std_logic;
signal \N__51421\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51395\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51370\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51355\ : std_logic;
signal \N__51348\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51334\ : std_logic;
signal \N__51329\ : std_logic;
signal \N__51306\ : std_logic;
signal \N__51303\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51297\ : std_logic;
signal \N__51294\ : std_logic;
signal \N__51291\ : std_logic;
signal \N__51288\ : std_logic;
signal \N__51285\ : std_logic;
signal \N__51282\ : std_logic;
signal \N__51279\ : std_logic;
signal \N__51276\ : std_logic;
signal \N__51273\ : std_logic;
signal \N__51272\ : std_logic;
signal \N__51271\ : std_logic;
signal \N__51270\ : std_logic;
signal \N__51269\ : std_logic;
signal \N__51268\ : std_logic;
signal \N__51267\ : std_logic;
signal \N__51266\ : std_logic;
signal \N__51263\ : std_logic;
signal \N__51262\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51260\ : std_logic;
signal \N__51259\ : std_logic;
signal \N__51258\ : std_logic;
signal \N__51257\ : std_logic;
signal \N__51254\ : std_logic;
signal \N__51253\ : std_logic;
signal \N__51252\ : std_logic;
signal \N__51249\ : std_logic;
signal \N__51248\ : std_logic;
signal \N__51247\ : std_logic;
signal \N__51246\ : std_logic;
signal \N__51243\ : std_logic;
signal \N__51242\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51240\ : std_logic;
signal \N__51239\ : std_logic;
signal \N__51236\ : std_logic;
signal \N__51233\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51229\ : std_logic;
signal \N__51226\ : std_logic;
signal \N__51223\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51217\ : std_logic;
signal \N__51216\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51210\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51203\ : std_logic;
signal \N__51200\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51188\ : std_logic;
signal \N__51185\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51181\ : std_logic;
signal \N__51178\ : std_logic;
signal \N__51175\ : std_logic;
signal \N__51172\ : std_logic;
signal \N__51169\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51165\ : std_logic;
signal \N__51164\ : std_logic;
signal \N__51159\ : std_logic;
signal \N__51158\ : std_logic;
signal \N__51157\ : std_logic;
signal \N__51156\ : std_logic;
signal \N__51155\ : std_logic;
signal \N__51152\ : std_logic;
signal \N__51147\ : std_logic;
signal \N__51140\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51138\ : std_logic;
signal \N__51135\ : std_logic;
signal \N__51134\ : std_logic;
signal \N__51133\ : std_logic;
signal \N__51132\ : std_logic;
signal \N__51127\ : std_logic;
signal \N__51122\ : std_logic;
signal \N__51119\ : std_logic;
signal \N__51112\ : std_logic;
signal \N__51105\ : std_logic;
signal \N__51102\ : std_logic;
signal \N__51101\ : std_logic;
signal \N__51100\ : std_logic;
signal \N__51099\ : std_logic;
signal \N__51096\ : std_logic;
signal \N__51087\ : std_logic;
signal \N__51084\ : std_logic;
signal \N__51083\ : std_logic;
signal \N__51082\ : std_logic;
signal \N__51081\ : std_logic;
signal \N__51080\ : std_logic;
signal \N__51079\ : std_logic;
signal \N__51078\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51072\ : std_logic;
signal \N__51069\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51063\ : std_logic;
signal \N__51060\ : std_logic;
signal \N__51057\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51051\ : std_logic;
signal \N__51048\ : std_logic;
signal \N__51045\ : std_logic;
signal \N__51042\ : std_logic;
signal \N__51041\ : std_logic;
signal \N__51040\ : std_logic;
signal \N__51037\ : std_logic;
signal \N__51034\ : std_logic;
signal \N__51031\ : std_logic;
signal \N__51028\ : std_logic;
signal \N__51027\ : std_logic;
signal \N__51026\ : std_logic;
signal \N__51025\ : std_logic;
signal \N__51024\ : std_logic;
signal \N__51017\ : std_logic;
signal \N__51010\ : std_logic;
signal \N__51007\ : std_logic;
signal \N__51004\ : std_logic;
signal \N__51001\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50991\ : std_logic;
signal \N__50988\ : std_logic;
signal \N__50987\ : std_logic;
signal \N__50986\ : std_logic;
signal \N__50983\ : std_logic;
signal \N__50982\ : std_logic;
signal \N__50981\ : std_logic;
signal \N__50978\ : std_logic;
signal \N__50975\ : std_logic;
signal \N__50972\ : std_logic;
signal \N__50967\ : std_logic;
signal \N__50956\ : std_logic;
signal \N__50953\ : std_logic;
signal \N__50944\ : std_logic;
signal \N__50941\ : std_logic;
signal \N__50938\ : std_logic;
signal \N__50929\ : std_logic;
signal \N__50926\ : std_logic;
signal \N__50923\ : std_logic;
signal \N__50920\ : std_logic;
signal \N__50917\ : std_logic;
signal \N__50914\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50898\ : std_logic;
signal \N__50895\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50889\ : std_logic;
signal \N__50886\ : std_logic;
signal \N__50883\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50881\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50873\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50867\ : std_logic;
signal \N__50860\ : std_logic;
signal \N__50857\ : std_logic;
signal \N__50846\ : std_logic;
signal \N__50835\ : std_logic;
signal \N__50828\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50819\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50801\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50789\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50771\ : std_logic;
signal \N__50770\ : std_logic;
signal \N__50769\ : std_logic;
signal \N__50766\ : std_logic;
signal \N__50763\ : std_logic;
signal \N__50762\ : std_logic;
signal \N__50761\ : std_logic;
signal \N__50758\ : std_logic;
signal \N__50755\ : std_logic;
signal \N__50754\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50747\ : std_logic;
signal \N__50744\ : std_logic;
signal \N__50741\ : std_logic;
signal \N__50740\ : std_logic;
signal \N__50735\ : std_logic;
signal \N__50734\ : std_logic;
signal \N__50733\ : std_logic;
signal \N__50732\ : std_logic;
signal \N__50729\ : std_logic;
signal \N__50726\ : std_logic;
signal \N__50725\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50723\ : std_logic;
signal \N__50714\ : std_logic;
signal \N__50711\ : std_logic;
signal \N__50710\ : std_logic;
signal \N__50709\ : std_logic;
signal \N__50708\ : std_logic;
signal \N__50707\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50701\ : std_logic;
signal \N__50698\ : std_logic;
signal \N__50695\ : std_logic;
signal \N__50694\ : std_logic;
signal \N__50693\ : std_logic;
signal \N__50692\ : std_logic;
signal \N__50691\ : std_logic;
signal \N__50688\ : std_logic;
signal \N__50687\ : std_logic;
signal \N__50686\ : std_logic;
signal \N__50685\ : std_logic;
signal \N__50682\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50678\ : std_logic;
signal \N__50677\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50675\ : std_logic;
signal \N__50674\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50672\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50665\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50659\ : std_logic;
signal \N__50656\ : std_logic;
signal \N__50653\ : std_logic;
signal \N__50650\ : std_logic;
signal \N__50647\ : std_logic;
signal \N__50638\ : std_logic;
signal \N__50635\ : std_logic;
signal \N__50632\ : std_logic;
signal \N__50629\ : std_logic;
signal \N__50626\ : std_logic;
signal \N__50625\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50619\ : std_logic;
signal \N__50616\ : std_logic;
signal \N__50613\ : std_logic;
signal \N__50608\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50602\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50600\ : std_logic;
signal \N__50599\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50593\ : std_logic;
signal \N__50592\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50585\ : std_logic;
signal \N__50584\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50582\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50577\ : std_logic;
signal \N__50576\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50574\ : std_logic;
signal \N__50573\ : std_logic;
signal \N__50572\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50564\ : std_logic;
signal \N__50561\ : std_logic;
signal \N__50560\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50542\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50534\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50504\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50497\ : std_logic;
signal \N__50494\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50488\ : std_logic;
signal \N__50485\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50476\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50467\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50461\ : std_logic;
signal \N__50458\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50451\ : std_logic;
signal \N__50448\ : std_logic;
signal \N__50445\ : std_logic;
signal \N__50442\ : std_logic;
signal \N__50439\ : std_logic;
signal \N__50432\ : std_logic;
signal \N__50423\ : std_logic;
signal \N__50422\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50369\ : std_logic;
signal \N__50360\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50352\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50327\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50242\ : std_logic;
signal \N__50241\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50231\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50221\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50210\ : std_logic;
signal \N__50207\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50197\ : std_logic;
signal \N__50194\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50180\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50174\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50161\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50144\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50124\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50112\ : std_logic;
signal \N__50109\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50094\ : std_logic;
signal \N__50093\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50090\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50084\ : std_logic;
signal \N__50081\ : std_logic;
signal \N__50080\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50078\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50074\ : std_logic;
signal \N__50063\ : std_logic;
signal \N__50060\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50044\ : std_logic;
signal \N__50039\ : std_logic;
signal \N__50036\ : std_logic;
signal \N__50033\ : std_logic;
signal \N__50030\ : std_logic;
signal \N__50027\ : std_logic;
signal \N__50026\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50024\ : std_logic;
signal \N__50023\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49984\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49885\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49870\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49836\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49826\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49823\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49799\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49787\ : std_logic;
signal \N__49786\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49784\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49769\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49766\ : std_logic;
signal \N__49765\ : std_logic;
signal \N__49762\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49737\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49720\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49702\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49689\ : std_logic;
signal \N__49686\ : std_logic;
signal \N__49677\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49668\ : std_logic;
signal \N__49665\ : std_logic;
signal \N__49662\ : std_logic;
signal \N__49661\ : std_logic;
signal \N__49652\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49646\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49592\ : std_logic;
signal \N__49591\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49587\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49579\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49575\ : std_logic;
signal \N__49574\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49572\ : std_logic;
signal \N__49571\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49415\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49400\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49377\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49367\ : std_logic;
signal \N__49364\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49358\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49355\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49346\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49328\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49319\ : std_logic;
signal \N__49316\ : std_logic;
signal \N__49313\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49307\ : std_logic;
signal \N__49306\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49291\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49285\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49276\ : std_logic;
signal \N__49273\ : std_logic;
signal \N__49270\ : std_logic;
signal \N__49267\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49261\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49254\ : std_logic;
signal \N__49251\ : std_logic;
signal \N__49248\ : std_logic;
signal \N__49241\ : std_logic;
signal \N__49238\ : std_logic;
signal \N__49235\ : std_logic;
signal \N__49232\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49226\ : std_logic;
signal \N__49223\ : std_logic;
signal \N__49222\ : std_logic;
signal \N__49219\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49207\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49199\ : std_logic;
signal \N__49190\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49181\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49177\ : std_logic;
signal \N__49172\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49166\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49160\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49152\ : std_logic;
signal \N__49149\ : std_logic;
signal \N__49146\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49106\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49092\ : std_logic;
signal \N__49091\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49085\ : std_logic;
signal \N__49082\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49076\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49068\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49057\ : std_logic;
signal \N__49052\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49028\ : std_logic;
signal \N__49025\ : std_logic;
signal \N__49022\ : std_logic;
signal \N__49019\ : std_logic;
signal \N__49016\ : std_logic;
signal \N__49009\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48993\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48989\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48982\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48930\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48897\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48882\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48843\ : std_logic;
signal \N__48842\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48835\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48832\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48818\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48813\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48744\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48669\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48664\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48634\ : std_logic;
signal \N__48633\ : std_logic;
signal \N__48630\ : std_logic;
signal \N__48627\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48621\ : std_logic;
signal \N__48618\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48600\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48552\ : std_logic;
signal \N__48549\ : std_logic;
signal \N__48546\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48540\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48433\ : std_logic;
signal \N__48428\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48312\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48306\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48294\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48274\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48255\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48230\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48124\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48062\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48031\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47975\ : std_logic;
signal \N__47972\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47960\ : std_logic;
signal \N__47949\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47926\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47920\ : std_logic;
signal \N__47917\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47899\ : std_logic;
signal \N__47896\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47884\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47856\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47767\ : std_logic;
signal \N__47766\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47748\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47720\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47717\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47715\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47334\ : std_logic;
signal \N__47331\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47300\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47235\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47187\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47144\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47130\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47126\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46998\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46868\ : std_logic;
signal \N__46865\ : std_logic;
signal \N__46862\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46759\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46738\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46702\ : std_logic;
signal \N__46699\ : std_logic;
signal \N__46690\ : std_logic;
signal \N__46687\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46574\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46565\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46532\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46486\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46451\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46414\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46398\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46365\ : std_logic;
signal \N__46362\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46283\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46247\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46190\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46141\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46123\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46088\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46069\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45938\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45910\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45892\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45889\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45883\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45880\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45828\ : std_logic;
signal \N__45825\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45817\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45808\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45780\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45706\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45690\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45521\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45518\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45496\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45440\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45421\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45372\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45300\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45291\ : std_logic;
signal \N__45288\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45258\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45189\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45168\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45009\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44993\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44981\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44912\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44855\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44825\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44794\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44759\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44750\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44637\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44594\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44511\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44319\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44307\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44126\ : std_logic;
signal \N__44123\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44110\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44067\ : std_logic;
signal \N__44064\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44030\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44023\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44008\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43989\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43941\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43935\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43875\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43868\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43846\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43843\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43832\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43792\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43765\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43759\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43731\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43689\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43675\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43662\ : std_logic;
signal \N__43659\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43564\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43551\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43503\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43479\ : std_logic;
signal \N__43476\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43396\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43216\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43208\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43191\ : std_logic;
signal \N__43190\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43178\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43130\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43026\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42971\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42919\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42732\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42611\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42529\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42526\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42476\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42338\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42292\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42240\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42234\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42000\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41845\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41839\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41710\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41556\ : std_logic;
signal \N__41553\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41421\ : std_logic;
signal \N__41418\ : std_logic;
signal \N__41415\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41205\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41175\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41118\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40980\ : std_logic;
signal \N__40977\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40695\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40677\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40630\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40513\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40402\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40399\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40396\ : std_logic;
signal \N__40395\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40360\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40348\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40334\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40301\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40283\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40062\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39669\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39267\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39000\ : std_logic;
signal \N__38997\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38370\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38000\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37970\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37937\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37572\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37182\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36347\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36116\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34997\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34606\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33305\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33278\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33256\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33221\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33191\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32792\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32614\ : std_logic;
signal \N__32611\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32423\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32380\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32279\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31993\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31952\ : std_logic;
signal \N__31949\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31616\ : std_logic;
signal \N__31613\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30919\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30903\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30652\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30248\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28670\ : std_logic;
signal \N__28667\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24823\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22164\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal clk_c : std_logic;
signal \pll128M2_inst.pll_clk64_0\ : std_logic;
signal \pll128M2_inst.pll_clk128\ : std_logic;
signal \VCCG0\ : std_logic;
signal button_mode_c : std_logic;
signal \button_mode_ibuf_RNIN5KZ0Z7\ : std_logic;
signal \DAC_cs_c\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i_cascade_\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \sRAM_pointer_read_cry_0\ : std_logic;
signal \sRAM_pointer_read_cry_1\ : std_logic;
signal \sRAM_pointer_read_cry_2\ : std_logic;
signal \sRAM_pointer_read_cry_3\ : std_logic;
signal \sRAM_pointer_read_cry_4\ : std_logic;
signal \sRAM_pointer_read_cry_5\ : std_logic;
signal \sRAM_pointer_read_cry_6\ : std_logic;
signal \sRAM_pointer_read_cry_7\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \sRAM_pointer_read_cry_8\ : std_logic;
signal \sRAM_pointer_read_cry_9\ : std_logic;
signal \sRAM_pointer_read_cry_10\ : std_logic;
signal \sRAM_pointer_read_cry_11\ : std_logic;
signal \sRAM_pointer_read_cry_12\ : std_logic;
signal \sRAM_pointer_read_cry_13\ : std_logic;
signal \sRAM_pointer_read_cry_14\ : std_logic;
signal \sRAM_pointer_read_cry_15\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \sRAM_pointer_read_cry_16\ : std_logic;
signal \sRAM_pointer_read_cry_17\ : std_logic;
signal \N_28_g\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_s_0\ : std_logic;
signal \bfn_3_3_0_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_s_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2\ : std_logic;
signal \bfn_3_4_0_\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO\ : std_logic;
signal \bfn_3_5_0_\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0\ : std_logic;
signal \DAC_mosi_c\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4\ : std_logic;
signal \DAC_sclk_c\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6\ : std_logic;
signal \spi_master_inst.o_sclk_RNIH6AC\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO\ : std_logic;
signal \bfn_5_5_0_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_i_cry_6\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_1666_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_48_cascade_\ : std_logic;
signal \spi_master_inst.ss_start_i\ : std_logic;
signal \sEEPonPoff_i_0\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \sEEPonPoff_i_1\ : std_logic;
signal un4_spoff_cry_0 : std_logic;
signal \sEEPonPoff_i_2\ : std_logic;
signal un4_spoff_cry_1 : std_logic;
signal \sEEPonPoff_i_3\ : std_logic;
signal un4_spoff_cry_2 : std_logic;
signal \sEEPonPoff_i_4\ : std_logic;
signal un4_spoff_cry_3 : std_logic;
signal \sEEPonPoff_i_5\ : std_logic;
signal un4_spoff_cry_4 : std_logic;
signal \sEEPonPoff_i_6\ : std_logic;
signal un4_spoff_cry_5 : std_logic;
signal \sEEPonPoff_i_7\ : std_logic;
signal un4_spoff_cry_6 : std_logic;
signal un4_spoff_cry_7 : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal un4_spoff_cry_8 : std_logic;
signal un4_spoff_cry_9 : std_logic;
signal un4_spoff_cry_10 : std_logic;
signal un4_spoff_cry_11 : std_logic;
signal un4_spoff_cry_12 : std_logic;
signal un4_spoff_cry_13 : std_logic;
signal un4_spoff_cry_14 : std_logic;
signal un4_spoff_cry_15 : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal un4_spoff_cry_16 : std_logic;
signal un4_spoff_cry_17 : std_logic;
signal un4_spoff_cry_18 : std_logic;
signal un4_spoff_cry_19 : std_logic;
signal un4_spoff_cry_20 : std_logic;
signal un4_spoff_cry_21 : std_logic;
signal un4_spoff_cry_22 : std_logic;
signal un4_spoff_cry_23 : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1423\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1416\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1415\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14_cascade_\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1419\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1422\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_1520\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_start_i_i\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15_cascade_\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.N_1412\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_1666\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_1515_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_36_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_48\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_5_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_count_start_iZ0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1\ : std_logic;
signal \sEEPonPoffZ0Z_0\ : std_logic;
signal \sEEPonPoffZ0Z_1\ : std_logic;
signal \sEEPonPoffZ0Z_2\ : std_logic;
signal \sEEPonPoffZ0Z_3\ : std_logic;
signal \sEEPonPoffZ0Z_4\ : std_logic;
signal \sEEPonPoffZ0Z_5\ : std_logic;
signal \sEEPonPoffZ0Z_6\ : std_logic;
signal \sEEPonPoffZ0Z_7\ : std_logic;
signal \sEEPonZ0Z_0\ : std_logic;
signal \sEEPon_i_0\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \sEEPonZ0Z_1\ : std_logic;
signal \sEEPon_i_1\ : std_logic;
signal un7_spon_cry_0 : std_logic;
signal \sEEPonZ0Z_2\ : std_logic;
signal \sEEPon_i_2\ : std_logic;
signal un7_spon_cry_1 : std_logic;
signal \sEEPonZ0Z_3\ : std_logic;
signal \sEEPon_i_3\ : std_logic;
signal un7_spon_cry_2 : std_logic;
signal \sEEPonZ0Z_4\ : std_logic;
signal \sEEPon_i_4\ : std_logic;
signal un7_spon_cry_3 : std_logic;
signal \sEEPonZ0Z_5\ : std_logic;
signal \sEEPon_i_5\ : std_logic;
signal un7_spon_cry_4 : std_logic;
signal \sEEPonZ0Z_6\ : std_logic;
signal \sEEPon_i_6\ : std_logic;
signal un7_spon_cry_5 : std_logic;
signal \sEEPonZ0Z_7\ : std_logic;
signal \sEEPon_i_7\ : std_logic;
signal un7_spon_cry_6 : std_logic;
signal un7_spon_cry_7 : std_logic;
signal \bfn_6_12_0_\ : std_logic;
signal un7_spon_cry_8 : std_logic;
signal un7_spon_cry_9 : std_logic;
signal un7_spon_cry_10 : std_logic;
signal un7_spon_cry_11 : std_logic;
signal un7_spon_cry_12 : std_logic;
signal un7_spon_cry_13 : std_logic;
signal un7_spon_cry_14 : std_logic;
signal un7_spon_cry_15 : std_logic;
signal \bfn_6_13_0_\ : std_logic;
signal un7_spon_cry_16 : std_logic;
signal un7_spon_cry_17 : std_logic;
signal un7_spon_cry_18 : std_logic;
signal un7_spon_cry_19 : std_logic;
signal un7_spon_cry_20 : std_logic;
signal un7_spon_cry_21 : std_logic;
signal un7_spon_cry_22 : std_logic;
signal un7_spon_cry_23 : std_logic;
signal \bfn_6_14_0_\ : std_logic;
signal \pon_obuf_RNOZ0\ : std_logic;
signal g1_0_5 : std_logic;
signal g1 : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1\ : std_logic;
signal \sEESingleContZ0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_1515\ : std_logic;
signal \sEESingleCont_1_sqmuxa\ : std_logic;
signal un3_trig_0_2 : std_logic;
signal un3_trig_0_1 : std_logic;
signal \g1_3_cascade_\ : std_logic;
signal \sEETrigInternal_prev_RNISEUGZ0_cascade_\ : std_logic;
signal \sTrigInternal_RNIOMLDZ0Z1_cascade_\ : std_logic;
signal \sTrigInternal_RNIOMLDZ0Z1\ : std_logic;
signal \sTrigInternal_RNOZ0Z_0_cascade_\ : std_logic;
signal un3_trig_0 : std_logic;
signal un3_trig_0_4 : std_logic;
signal un1_reset_rpi_inv_2_i_o3_8 : std_logic;
signal \un1_reset_rpi_inv_2_i_o3_18_cascade_\ : std_logic;
signal un3_trig_0_5 : std_logic;
signal un1_reset_rpi_inv_2_i_o3_13 : std_logic;
signal g0_2_0_3 : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_22_cascade_\ : std_logic;
signal \sbuttonModeStatusZ0\ : std_logic;
signal g1_0_0_3 : std_logic;
signal un1_reset_rpi_inv_2_i_o3_16 : std_logic;
signal g0_2_0_4 : std_logic;
signal g2_0_4 : std_logic;
signal g2_0_3 : std_logic;
signal \g1_0_1_1_cascade_\ : std_logic;
signal g1_0_4 : std_logic;
signal op_gt_op_gt_un13_striginternallto23_13 : std_logic;
signal \op_gt_op_gt_un13_striginternal_0_cascade_\ : std_logic;
signal \op_gt_op_gt_un13_striginternallto23_11_cascade_\ : std_logic;
signal op_gt_op_gt_un13_striginternallto23_16 : std_logic;
signal \sTrigInternalZ0\ : std_logic;
signal op_gt_op_gt_un13_striginternal_0 : std_logic;
signal \LED_ACQ_obuf_RNOZ0\ : std_logic;
signal op_gt_op_gt_un13_striginternallto23_18 : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \sCounterRAM_cry_0\ : std_logic;
signal \sCounterRAM_cry_1\ : std_logic;
signal \sCounterRAM_cry_2\ : std_logic;
signal \sCounterRAM_cry_3\ : std_logic;
signal \sCounterRAM_cry_4\ : std_logic;
signal \sCounterRAM_cry_5\ : std_logic;
signal \un1_spi_data_miso_0_sqmuxa_1_i_0_N_3_0\ : std_logic;
signal \sCounterRAM_cry_6\ : std_logic;
signal \sSPI_MSB0LSB1_RNIO3VPZ0Z1\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_16\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_14\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_15\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_150_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_36\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.div_clk_iZ0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.delay_clk_iZ0\ : std_logic;
signal g0_2_0_2 : std_logic;
signal g1_1 : std_logic;
signal \g2_0_2_cascade_\ : std_logic;
signal g1_0_3 : std_logic;
signal g0_2_0_1 : std_logic;
signal \g2_0_1_cascade_\ : std_logic;
signal g1_2 : std_logic;
signal g1_0_0_1 : std_logic;
signal g1_0_2 : std_logic;
signal g0_2_0_0 : std_logic;
signal \g2_0_0_cascade_\ : std_logic;
signal g1_0_0_0 : std_logic;
signal g1_0_1 : std_logic;
signal g0_2_0 : std_logic;
signal g1_4 : std_logic;
signal \g2_0_cascade_\ : std_logic;
signal \sEEPeriodZ0Z_0\ : std_logic;
signal \sEEPeriod_i_0\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \sEEPeriodZ0Z_1\ : std_logic;
signal \sEEPeriod_i_1\ : std_logic;
signal un4_speriod_cry_0 : std_logic;
signal \sEEPeriodZ0Z_2\ : std_logic;
signal \sEEPeriod_i_2\ : std_logic;
signal un4_speriod_cry_1 : std_logic;
signal \sEEPeriodZ0Z_3\ : std_logic;
signal \sEEPeriod_i_3\ : std_logic;
signal un4_speriod_cry_2 : std_logic;
signal \sEEPeriodZ0Z_4\ : std_logic;
signal \sEEPeriod_i_4\ : std_logic;
signal un4_speriod_cry_3 : std_logic;
signal \sEEPeriodZ0Z_5\ : std_logic;
signal \sEEPeriod_i_5\ : std_logic;
signal un4_speriod_cry_4 : std_logic;
signal \sEEPeriodZ0Z_6\ : std_logic;
signal \sEEPeriod_i_6\ : std_logic;
signal un4_speriod_cry_5 : std_logic;
signal \sEEPeriodZ0Z_7\ : std_logic;
signal \sEEPeriod_i_7\ : std_logic;
signal un4_speriod_cry_6 : std_logic;
signal un4_speriod_cry_7 : std_logic;
signal \sEEPeriod_i_8\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \sEEPeriod_i_9\ : std_logic;
signal un4_speriod_cry_8 : std_logic;
signal \sEEPeriod_i_10\ : std_logic;
signal un4_speriod_cry_9 : std_logic;
signal \sEEPeriod_i_11\ : std_logic;
signal un4_speriod_cry_10 : std_logic;
signal \sEEPeriod_i_12\ : std_logic;
signal un4_speriod_cry_11 : std_logic;
signal \sEEPeriod_i_13\ : std_logic;
signal un4_speriod_cry_12 : std_logic;
signal \sEEPeriod_i_14\ : std_logic;
signal un4_speriod_cry_13 : std_logic;
signal \sEEPeriod_i_15\ : std_logic;
signal un4_speriod_cry_14 : std_logic;
signal un4_speriod_cry_15 : std_logic;
signal \sEEPeriodZ0Z_16\ : std_logic;
signal \sEEPeriod_i_16\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \sEEPeriodZ0Z_17\ : std_logic;
signal \sEEPeriod_i_17\ : std_logic;
signal un4_speriod_cry_16 : std_logic;
signal \sEEPeriodZ0Z_18\ : std_logic;
signal \sEEPeriod_i_18\ : std_logic;
signal un4_speriod_cry_17 : std_logic;
signal \sEEPeriodZ0Z_19\ : std_logic;
signal \sEEPeriod_i_19\ : std_logic;
signal un4_speriod_cry_18 : std_logic;
signal \sEEPeriodZ0Z_20\ : std_logic;
signal \sEEPeriod_i_20\ : std_logic;
signal un4_speriod_cry_19 : std_logic;
signal \sEEPeriodZ0Z_21\ : std_logic;
signal \sEEPeriod_i_21\ : std_logic;
signal un4_speriod_cry_20 : std_logic;
signal \sEEPeriodZ0Z_22\ : std_logic;
signal \sEEPeriod_i_22\ : std_logic;
signal un4_speriod_cry_21 : std_logic;
signal \sEEPeriodZ0Z_23\ : std_logic;
signal \sEEPeriod_i_23\ : std_logic;
signal un4_speriod_cry_22 : std_logic;
signal un4_speriod_cry_23 : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal un1_reset_rpi_inv_2_i_o3_15 : std_logic;
signal un1_reset_rpi_inv_2_i_o3_11 : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_17\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \sCounter_cry_0\ : std_logic;
signal \sCounter_cry_1\ : std_logic;
signal \sCounter_cry_2\ : std_logic;
signal \sCounter_cry_3\ : std_logic;
signal \sCounter_cry_4\ : std_logic;
signal \sCounter_cry_5\ : std_logic;
signal \sCounter_cry_6\ : std_logic;
signal \sCounter_cry_7\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \sCounter_cry_8\ : std_logic;
signal \sCounter_cry_9\ : std_logic;
signal \sCounter_cry_10\ : std_logic;
signal \sCounter_cry_11\ : std_logic;
signal \sCounter_cry_12\ : std_logic;
signal \sCounter_cry_13\ : std_logic;
signal \sCounter_cry_14\ : std_logic;
signal \sCounter_cry_15\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \sCounter_cry_16\ : std_logic;
signal \sCounter_cry_17\ : std_logic;
signal \sCounter_cry_18\ : std_logic;
signal \sCounter_cry_19\ : std_logic;
signal \sCounter_cry_20\ : std_logic;
signal \sCounter_cry_21\ : std_logic;
signal \LED_ACQ_c_i\ : std_logic;
signal \sCounter_cry_22\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal un1_button_debounce_counter_cry_1 : std_logic;
signal un1_button_debounce_counter_cry_2 : std_logic;
signal un1_button_debounce_counter_cry_3 : std_logic;
signal un1_button_debounce_counter_cry_4 : std_logic;
signal \button_debounce_counterZ0Z_6\ : std_logic;
signal un1_button_debounce_counter_cry_5 : std_logic;
signal \button_debounce_counterZ0Z_7\ : std_logic;
signal un1_button_debounce_counter_cry_6 : std_logic;
signal \button_debounce_counterZ0Z_8\ : std_logic;
signal un1_button_debounce_counter_cry_7 : std_logic;
signal un1_button_debounce_counter_cry_8 : std_logic;
signal \button_debounce_counterZ0Z_9\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \button_debounce_counterZ0Z_10\ : std_logic;
signal un1_button_debounce_counter_cry_9 : std_logic;
signal \button_debounce_counterZ0Z_11\ : std_logic;
signal un1_button_debounce_counter_cry_10 : std_logic;
signal \button_debounce_counterZ0Z_12\ : std_logic;
signal un1_button_debounce_counter_cry_11 : std_logic;
signal \button_debounce_counterZ0Z_13\ : std_logic;
signal un1_button_debounce_counter_cry_12 : std_logic;
signal \button_debounce_counterZ0Z_14\ : std_logic;
signal un1_button_debounce_counter_cry_13 : std_logic;
signal \button_debounce_counterZ0Z_15\ : std_logic;
signal un1_button_debounce_counter_cry_14 : std_logic;
signal \button_debounce_counterZ0Z_16\ : std_logic;
signal un1_button_debounce_counter_cry_15 : std_logic;
signal un1_button_debounce_counter_cry_16 : std_logic;
signal \button_debounce_counterZ0Z_17\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \button_debounce_counterZ0Z_18\ : std_logic;
signal un1_button_debounce_counter_cry_17 : std_logic;
signal \button_debounce_counterZ0Z_19\ : std_logic;
signal un1_button_debounce_counter_cry_18 : std_logic;
signal \button_debounce_counterZ0Z_20\ : std_logic;
signal un1_button_debounce_counter_cry_19 : std_logic;
signal un1_button_debounce_counter_cry_20 : std_logic;
signal un1_button_debounce_counter_cry_21 : std_logic;
signal un1_button_debounce_counter_cry_22 : std_logic;
signal \un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO\ : std_logic;
signal \un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \button_debounce_counterZ0Z_23\ : std_logic;
signal \bfn_9_3_0_\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_158_7\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.N_158_7_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.falling_count_start_iZ0\ : std_logic;
signal un3_trig_0_0 : std_logic;
signal \un3_trig_0_0_cascade_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2\ : std_logic;
signal trig_ext_c : std_logic;
signal trig_rpi_c : std_logic;
signal trig_ft_c : std_logic;
signal \un8_trig_prev_0_c5_a0_0_0_cascade_\ : std_logic;
signal \un8_trig_prev_0_c4_a0_1_cascade_\ : std_logic;
signal \sEETrigCounterZ0Z_5\ : std_logic;
signal \sEETrigCounterZ0Z_6\ : std_logic;
signal \sEETrigCounterZ0Z_7\ : std_logic;
signal \un8_trig_prev_0_c7_a0_1_cascade_\ : std_logic;
signal un8_trig_prev_0_c4_a0_1 : std_logic;
signal \sEETrigCounterZ0Z_4\ : std_logic;
signal un8_trig_prev_0_c5_a0_0 : std_logic;
signal \sTrigCounter_i_0\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \sTrigCounter_i_1\ : std_logic;
signal un10_trig_prev_cry_0 : std_logic;
signal \sTrigCounter_i_2\ : std_logic;
signal un10_trig_prev_cry_1 : std_logic;
signal \sTrigCounter_i_3\ : std_logic;
signal un10_trig_prev_cry_2 : std_logic;
signal un10_trig_prev_4 : std_logic;
signal \sTrigCounter_i_4\ : std_logic;
signal un10_trig_prev_cry_3 : std_logic;
signal un10_trig_prev_5 : std_logic;
signal \sTrigCounter_i_5\ : std_logic;
signal un10_trig_prev_cry_4 : std_logic;
signal un10_trig_prev_6 : std_logic;
signal \sTrigCounter_i_6\ : std_logic;
signal un10_trig_prev_cry_5 : std_logic;
signal un10_trig_prev_7 : std_logic;
signal \sTrigCounter_i_7\ : std_logic;
signal un10_trig_prev_cry_6 : std_logic;
signal un10_trig_prev_cry_7 : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \sAddress_RNI9IH12_1Z0Z_1\ : std_logic;
signal \trig_prevZ0\ : std_logic;
signal un3_trig_0_3 : std_logic;
signal g1_0_0_2 : std_logic;
signal g1_0_0 : std_logic;
signal g1_0 : std_logic;
signal \sPeriod_prevZ0\ : std_logic;
signal \LED_MODE_c\ : std_logic;
signal \sTrigCounterZ0Z_4\ : std_logic;
signal \sTrigCounterZ0Z_3\ : std_logic;
signal \un1_sTrigCounter_ac0_0_0_cascade_\ : std_logic;
signal un1_reset_rpi_inv_2_i_o3_0_0 : std_logic;
signal \un1_sTrigCounter_ac0_0_2_0_cascade_\ : std_logic;
signal \un10_trig_prev_cry_7_THRU_CO\ : std_logic;
signal \sTrigCounterZ0Z_5\ : std_logic;
signal \un1_sTrigCounter_ac0_0_2\ : std_logic;
signal \un1_sTrigCounter_ac0_3_out_cascade_\ : std_logic;
signal \sTrigCounterZ0Z_2\ : std_logic;
signal g1_0_1_0 : std_logic;
signal g1_3_0 : std_logic;
signal \sEEPeriodZ0Z_10\ : std_logic;
signal \sEEPeriodZ0Z_11\ : std_logic;
signal \sEEPeriodZ0Z_12\ : std_logic;
signal \sEEPeriodZ0Z_13\ : std_logic;
signal \sEEPeriodZ0Z_14\ : std_logic;
signal \sEEPeriodZ0Z_15\ : std_logic;
signal \sEEPeriodZ0Z_8\ : std_logic;
signal \sEEPeriodZ0Z_9\ : std_logic;
signal op_gt_op_gt_un13_striginternallto23_12 : std_logic;
signal un1_reset_rpi_inv_2_i_o3_12 : std_logic;
signal op_gt_op_gt_un13_striginternallto23_15 : std_logic;
signal \sEETrigInternal_prevZ0\ : std_logic;
signal \N_5_0\ : std_logic;
signal \un4_speriod_cry_23_THRU_CO\ : std_logic;
signal \un1_reset_rpi_inv_2_i_1_1_0_cascade_\ : std_logic;
signal \un1_reset_rpi_inv_2_i_1_cascade_\ : std_logic;
signal \un1_sTrigCounter_ac0_0_4\ : std_logic;
signal \sTrigCounterZ0Z_6\ : std_logic;
signal \un1_sTrigCounter_axbxc7_m7_0_a2_2\ : std_logic;
signal un1_reset_rpi_inv_2_i_1 : std_logic;
signal \N_123\ : std_logic;
signal \sTrigCounterZ0Z_7\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal un1_spoff_cry_0 : std_logic;
signal un1_spoff_cry_1 : std_logic;
signal un1_spoff_cry_2 : std_logic;
signal un1_spoff_cry_3 : std_logic;
signal un1_spoff_cry_4 : std_logic;
signal un1_spoff_cry_5 : std_logic;
signal un1_spoff_cry_6 : std_logic;
signal un1_spoff_cry_7 : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal un1_spoff_cry_8 : std_logic;
signal un1_spoff_cry_9 : std_logic;
signal un1_spoff_cry_10 : std_logic;
signal un1_spoff_cry_11 : std_logic;
signal un1_spoff_cry_12 : std_logic;
signal un1_spoff_cry_13 : std_logic;
signal un1_spoff_cry_14 : std_logic;
signal un1_spoff_cry_15 : std_logic;
signal \sCounter_i_16\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \sCounter_i_17\ : std_logic;
signal un1_spoff_cry_16 : std_logic;
signal \sCounter_i_18\ : std_logic;
signal un1_spoff_cry_17 : std_logic;
signal \sCounter_i_19\ : std_logic;
signal un1_spoff_cry_18 : std_logic;
signal \sCounter_i_20\ : std_logic;
signal un1_spoff_cry_19 : std_logic;
signal \sCounter_i_21\ : std_logic;
signal un1_spoff_cry_20 : std_logic;
signal \sCounter_i_22\ : std_logic;
signal un1_spoff_cry_21 : std_logic;
signal \sCounter_i_23\ : std_logic;
signal un1_spoff_cry_22 : std_logic;
signal un1_spoff_cry_23 : std_logic;
signal \un4_spoff_cry_23_THRU_CO\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \N_1612_i\ : std_logic;
signal \sCounterRAMZ0Z_6\ : std_logic;
signal \sCounterRAMZ0Z_3\ : std_logic;
signal \button_debounce_counterZ0Z_21\ : std_logic;
signal \button_debounce_counterZ0Z_22\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_0\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_18\ : std_logic;
signal \button_debounce_counterZ0Z_4\ : std_logic;
signal \button_debounce_counterZ0Z_3\ : std_logic;
signal \button_debounce_counterZ0Z_5\ : std_logic;
signal \button_debounce_counterZ0Z_2\ : std_logic;
signal \sbuttonModeStatus_0_sqmuxa_13\ : std_logic;
signal \sEEDelayACQ_i_0\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \sEEDelayACQ_i_1\ : std_logic;
signal un4_sacqtime_cry_0 : std_logic;
signal \sEEDelayACQ_i_2\ : std_logic;
signal un4_sacqtime_cry_1 : std_logic;
signal \sEEDelayACQ_i_3\ : std_logic;
signal un4_sacqtime_cry_2 : std_logic;
signal \sEEDelayACQ_i_4\ : std_logic;
signal un4_sacqtime_cry_3 : std_logic;
signal \sEEDelayACQ_i_5\ : std_logic;
signal un4_sacqtime_cry_4 : std_logic;
signal \sEEDelayACQ_i_6\ : std_logic;
signal un4_sacqtime_cry_5 : std_logic;
signal \sEEDelayACQ_i_7\ : std_logic;
signal un4_sacqtime_cry_6 : std_logic;
signal un4_sacqtime_cry_7 : std_logic;
signal \sEEDelayACQ_i_8\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \sEEDelayACQ_i_9\ : std_logic;
signal un4_sacqtime_cry_8 : std_logic;
signal \sEEDelayACQ_i_10\ : std_logic;
signal un4_sacqtime_cry_9 : std_logic;
signal \sEEDelayACQ_i_11\ : std_logic;
signal un4_sacqtime_cry_10 : std_logic;
signal \sEEDelayACQ_i_12\ : std_logic;
signal un4_sacqtime_cry_11 : std_logic;
signal \sEEDelayACQ_i_13\ : std_logic;
signal un4_sacqtime_cry_12 : std_logic;
signal \sEEDelayACQ_i_14\ : std_logic;
signal un4_sacqtime_cry_13 : std_logic;
signal \sEEDelayACQ_i_15\ : std_logic;
signal un4_sacqtime_cry_14 : std_logic;
signal un4_sacqtime_cry_15 : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal un4_sacqtime_cry_16 : std_logic;
signal un4_sacqtime_cry_17 : std_logic;
signal un4_sacqtime_cry_18 : std_logic;
signal un4_sacqtime_cry_19 : std_logic;
signal op_gt_op_gt_un13_striginternallto23_8 : std_logic;
signal un4_sacqtime_cry_20 : std_logic;
signal un4_sacqtime_cry_21 : std_logic;
signal un4_sacqtime_cry_22 : std_logic;
signal un4_sacqtime_cry_23 : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \LED3_c_0\ : std_logic;
signal \bfn_10_2_0_\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3\ : std_logic;
signal \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4\ : std_logic;
signal \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_i6_3_cascade_\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_5\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.un23_i_ssn_3_cascade_\ : std_logic;
signal \spi_slave_inst.un23_i_ssn\ : std_logic;
signal \spi_slave_inst.un23_i_ssn_cascade_\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa\ : std_logic;
signal \spi_slave_inst.un23_i_ssn_3\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5\ : std_logic;
signal \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_6\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_1\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_2\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_11\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_12\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_3\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_14\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_15\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0\ : std_logic;
signal \bfn_10_6_0_\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.falling_count_start_i_i\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i\ : std_logic;
signal \sEETrigCounterZ0Z_3\ : std_logic;
signal un10_trig_prev_3 : std_logic;
signal \sEETrigCounterZ0Z_2\ : std_logic;
signal un10_trig_prev_2 : std_logic;
signal un10_trig_prev_0 : std_logic;
signal \sEETrigCounterZ0Z_0\ : std_logic;
signal \sEETrigCounterZ0Z_1\ : std_logic;
signal un10_trig_prev_1 : std_logic;
signal \spi_slave_inst.rx_done_reg3_iZ0\ : std_logic;
signal \spi_slave_inst.rx_ready_i_RNOZ0Z_0_cascade_\ : std_logic;
signal \spi_slave_inst.un4_tx_done_reg2_i_cascade_\ : std_logic;
signal \button_debounce_counterZ0Z_0\ : std_logic;
signal \button_debounce_counterZ0Z_1\ : std_logic;
signal \N_3089_g\ : std_logic;
signal \spi_mosi_ready_prevZ0Z2\ : std_logic;
signal \spi_mosi_ready_prevZ0\ : std_logic;
signal \spi_mosi_ready_prevZ0Z3\ : std_logic;
signal \spi_mosi_ready_prev3_RNILKERZ0_cascade_\ : std_logic;
signal \spi_slave_inst.tx_ready_iZ0\ : std_logic;
signal \sCounter_i_0\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \sCounter_i_1\ : std_logic;
signal un1_sacqtime_cry_0 : std_logic;
signal \sCounter_i_2\ : std_logic;
signal un1_sacqtime_cry_1 : std_logic;
signal \sCounter_i_3\ : std_logic;
signal un1_sacqtime_cry_2 : std_logic;
signal \sCounter_i_4\ : std_logic;
signal un1_sacqtime_cry_3 : std_logic;
signal \sCounter_i_5\ : std_logic;
signal un1_sacqtime_cry_4 : std_logic;
signal \sCounter_i_6\ : std_logic;
signal un1_sacqtime_cry_5 : std_logic;
signal \sCounter_i_7\ : std_logic;
signal un1_sacqtime_cry_6 : std_logic;
signal un1_sacqtime_cry_7 : std_logic;
signal \sCounter_i_8\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \sCounter_i_9\ : std_logic;
signal un1_sacqtime_cry_8 : std_logic;
signal \sCounter_i_10\ : std_logic;
signal un1_sacqtime_cry_9 : std_logic;
signal \sCounter_i_11\ : std_logic;
signal un1_sacqtime_cry_10 : std_logic;
signal \sCounter_i_12\ : std_logic;
signal un1_sacqtime_cry_11 : std_logic;
signal \sCounter_i_13\ : std_logic;
signal un1_sacqtime_cry_12 : std_logic;
signal \sCounter_i_14\ : std_logic;
signal un1_sacqtime_cry_13 : std_logic;
signal \sCounter_i_15\ : std_logic;
signal un1_sacqtime_cry_14 : std_logic;
signal un1_sacqtime_cry_15 : std_logic;
signal un1_sacqtime_cry_16_sf : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal un1_sacqtime_cry_17_sf : std_logic;
signal un1_sacqtime_cry_16 : std_logic;
signal un1_sacqtime_cry_18_sf : std_logic;
signal un1_sacqtime_cry_17 : std_logic;
signal un1_sacqtime_cry_19_sf : std_logic;
signal un1_sacqtime_cry_18 : std_logic;
signal un1_sacqtime_cry_20_sf : std_logic;
signal un1_sacqtime_cry_19 : std_logic;
signal un1_sacqtime_cry_21_sf : std_logic;
signal un1_sacqtime_cry_20 : std_logic;
signal un1_sacqtime_cry_22_sf : std_logic;
signal un1_sacqtime_cry_21 : std_logic;
signal un1_sacqtime_cry_23_sf : std_logic;
signal un1_sacqtime_cry_22 : std_logic;
signal un1_sacqtime_cry_23 : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \RAM_DATA_cl_10Z0Z_15\ : std_logic;
signal \N_106\ : std_logic;
signal \N_26\ : std_logic;
signal \N_76_i\ : std_logic;
signal \N_71_cascade_\ : std_logic;
signal \sEEDelayACQZ0Z_0\ : std_logic;
signal \sEEDelayACQZ0Z_1\ : std_logic;
signal \sEEDelayACQZ0Z_2\ : std_logic;
signal \sEEDelayACQZ0Z_3\ : std_logic;
signal \sEEDelayACQZ0Z_4\ : std_logic;
signal \sEEDelayACQZ0Z_5\ : std_logic;
signal \sEEDelayACQZ0Z_6\ : std_logic;
signal \sEEDelayACQZ0Z_7\ : std_logic;
signal \sEEDelayACQZ0Z_10\ : std_logic;
signal \sEEDelayACQZ0Z_11\ : std_logic;
signal \sEEDelayACQZ0Z_12\ : std_logic;
signal \sEEDelayACQZ0Z_13\ : std_logic;
signal \sEEDelayACQZ0Z_14\ : std_logic;
signal \sEEDelayACQZ0Z_15\ : std_logic;
signal \sEEDelayACQZ0Z_8\ : std_logic;
signal \sEEDelayACQZ0Z_9\ : std_logic;
signal \sAddress_RNIA6242Z0Z_0\ : std_logic;
signal \N_99_cascade_\ : std_logic;
signal \RAM_DATA_cl_12Z0Z_15\ : std_logic;
signal \N_94_cascade_\ : std_logic;
signal \RAM_DATA_cl_11Z0Z_15\ : std_logic;
signal \N_104_cascade_\ : std_logic;
signal \RAM_DATA_cl_14Z0Z_15\ : std_logic;
signal \sDAC_dataZ0Z_2\ : std_logic;
signal \spi_slave_inst.rx_data_count_neg_sclk_i6\ : std_logic;
signal \INVspi_slave_inst.rx_done_neg_sclk_iC_net\ : std_logic;
signal \spi_slave_inst.rx_done_neg_sclk_iZ0\ : std_logic;
signal \spi_slave_inst.rx_done_pos_sclk_iZ0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0\ : std_logic;
signal \spi_master_inst.sclk_gen_u0.spi_start_iZ0\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3_cascade_\ : std_logic;
signal \spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0\ : std_logic;
signal \spi_slave_inst.N_1394\ : std_logic;
signal \spi_slave_inst.N_1397_cascade_\ : std_logic;
signal \spi_slave_inst.tx_done_reg1_iZ0\ : std_logic;
signal \spi_slave_inst.tx_done_reg2_iZ0\ : std_logic;
signal \spi_slave_inst.tx_done_reg3_iZ0\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_0\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_7\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_5\ : std_logic;
signal \spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_1\ : std_logic;
signal \spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_2\ : std_logic;
signal \spi_slave_inst.txdata_reg_iZ0Z_6\ : std_logic;
signal \N_206\ : std_logic;
signal \N_206_cascade_\ : std_logic;
signal \sAddress_RNIA6242_1Z0Z_0\ : std_logic;
signal \spi_mosi_ready64_prevZ0Z2\ : std_logic;
signal \spi_mosi_ready64_prevZ0\ : std_logic;
signal \spi_mosi_ready64_prevZ0Z3\ : std_logic;
signal spi_mosi_ready : std_logic;
signal \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_\ : std_logic;
signal \LED3_c_i\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_0\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_1\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_2\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_5\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_6\ : std_logic;
signal \spi_slave_inst.data_in_reg_iZ0Z_7\ : std_logic;
signal \spi_slave_inst.un4_i_wr\ : std_logic;
signal \RAM_DATA_in_6\ : std_logic;
signal \RAM_DATA_in_14\ : std_logic;
signal \spi_data_misoZ0Z_6\ : std_logic;
signal \RAM_DATA_in_7\ : std_logic;
signal \RAM_DATA_in_15\ : std_logic;
signal \spi_data_misoZ0Z_7\ : std_logic;
signal \RAM_nWE_0_i\ : std_logic;
signal \sADC_clk_prevZ0\ : std_logic;
signal \ADC_clk_c\ : std_logic;
signal \N_127\ : std_logic;
signal \N_1470_i\ : std_logic;
signal \N_86\ : std_logic;
signal \sRead_dataZ0\ : std_logic;
signal \sCounterRAMZ0Z_5\ : std_logic;
signal \sCounterRAMZ0Z_4\ : std_logic;
signal \sCounterRAMZ0Z_7\ : std_logic;
signal \sCounterRAMZ0Z_0\ : std_logic;
signal \sCounterRAMZ0Z_2\ : std_logic;
signal \sCounterRAMZ0Z_1\ : std_logic;
signal \spi_data_miso_0_sqmuxa_2_i_o2_5_cascade_\ : std_logic;
signal spi_data_miso_0_sqmuxa_2_i_o2_4 : std_logic;
signal \N_75_cascade_\ : std_logic;
signal \sSPI_MSB0LSBZ0Z1\ : std_logic;
signal \spi_mosi_ready_prev3_RNILKERZ0\ : std_logic;
signal \N_88\ : std_logic;
signal \N_88_cascade_\ : std_logic;
signal \N_28\ : std_logic;
signal \N_93_cascade_\ : std_logic;
signal \RAM_DATA_cl_9Z0Z_15\ : std_logic;
signal \N_98_cascade_\ : std_logic;
signal \RAM_DATA_clZ0Z_15\ : std_logic;
signal \N_96_cascade_\ : std_logic;
signal \RAM_DATA_cl_8Z0Z_15\ : std_logic;
signal \sRAM_pointer_readZ0Z_14\ : std_logic;
signal \RAM_ADD_c_14\ : std_logic;
signal \sRAM_pointer_readZ0Z_15\ : std_logic;
signal \RAM_ADD_c_15\ : std_logic;
signal \sRAM_pointer_readZ0Z_16\ : std_logic;
signal \RAM_ADD_c_16\ : std_logic;
signal \sRAM_pointer_readZ0Z_17\ : std_logic;
signal \RAM_ADD_c_17\ : std_logic;
signal \sRAM_pointer_readZ0Z_18\ : std_logic;
signal \RAM_ADD_c_18\ : std_logic;
signal \sRAM_pointer_readZ0Z_2\ : std_logic;
signal \RAM_ADD_c_2\ : std_logic;
signal \sRAM_pointer_readZ0Z_3\ : std_logic;
signal \RAM_ADD_c_3\ : std_logic;
signal \sRAM_pointer_readZ0Z_4\ : std_logic;
signal \RAM_ADD_c_4\ : std_logic;
signal \sRAM_pointer_readZ0Z_5\ : std_logic;
signal \RAM_ADD_c_5\ : std_logic;
signal \sRAM_pointer_readZ0Z_6\ : std_logic;
signal \RAM_ADD_c_6\ : std_logic;
signal \sRAM_pointer_readZ0Z_7\ : std_logic;
signal \RAM_ADD_c_7\ : std_logic;
signal \sRAM_pointer_readZ0Z_8\ : std_logic;
signal \RAM_ADD_c_8\ : std_logic;
signal \sRAM_pointer_readZ0Z_9\ : std_logic;
signal \RAM_ADD_c_9\ : std_logic;
signal \N_102\ : std_logic;
signal \RAM_DATA_cl_15Z0Z_15\ : std_logic;
signal spi_sclk_ft_c : std_logic;
signal spi_sclk : std_logic;
signal \spi_slave_inst.rx_done_reg1_iZ0\ : std_logic;
signal \spi_slave_inst.rx_done_reg2_iZ0\ : std_logic;
signal \spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_10\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_13\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_4\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_5\ : std_logic;
signal \sDAC_dataZ0Z_0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_0\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_7\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_8\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.data_inZ0Z_9\ : std_logic;
signal \spi_master_inst.spi_data_path_u1.tx_ready_iZ0\ : std_logic;
signal \un1_spointer11_5_0_2_cascade_\ : std_logic;
signal \sAddress_RNIA6242_0Z0Z_2\ : std_logic;
signal \sDAC_mem_23_1_sqmuxa\ : std_logic;
signal \N_275_cascade_\ : std_logic;
signal \N_360_cascade_\ : std_logic;
signal \N_269\ : std_logic;
signal \N_132\ : std_logic;
signal \sAddress_RNIA6242_0Z0Z_0\ : std_logic;
signal un1_spointer11_7_0_tz : std_logic;
signal \un1_spointer11_7_0_tz_cascade_\ : std_logic;
signal \sAddress_RNID9242Z0Z_3\ : std_logic;
signal \spi_slave_inst.un1_spointer11_2_0_a2_0_6_4\ : std_logic;
signal \spi_slave_inst.un1_spointer11_2_0_a2_0_6_5_cascade_\ : std_logic;
signal un1_spointer11_2_0 : std_logic;
signal \N_285_cascade_\ : std_logic;
signal \sPointerZ0Z_0\ : std_logic;
signal \N_116_cascade_\ : std_logic;
signal \N_159\ : std_logic;
signal \N_117_cascade_\ : std_logic;
signal \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1\ : std_logic;
signal \sEETrigInternalZ0\ : std_logic;
signal \sEEPoffZ0Z_0\ : std_logic;
signal \sEEPoffZ0Z_1\ : std_logic;
signal \sEEPoffZ0Z_2\ : std_logic;
signal \sEEPoffZ0Z_3\ : std_logic;
signal \sEEPoffZ0Z_4\ : std_logic;
signal \sEEPoffZ0Z_5\ : std_logic;
signal \sEEPoffZ0Z_6\ : std_logic;
signal \sEEPoffZ0Z_7\ : std_logic;
signal \sEEPoffZ0Z_10\ : std_logic;
signal \sEEPoffZ0Z_11\ : std_logic;
signal \sEEPoffZ0Z_12\ : std_logic;
signal \sEEPoffZ0Z_13\ : std_logic;
signal \sEEPoffZ0Z_14\ : std_logic;
signal \sEEPoffZ0Z_15\ : std_logic;
signal \sEEPoffZ0Z_8\ : std_logic;
signal \sEEPoffZ0Z_9\ : std_logic;
signal \sAddress_RNIA6242_1Z0Z_2\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \sCounterADC_cry_0\ : std_logic;
signal \sCounterADC_cry_1\ : std_logic;
signal \sCounterADC_cry_2\ : std_logic;
signal \sCounterADC_cry_3\ : std_logic;
signal \sCounterADC_cry_4\ : std_logic;
signal \sCounterADC_cry_5\ : std_logic;
signal \sCounterADC_cry_6\ : std_logic;
signal \RAM_DATA_in_8\ : std_logic;
signal \RAM_DATA_in_0\ : std_logic;
signal \spi_data_misoZ0Z_0\ : std_logic;
signal \RAM_DATA_in_9\ : std_logic;
signal \RAM_DATA_in_1\ : std_logic;
signal \spi_data_misoZ0Z_1\ : std_logic;
signal \RAM_DATA_in_10\ : std_logic;
signal \RAM_DATA_in_2\ : std_logic;
signal \spi_data_misoZ0Z_2\ : std_logic;
signal \RAM_DATA_in_11\ : std_logic;
signal \RAM_DATA_in_3\ : std_logic;
signal \spi_data_misoZ0Z_3\ : std_logic;
signal \RAM_DATA_in_12\ : std_logic;
signal \RAM_DATA_in_4\ : std_logic;
signal \spi_data_misoZ0Z_4\ : std_logic;
signal \un4_sacqtime_cry_23_c_RNITTSZ0Z3\ : std_logic;
signal \RAM_DATA_in_5\ : std_logic;
signal \N_75\ : std_logic;
signal \RAM_DATA_in_13\ : std_logic;
signal \spi_data_misoZ0Z_5\ : std_logic;
signal \N_6\ : std_logic;
signal \sRAM_pointer_readZ0Z_0\ : std_logic;
signal \RAM_ADD_c_0\ : std_logic;
signal \reset_rpi_ibuf_RNI7JCVZ0\ : std_logic;
signal \sRAM_ADD_0_sqmuxa_i_0\ : std_logic;
signal \sRAM_pointer_readZ0Z_1\ : std_logic;
signal \RAM_ADD_c_1\ : std_logic;
signal \sRAM_pointer_readZ0Z_10\ : std_logic;
signal \RAM_ADD_c_10\ : std_logic;
signal \sRAM_pointer_readZ0Z_11\ : std_logic;
signal \RAM_ADD_c_11\ : std_logic;
signal \sRAM_pointer_readZ0Z_12\ : std_logic;
signal \RAM_ADD_c_12\ : std_logic;
signal \sRAM_pointer_readZ0Z_13\ : std_logic;
signal \RAM_ADD_c_13\ : std_logic;
signal \N_67_i\ : std_logic;
signal \ADC3_c\ : std_logic;
signal \RAM_DATA_1Z0Z_3\ : std_logic;
signal \ADC0_c\ : std_logic;
signal \RAM_DATA_1Z0Z_0\ : std_logic;
signal \ADC5_c\ : std_logic;
signal \RAM_DATA_1Z0Z_5\ : std_logic;
signal \ADC1_c\ : std_logic;
signal \RAM_DATA_1Z0Z_1\ : std_logic;
signal \ADC7_c\ : std_logic;
signal \RAM_DATA_1Z0Z_8\ : std_logic;
signal \ADC8_c\ : std_logic;
signal \RAM_DATA_1Z0Z_9\ : std_logic;
signal \RAM_DATA_1Z0Z_15\ : std_logic;
signal \RAM_DATA_1Z0Z_7\ : std_logic;
signal \RAM_DATA_cl_1Z0Z_15\ : std_logic;
signal \N_100\ : std_logic;
signal \RAM_DATA_cl_13Z0Z_15\ : std_logic;
signal \N_97\ : std_logic;
signal \RAM_DATA_cl_2Z0Z_15\ : std_logic;
signal \N_101\ : std_logic;
signal \N_103\ : std_logic;
signal \RAM_DATA_cl_3Z0Z_15\ : std_logic;
signal spi_mosi_ft_c : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6\ : std_logic;
signal \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7\ : std_logic;
signal spi_sclk_g : std_logic;
signal \spi_slave_inst.spi_cs_iZ0\ : std_logic;
signal \sDAC_mem_23Z0Z_2\ : std_logic;
signal \sDAC_mem_22Z0Z_2\ : std_logic;
signal \sDAC_mem_23Z0Z_3\ : std_logic;
signal \sDAC_mem_22Z0Z_3\ : std_logic;
signal \sDAC_mem_23Z0Z_4\ : std_logic;
signal \sDAC_mem_22Z0Z_4\ : std_logic;
signal \N_291_cascade_\ : std_logic;
signal \sEEPonPoff_1_sqmuxa\ : std_logic;
signal \sAddressZ0Z_6\ : std_logic;
signal \sAddressZ0Z_7\ : std_logic;
signal \sEEPonPoff_1_sqmuxa_0_a2_1\ : std_logic;
signal \sEEPon_1_sqmuxa\ : std_logic;
signal \N_291\ : std_logic;
signal \sDAC_mem_33_1_sqmuxa\ : std_logic;
signal \sDAC_mem_17_1_sqmuxa\ : std_logic;
signal \sDAC_mem_32_1_sqmuxa\ : std_logic;
signal \N_141\ : std_logic;
signal \sEETrigCounter_1_sqmuxa\ : std_logic;
signal \N_1480_cascade_\ : std_logic;
signal un1_spointer11_5_0_2 : std_logic;
signal \sAddress_RNIA6242_2Z0Z_2\ : std_logic;
signal \N_280_cascade_\ : std_logic;
signal \sDAC_mem_19_1_sqmuxa\ : std_logic;
signal \sDAC_mem_19Z0Z_4\ : std_logic;
signal \sDAC_mem_18Z0Z_4\ : std_logic;
signal \sDAC_mem_19Z0Z_5\ : std_logic;
signal \sDAC_mem_18Z0Z_5\ : std_logic;
signal \sDAC_mem_19Z0Z_6\ : std_logic;
signal \sDAC_mem_18Z0Z_6\ : std_logic;
signal \sAddress_RNIA6242Z0Z_2\ : std_logic;
signal \ADC4_c\ : std_logic;
signal \RAM_DATA_1Z0Z_4\ : std_logic;
signal \ADC6_c\ : std_logic;
signal \RAM_DATA_1Z0Z_6\ : std_logic;
signal \ADC9_c\ : std_logic;
signal \RAM_DATA_1Z0Z_10\ : std_logic;
signal top_tour1_c : std_logic;
signal \RAM_DATA_1Z0Z_11\ : std_logic;
signal top_tour2_c : std_logic;
signal \RAM_DATA_1Z0Z_12\ : std_logic;
signal \sTrigCounterZ0Z_0\ : std_logic;
signal \RAM_DATA_1Z0Z_13\ : std_logic;
signal \sTrigCounterZ0Z_1\ : std_logic;
signal \RAM_DATA_1Z0Z_14\ : std_logic;
signal \ADC2_c\ : std_logic;
signal \RAM_DATA_1Z0Z_2\ : std_logic;
signal \N_31_i\ : std_logic;
signal \N_107_cascade_\ : std_logic;
signal \RAM_DATA_cl_5Z0Z_15\ : std_logic;
signal \N_108_cascade_\ : std_logic;
signal \RAM_DATA_cl_6Z0Z_15\ : std_logic;
signal \LED3_c\ : std_logic;
signal \un4_sacqtime_cry_23_THRU_CO\ : std_logic;
signal \N_95_cascade_\ : std_logic;
signal \un1_sacqtime_cry_23_THRU_CO\ : std_logic;
signal \RAM_DATA_cl_7Z0Z_15\ : std_logic;
signal \RAM_DATA_cl_4Z0Z_15\ : std_logic;
signal \N_71\ : std_logic;
signal \N_105\ : std_logic;
signal \sRAM_pointer_writeZ0Z_0\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \sRAM_pointer_writeZ0Z_1\ : std_logic;
signal \sRAM_pointer_write_cry_0\ : std_logic;
signal \sRAM_pointer_writeZ0Z_2\ : std_logic;
signal \sRAM_pointer_write_cry_1\ : std_logic;
signal \sRAM_pointer_writeZ0Z_3\ : std_logic;
signal \sRAM_pointer_write_cry_2\ : std_logic;
signal \sRAM_pointer_writeZ0Z_4\ : std_logic;
signal \sRAM_pointer_write_cry_3\ : std_logic;
signal \sRAM_pointer_writeZ0Z_5\ : std_logic;
signal \sRAM_pointer_write_cry_4\ : std_logic;
signal \sRAM_pointer_writeZ0Z_6\ : std_logic;
signal \sRAM_pointer_write_cry_5\ : std_logic;
signal \sRAM_pointer_writeZ0Z_7\ : std_logic;
signal \sRAM_pointer_write_cry_6\ : std_logic;
signal \sRAM_pointer_write_cry_7\ : std_logic;
signal \sRAM_pointer_writeZ0Z_8\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \sRAM_pointer_writeZ0Z_9\ : std_logic;
signal \sRAM_pointer_write_cry_8\ : std_logic;
signal \sRAM_pointer_writeZ0Z_10\ : std_logic;
signal \sRAM_pointer_write_cry_9\ : std_logic;
signal \sRAM_pointer_writeZ0Z_11\ : std_logic;
signal \sRAM_pointer_write_cry_10\ : std_logic;
signal \sRAM_pointer_writeZ0Z_12\ : std_logic;
signal \sRAM_pointer_write_cry_11\ : std_logic;
signal \sRAM_pointer_writeZ0Z_13\ : std_logic;
signal \sRAM_pointer_write_cry_12\ : std_logic;
signal \sRAM_pointer_writeZ0Z_14\ : std_logic;
signal \sRAM_pointer_write_cry_13\ : std_logic;
signal \sRAM_pointer_writeZ0Z_15\ : std_logic;
signal \sRAM_pointer_write_cry_14\ : std_logic;
signal \sRAM_pointer_write_cry_15\ : std_logic;
signal \sRAM_pointer_writeZ0Z_16\ : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal \sRAM_pointer_writeZ0Z_17\ : std_logic;
signal \sRAM_pointer_write_cry_16\ : std_logic;
signal \sEEPointerResetZ0\ : std_logic;
signal \sRAM_pointer_write_cry_17\ : std_logic;
signal \sRAM_pointer_writeZ0Z_18\ : std_logic;
signal \N_26_g\ : std_logic;
signal spi_cs_ft_c : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_\ : std_logic;
signal \spi_slave_inst.spi_csZ0\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_\ : std_logic;
signal \spi_slave_inst.tx_done_neg_sclk_iZ0\ : std_logic;
signal \INVspi_slave_inst.tx_done_neg_sclk_iC_net\ : std_logic;
signal spi_miso_flash_c : std_logic;
signal spi_miso_rpi_c : std_logic;
signal \sDAC_data_2_13_bm_1_3_cascade_\ : std_logic;
signal \sDAC_mem_6Z0Z_0\ : std_logic;
signal \sDAC_mem_38Z0Z_1\ : std_logic;
signal \sDAC_data_2_13_bm_1_4_cascade_\ : std_logic;
signal \sDAC_mem_6Z0Z_1\ : std_logic;
signal \sDAC_mem_6Z0Z_2\ : std_logic;
signal \sDAC_data_2_13_bm_1_5_cascade_\ : std_logic;
signal \sDAC_data_2_13_am_1_5_cascade_\ : std_logic;
signal \sDAC_mem_4Z0Z_2\ : std_logic;
signal \sDAC_data_2_13_am_1_6_cascade_\ : std_logic;
signal \sDAC_mem_4Z0Z_3\ : std_logic;
signal \sDAC_mem_4Z0Z_4\ : std_logic;
signal \sDAC_data_2_13_am_1_7_cascade_\ : std_logic;
signal \sDAC_mem_2Z0Z_0\ : std_logic;
signal \sDAC_data_2_6_bm_1_3_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_0\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_5_cascade_\ : std_logic;
signal \sDAC_data_2_20_am_1_5_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_5_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_5_cascade_\ : std_logic;
signal \sDAC_data_2_32_ns_1_5\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_5\ : std_logic;
signal \sDAC_data_2_14_ns_1_5_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_5_cascade_\ : std_logic;
signal \sDAC_data_2_41_ns_1_5\ : std_logic;
signal \sDAC_data_2_5_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_5\ : std_logic;
signal \sDAC_mem_2Z0Z_2\ : std_logic;
signal \sDAC_data_2_6_bm_1_5_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_5\ : std_logic;
signal \sDAC_data_2_20_am_1_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_7\ : std_logic;
signal \sDAC_mem_33Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_27Z0Z_8_cascade_\ : std_logic;
signal \sDAC_mem_32Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_8\ : std_logic;
signal \sDAC_mem_1Z0Z_5\ : std_logic;
signal \sDAC_mem_33Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_9_cascade_\ : std_logic;
signal \sDAC_mem_32Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_27Z0Z_9\ : std_logic;
signal \sDAC_mem_1Z0Z_6\ : std_logic;
signal \sDAC_mem_2Z0Z_6\ : std_logic;
signal \sDAC_data_2_6_bm_1_9_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_6\ : std_logic;
signal \sDAC_mem_33Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_4_cascade_\ : std_logic;
signal \sDAC_mem_1Z0Z_1\ : std_logic;
signal \sDAC_mem_32Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_27Z0Z_4\ : std_logic;
signal \sDAC_mem_33Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_5_cascade_\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_5\ : std_logic;
signal \sDAC_mem_32Z0Z_2\ : std_logic;
signal \sDAC_mem_1Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_27Z0Z_5\ : std_logic;
signal \op_le_op_le_un15_sdacdynlt4_cascade_\ : std_logic;
signal un17_sdacdyn_0 : std_logic;
signal \sDAC_mem_10Z0Z_7\ : std_logic;
signal \sDAC_mem_19Z0Z_7\ : std_logic;
signal \sDAC_mem_18Z0Z_7\ : std_logic;
signal \sDAC_mem_19Z0Z_0\ : std_logic;
signal \sDAC_mem_18Z0Z_0\ : std_logic;
signal \sDAC_mem_19Z0Z_1\ : std_logic;
signal \sDAC_mem_18Z0Z_1\ : std_logic;
signal \sDAC_mem_19Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_5\ : std_logic;
signal \sDAC_mem_18Z0Z_2\ : std_logic;
signal \sDAC_mem_18_1_sqmuxa\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_5_cascade_\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_5\ : std_logic;
signal \sDAC_data_2_24_ns_1_5\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_6\ : std_logic;
signal \sDAC_mem_12Z0Z_2\ : std_logic;
signal \sDAC_mem_12Z0Z_3\ : std_logic;
signal \sDAC_mem_31_1_sqmuxa\ : std_logic;
signal \sCounterADCZ0Z_3\ : std_logic;
signal \sCounterADCZ0Z_2\ : std_logic;
signal \sEEADC_freqZ0Z_2\ : std_logic;
signal \sEEADC_freqZ0Z_3\ : std_logic;
signal \sCounterADCZ0Z_5\ : std_logic;
signal \sCounterADCZ0Z_4\ : std_logic;
signal \sEEADC_freqZ0Z_4\ : std_logic;
signal \sEEADC_freqZ0Z_5\ : std_logic;
signal \sCounterADCZ0Z_6\ : std_logic;
signal \sCounterADCZ0Z_7\ : std_logic;
signal un7_spon_0 : std_logic;
signal \sEEACQZ0Z_0\ : std_logic;
signal \sEEACQ_i_0\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \sEEACQZ0Z_1\ : std_logic;
signal un7_spon_1 : std_logic;
signal \sEEACQ_i_1\ : std_logic;
signal un5_sdacdyn_cry_0 : std_logic;
signal un7_spon_2 : std_logic;
signal \sEEACQZ0Z_2\ : std_logic;
signal \sEEACQ_i_2\ : std_logic;
signal un5_sdacdyn_cry_1 : std_logic;
signal un7_spon_3 : std_logic;
signal \sEEACQZ0Z_3\ : std_logic;
signal \sEEACQ_i_3\ : std_logic;
signal un5_sdacdyn_cry_2 : std_logic;
signal \sEEACQZ0Z_4\ : std_logic;
signal \sEEACQ_i_4\ : std_logic;
signal un5_sdacdyn_cry_3 : std_logic;
signal un7_spon_5 : std_logic;
signal \sEEACQZ0Z_5\ : std_logic;
signal \sEEACQ_i_5\ : std_logic;
signal un5_sdacdyn_cry_4 : std_logic;
signal un7_spon_6 : std_logic;
signal \sEEACQZ0Z_6\ : std_logic;
signal \sEEACQ_i_6\ : std_logic;
signal un5_sdacdyn_cry_5 : std_logic;
signal un7_spon_7 : std_logic;
signal \sEEACQZ0Z_7\ : std_logic;
signal \sEEACQ_i_7\ : std_logic;
signal un5_sdacdyn_cry_6 : std_logic;
signal un5_sdacdyn_cry_7 : std_logic;
signal un7_spon_8 : std_logic;
signal \sEEACQZ0Z_8\ : std_logic;
signal \sEEACQ_i_8\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal un7_spon_9 : std_logic;
signal \sEEACQZ0Z_9\ : std_logic;
signal \sEEACQ_i_9\ : std_logic;
signal un5_sdacdyn_cry_8 : std_logic;
signal un7_spon_10 : std_logic;
signal \sEEACQZ0Z_10\ : std_logic;
signal \sEEACQ_i_10\ : std_logic;
signal un5_sdacdyn_cry_9 : std_logic;
signal un7_spon_11 : std_logic;
signal \sEEACQZ0Z_11\ : std_logic;
signal \sEEACQ_i_11\ : std_logic;
signal un5_sdacdyn_cry_10 : std_logic;
signal \sEEACQZ0Z_12\ : std_logic;
signal un7_spon_12 : std_logic;
signal \sEEACQ_i_12\ : std_logic;
signal un5_sdacdyn_cry_11 : std_logic;
signal un7_spon_13 : std_logic;
signal \sEEACQZ0Z_13\ : std_logic;
signal \sEEACQ_i_13\ : std_logic;
signal un5_sdacdyn_cry_12 : std_logic;
signal un7_spon_14 : std_logic;
signal \sEEACQZ0Z_14\ : std_logic;
signal \sEEACQ_i_14\ : std_logic;
signal un5_sdacdyn_cry_13 : std_logic;
signal un7_spon_15 : std_logic;
signal \sEEACQZ0Z_15\ : std_logic;
signal \sEEACQ_i_15\ : std_logic;
signal un5_sdacdyn_cry_14 : std_logic;
signal un5_sdacdyn_cry_15 : std_logic;
signal un7_spon_16 : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal un7_spon_17 : std_logic;
signal un5_sdacdyn_cry_16 : std_logic;
signal un7_spon_18 : std_logic;
signal un5_sdacdyn_cry_17 : std_logic;
signal un7_spon_19 : std_logic;
signal un5_sdacdyn_cry_18 : std_logic;
signal un7_spon_20 : std_logic;
signal un5_sdacdyn_cry_19 : std_logic;
signal un7_spon_21 : std_logic;
signal un5_sdacdyn_cry_20 : std_logic;
signal un7_spon_22 : std_logic;
signal un5_sdacdyn_cry_21 : std_logic;
signal un7_spon_23 : std_logic;
signal un5_sdacdyn_cry_22 : std_logic;
signal un5_sdacdyn_cry_23 : std_logic;
signal un17_sdacdyn_1 : std_logic;
signal \N_1479\ : std_logic;
signal un7_spon_4 : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \sDAC_mem_24Z0Z_3\ : std_logic;
signal \sDAC_mem_24Z0Z_6\ : std_logic;
signal \sDAC_mem_17Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_5\ : std_logic;
signal \sDAC_mem_16Z0Z_2\ : std_logic;
signal \sDAC_mem_pointerZ0Z_6\ : std_logic;
signal \sDAC_mem_pointerZ0Z_7\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0\ : std_logic;
signal \bfn_15_2_0_\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1\ : std_logic;
signal \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_i6\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2\ : std_logic;
signal \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3\ : std_logic;
signal \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4\ : std_logic;
signal \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3\ : std_logic;
signal \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4\ : std_logic;
signal \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5\ : std_logic;
signal \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\ : std_logic;
signal \sDAC_mem_34Z0Z_0\ : std_logic;
signal \sDAC_mem_34Z0Z_2\ : std_logic;
signal \sDAC_mem_34Z0Z_6\ : std_logic;
signal \sDAC_mem_7Z0Z_0\ : std_logic;
signal \sDAC_mem_7Z0Z_1\ : std_logic;
signal \sDAC_mem_7Z0Z_2\ : std_logic;
signal \sDAC_mem_5Z0Z_2\ : std_logic;
signal \sDAC_mem_5Z0Z_3\ : std_logic;
signal \sDAC_mem_5Z0Z_4\ : std_logic;
signal \sDAC_mem_2_1_sqmuxa\ : std_logic;
signal \sDAC_mem_5_1_sqmuxa\ : std_logic;
signal \sDAC_mem_7_1_sqmuxa\ : std_logic;
signal \N_279\ : std_logic;
signal \N_279_cascade_\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_7\ : std_logic;
signal \sDAC_data_2_14_ns_1_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_7\ : std_logic;
signal \sDAC_data_2_41_ns_1_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_7\ : std_logic;
signal \sDAC_data_2_7_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_7\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_9_cascade_\ : std_logic;
signal \sDAC_data_2_20_am_1_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_9\ : std_logic;
signal \sDAC_mem_17Z0Z_4\ : std_logic;
signal \sDAC_mem_16Z0Z_4\ : std_logic;
signal \sDAC_mem_17Z0Z_5\ : std_logic;
signal \sDAC_mem_16Z0Z_5\ : std_logic;
signal \sDAC_mem_17Z0Z_6\ : std_logic;
signal \sDAC_mem_16Z0Z_6\ : std_logic;
signal \bfn_15_10_0_\ : std_logic;
signal \sDAC_mem_pointer_0_cry_1\ : std_logic;
signal \sDAC_mem_pointer_0_cry_2\ : std_logic;
signal \sDAC_mem_pointer_0_cry_3\ : std_logic;
signal \sDAC_mem_pointer_0_cry_4\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_10\ : std_logic;
signal \sDAC_data_2_24_ns_1_10\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_10_cascade_\ : std_logic;
signal \sDAC_data_2_20_am_1_10_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_10\ : std_logic;
signal \sDAC_mem_28Z0Z_6\ : std_logic;
signal \sDAC_dataZ0Z_1\ : std_logic;
signal \sDAC_dataZ0Z_11\ : std_logic;
signal \sDAC_dataZ0Z_12\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \sDAC_dataZ0Z_13\ : std_logic;
signal \sDAC_dataZ0Z_14\ : std_logic;
signal \GNDG0\ : std_logic;
signal \sDAC_dataZ0Z_15\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_8_cascade_\ : std_logic;
signal \sDAC_data_2_39_ns_1_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_32Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_8\ : std_logic;
signal \sDAC_mem_31Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_8\ : std_logic;
signal \sDAC_mem_24Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_9\ : std_logic;
signal \sDAC_data_RNO_32Z0Z_9\ : std_logic;
signal \sDAC_data_2_39_ns_1_9\ : std_logic;
signal \sDAC_mem_26Z0Z_0\ : std_logic;
signal \sDAC_mem_26Z0Z_5\ : std_logic;
signal \sDAC_mem_26Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_9\ : std_logic;
signal \sDAC_data_2_24_ns_1_9\ : std_logic;
signal \sCounterADCZ0Z_1\ : std_logic;
signal \sCounterADCZ0Z_0\ : std_logic;
signal \un11_sacqtime_NE_3\ : std_logic;
signal \un11_sacqtime_NE_2\ : std_logic;
signal \un11_sacqtime_NE_0_0_cascade_\ : std_logic;
signal \un11_sacqtime_NE_1\ : std_logic;
signal \un11_sacqtime_NE_0\ : std_logic;
signal \sDAC_mem_31Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_9\ : std_logic;
signal \sDAC_mem_29Z0Z_5\ : std_logic;
signal \sDAC_mem_29Z0Z_6\ : std_logic;
signal \sDAC_mem_29_1_sqmuxa\ : std_logic;
signal \sDAC_mem_29Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_6\ : std_logic;
signal \sDAC_mem_24Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_7_cascade_\ : std_logic;
signal \sDAC_data_2_39_ns_1_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_7\ : std_logic;
signal \sDAC_mem_28Z0Z_3\ : std_logic;
signal \sDAC_mem_26Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_32Z0Z_7\ : std_logic;
signal \sDAC_mem_31Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_5_cascade_\ : std_logic;
signal \sDAC_data_2_39_ns_1_5_cascade_\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_5\ : std_logic;
signal \sDAC_mem_26Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_32Z0Z_5\ : std_logic;
signal \sDAC_mem_29Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_5\ : std_logic;
signal \sDAC_mem_31Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_5\ : std_logic;
signal \sDAC_mem_24Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_6\ : std_logic;
signal \sDAC_data_2_39_ns_1_6\ : std_logic;
signal \sDAC_mem_29Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_7\ : std_logic;
signal \sDAC_mem_26Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_32Z0Z_6\ : std_logic;
signal \sDAC_mem_24Z0Z_0\ : std_logic;
signal \sDAC_mem_17Z0Z_3\ : std_logic;
signal \spi_slave_inst.spi_miso\ : std_logic;
signal spi_select_c : std_logic;
signal spi_miso_ft_c : std_logic;
signal \sDAC_mem_36Z0Z_2\ : std_logic;
signal \sDAC_mem_36Z0Z_3\ : std_logic;
signal \sDAC_mem_36Z0Z_4\ : std_logic;
signal \sDAC_mem_37Z0Z_2\ : std_logic;
signal \sDAC_mem_37Z0Z_3\ : std_logic;
signal \sDAC_mem_37Z0Z_4\ : std_logic;
signal \sDAC_mem_8Z0Z_2\ : std_logic;
signal \sDAC_mem_8Z0Z_4\ : std_logic;
signal \sDAC_mem_8Z0Z_6\ : std_logic;
signal \sDAC_mem_8Z0Z_7\ : std_logic;
signal \sDAC_mem_8_1_sqmuxa\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_7\ : std_logic;
signal \sDAC_mem_20Z0Z_4\ : std_logic;
signal \sDAC_mem_20Z0Z_5\ : std_logic;
signal \sDAC_mem_20Z0Z_6\ : std_logic;
signal \sDAC_mem_23Z0Z_7\ : std_logic;
signal \sDAC_mem_22Z0Z_7\ : std_logic;
signal \sDAC_mem_23Z0Z_0\ : std_logic;
signal \sDAC_mem_22Z0Z_0\ : std_logic;
signal \sDAC_data_2_13_bm_1_7_cascade_\ : std_logic;
signal \sDAC_mem_7Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_7\ : std_logic;
signal \sDAC_data_2_32_ns_1_7\ : std_logic;
signal \sDAC_mem_34Z0Z_4\ : std_logic;
signal \sDAC_mem_2Z0Z_4\ : std_logic;
signal \sDAC_mem_3Z0Z_4\ : std_logic;
signal \sDAC_data_2_6_bm_1_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_7\ : std_logic;
signal \sDAC_mem_36Z0Z_5\ : std_logic;
signal \sDAC_mem_37Z0Z_5\ : std_logic;
signal \sDAC_data_2_13_am_1_8_cascade_\ : std_logic;
signal \sDAC_mem_5Z0Z_5\ : std_logic;
signal \sDAC_mem_4Z0Z_5\ : std_logic;
signal \sDAC_mem_36Z0Z_6\ : std_logic;
signal \sDAC_mem_37Z0Z_6\ : std_logic;
signal \sDAC_data_2_13_am_1_9_cascade_\ : std_logic;
signal \sDAC_mem_5Z0Z_6\ : std_logic;
signal \sDAC_mem_4Z0Z_6\ : std_logic;
signal \sDAC_mem_6Z0Z_7\ : std_logic;
signal \sDAC_data_2_13_bm_1_10_cascade_\ : std_logic;
signal \sDAC_mem_7Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_9\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_9\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_9_cascade_\ : std_logic;
signal \sDAC_data_2_9_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_9\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_9\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_9\ : std_logic;
signal \sDAC_data_2_14_ns_1_9\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_9\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_9\ : std_logic;
signal \sDAC_data_2_32_ns_1_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_9\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_9_cascade_\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_9\ : std_logic;
signal \sDAC_data_2_41_ns_1_9\ : std_logic;
signal \sDAC_mem_2Z0Z_5\ : std_logic;
signal \sDAC_mem_34Z0Z_5\ : std_logic;
signal \sDAC_data_2_6_bm_1_8_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_5\ : std_logic;
signal \sDAC_mem_33Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_10_cascade_\ : std_logic;
signal \sDAC_mem_1Z0Z_7\ : std_logic;
signal \sDAC_mem_32Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_27Z0Z_10\ : std_logic;
signal \sDAC_mem_1Z0Z_0\ : std_logic;
signal \sDAC_mem_32Z0Z_0\ : std_logic;
signal \sDAC_mem_33Z0Z_0\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_27Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_10\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_10\ : std_logic;
signal \sDAC_data_2_32_ns_1_10\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_10\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_10\ : std_logic;
signal \sDAC_data_2_14_ns_1_10_cascade_\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_10\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_10\ : std_logic;
signal \sDAC_data_2_41_ns_1_10_cascade_\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_10\ : std_logic;
signal \sDAC_data_2_10_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_10\ : std_logic;
signal \sDAC_mem_36Z0Z_7\ : std_logic;
signal \sDAC_mem_37Z0Z_7\ : std_logic;
signal \sDAC_data_2_13_am_1_10_cascade_\ : std_logic;
signal \sDAC_mem_5Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_10\ : std_logic;
signal \sDAC_mem_4Z0Z_7\ : std_logic;
signal \sDAC_mem_36Z0Z_0\ : std_logic;
signal \sDAC_mem_37Z0Z_0\ : std_logic;
signal \sDAC_data_2_13_am_1_3_cascade_\ : std_logic;
signal \sDAC_mem_5Z0Z_0\ : std_logic;
signal \sDAC_mem_4Z0Z_0\ : std_logic;
signal \sDAC_mem_4_1_sqmuxa\ : std_logic;
signal \sDAC_mem_36Z0Z_1\ : std_logic;
signal \sDAC_mem_4Z0Z_1\ : std_logic;
signal \sDAC_mem_37Z0Z_1\ : std_logic;
signal \sDAC_data_2_13_am_1_4_cascade_\ : std_logic;
signal \sDAC_mem_5Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_10\ : std_logic;
signal \sDAC_mem_26_1_sqmuxa\ : std_logic;
signal \N_142_cascade_\ : std_logic;
signal \sDAC_mem_30Z0Z_2\ : std_logic;
signal \sDAC_mem_30Z0Z_3\ : std_logic;
signal \sDAC_mem_30Z0Z_5\ : std_logic;
signal \sDAC_mem_30Z0Z_6\ : std_logic;
signal \sDAC_mem_30_1_sqmuxa\ : std_logic;
signal \sDAC_mem_23Z0Z_5\ : std_logic;
signal \sDAC_mem_22Z0Z_5\ : std_logic;
signal \sDAC_mem_23Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_9\ : std_logic;
signal \sDAC_mem_22Z0Z_6\ : std_logic;
signal \sDAC_mem_22_1_sqmuxa\ : std_logic;
signal \sDAC_mem_29Z0Z_1\ : std_logic;
signal \sDAC_mem_30Z0Z_1\ : std_logic;
signal \sDAC_mem_31Z0Z_1\ : std_logic;
signal \sDAC_mem_31Z0Z_4\ : std_logic;
signal \sDAC_mem_30Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_10_cascade_\ : std_logic;
signal \sDAC_data_2_39_ns_1_10_cascade_\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_10\ : std_logic;
signal \sDAC_mem_26Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_32Z0Z_10\ : std_logic;
signal \sDAC_mem_29Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_10\ : std_logic;
signal \sDAC_mem_31Z0Z_7\ : std_logic;
signal \sDAC_mem_30Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_10\ : std_logic;
signal \sDAC_mem_24Z0Z_7\ : std_logic;
signal \sDAC_mem_24_1_sqmuxa\ : std_logic;
signal \sDAC_data_RNO_32Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_3\ : std_logic;
signal \sDAC_mem_25Z0Z_4\ : std_logic;
signal \sDAC_mem_25Z0Z_7\ : std_logic;
signal \sDAC_mem_25Z0Z_2\ : std_logic;
signal \sDAC_mem_25Z0Z_5\ : std_logic;
signal \sDAC_mem_25Z0Z_0\ : std_logic;
signal \sDAC_mem_25Z0Z_6\ : std_logic;
signal \sDAC_mem_25Z0Z_3\ : std_logic;
signal \sDAC_mem_34_1_sqmuxa\ : std_logic;
signal \sDAC_mem_39Z0Z_0\ : std_logic;
signal \sDAC_mem_39Z0Z_1\ : std_logic;
signal \sDAC_mem_39Z0Z_2\ : std_logic;
signal \sDAC_mem_39Z0Z_4\ : std_logic;
signal \sDAC_mem_39Z0Z_7\ : std_logic;
signal \sDAC_mem_37_1_sqmuxa\ : std_logic;
signal \sDAC_mem_39_1_sqmuxa\ : std_logic;
signal \sDAC_mem_36_1_sqmuxa\ : std_logic;
signal \N_288\ : std_logic;
signal \sAddressZ0Z_3\ : std_logic;
signal \N_288_cascade_\ : std_logic;
signal \sAddressZ0Z_0\ : std_logic;
signal \sDAC_mem_35Z0Z_0\ : std_logic;
signal \sDAC_mem_35Z0Z_2\ : std_logic;
signal \sDAC_mem_35Z0Z_4\ : std_logic;
signal \sDAC_mem_35Z0Z_5\ : std_logic;
signal \sDAC_mem_35Z0Z_6\ : std_logic;
signal \sDAC_mem_35_1_sqmuxa\ : std_logic;
signal \sDAC_mem_21Z0Z_4\ : std_logic;
signal \sDAC_mem_21Z0Z_5\ : std_logic;
signal \sDAC_mem_21Z0Z_6\ : std_logic;
signal \sDAC_mem_21Z0Z_7\ : std_logic;
signal \sDAC_mem_21_1_sqmuxa\ : std_logic;
signal \sDAC_mem_7Z0Z_3\ : std_logic;
signal \sDAC_data_2_13_bm_1_6_cascade_\ : std_logic;
signal \sDAC_mem_39Z0Z_3\ : std_logic;
signal \sDAC_mem_6Z0Z_3\ : std_logic;
signal \sDAC_mem_6Z0Z_4\ : std_logic;
signal \sDAC_mem_6Z0Z_5\ : std_logic;
signal \sDAC_mem_7Z0Z_5\ : std_logic;
signal \sDAC_data_2_13_bm_1_8_cascade_\ : std_logic;
signal \sDAC_mem_39Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_8\ : std_logic;
signal \sDAC_data_2_32_ns_1_8\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_8\ : std_logic;
signal \sDAC_data_2_14_ns_1_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_8\ : std_logic;
signal \sDAC_data_2_41_ns_1_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_8\ : std_logic;
signal \sDAC_data_2_8_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_8\ : std_logic;
signal \sDAC_mem_2Z0Z_1\ : std_logic;
signal \sDAC_mem_34Z0Z_1\ : std_logic;
signal \sDAC_mem_35Z0Z_1\ : std_logic;
signal \sDAC_data_2_6_bm_1_4_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_6_cascade_\ : std_logic;
signal \sDAC_mem_8Z0Z_3\ : std_logic;
signal \sDAC_data_2_20_am_1_6_cascade_\ : std_logic;
signal \sDAC_data_2_24_ns_1_6\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_4\ : std_logic;
signal \sDAC_data_2_32_ns_1_4\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_4\ : std_logic;
signal \sDAC_data_2_14_ns_1_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_2_41_ns_1_4\ : std_logic;
signal \sDAC_data_2_4_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_4\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_3\ : std_logic;
signal \sDAC_data_2_32_ns_1_3\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_3\ : std_logic;
signal \sDAC_data_2_14_ns_1_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \sDAC_data_2_41_ns_1_3\ : std_logic;
signal \sDAC_data_2_3_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_3\ : std_logic;
signal \sDAC_mem_16Z0Z_7\ : std_logic;
signal \sDAC_mem_17Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_10\ : std_logic;
signal \sDAC_mem_19Z0Z_3\ : std_logic;
signal \sDAC_mem_18Z0Z_3\ : std_logic;
signal \sDAC_mem_23Z0Z_1\ : std_logic;
signal \sDAC_mem_22Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_4\ : std_logic;
signal \sDAC_mem_27Z0Z_2\ : std_logic;
signal \sDAC_mem_27Z0Z_3\ : std_logic;
signal \sDAC_mem_27Z0Z_4\ : std_logic;
signal \sDAC_mem_27Z0Z_5\ : std_logic;
signal \sDAC_mem_27Z0Z_6\ : std_logic;
signal \sDAC_mem_27Z0Z_7\ : std_logic;
signal \sEEADC_freqZ0Z_0\ : std_logic;
signal \sEEADC_freqZ0Z_6\ : std_logic;
signal \sEEADC_freqZ0Z_7\ : std_logic;
signal \sDAC_mem_31Z0Z_0\ : std_logic;
signal \sDAC_mem_30Z0Z_0\ : std_logic;
signal \sDAC_mem_29Z0Z_0\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_3_cascade_\ : std_logic;
signal \sDAC_data_2_39_ns_1_3\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_3\ : std_logic;
signal \sDAC_mem_28Z0Z_0\ : std_logic;
signal \sDAC_mem_24Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_31Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_24Z0Z_4\ : std_logic;
signal \sDAC_data_2_39_ns_1_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_23Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_4\ : std_logic;
signal \sDAC_mem_26Z0Z_1\ : std_logic;
signal \sDAC_mem_27Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_32Z0Z_4\ : std_logic;
signal \sDAC_mem_28Z0Z_1\ : std_logic;
signal \sDAC_mem_28Z0Z_2\ : std_logic;
signal \sDAC_mem_28Z0Z_4\ : std_logic;
signal \sDAC_mem_28Z0Z_5\ : std_logic;
signal \sDAC_mem_28Z0Z_7\ : std_logic;
signal \sDAC_mem_28_1_sqmuxa\ : std_logic;
signal \sDAC_mem_25Z0Z_1\ : std_logic;
signal \sDAC_mem_25_1_sqmuxa\ : std_logic;
signal \sDAC_mem_17Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_4\ : std_logic;
signal \sDAC_mem_38Z0Z_0\ : std_logic;
signal \sDAC_mem_38Z0Z_2\ : std_logic;
signal \sDAC_mem_38Z0Z_3\ : std_logic;
signal \sDAC_mem_38Z0Z_4\ : std_logic;
signal \sDAC_mem_38Z0Z_5\ : std_logic;
signal \sDAC_mem_38Z0Z_7\ : std_logic;
signal \sDAC_mem_38_1_sqmuxa\ : std_logic;
signal \sDAC_mem_40Z0Z_2\ : std_logic;
signal \sDAC_mem_40Z0Z_3\ : std_logic;
signal \sDAC_mem_40Z0Z_4\ : std_logic;
signal \sDAC_mem_40Z0Z_6\ : std_logic;
signal \sDAC_mem_40Z0Z_7\ : std_logic;
signal \sDAC_mem_40_1_sqmuxa\ : std_logic;
signal \sDAC_mem_21Z0Z_0\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_3\ : std_logic;
signal \sDAC_mem_20Z0Z_0\ : std_logic;
signal \sDAC_mem_21Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_4\ : std_logic;
signal \sDAC_mem_20Z0Z_1\ : std_logic;
signal \sDAC_mem_21Z0Z_2\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_5\ : std_logic;
signal \sDAC_mem_20Z0Z_2\ : std_logic;
signal \sDAC_mem_21Z0Z_3\ : std_logic;
signal \sDAC_mem_20Z0Z_3\ : std_logic;
signal \sDAC_mem_33Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_6_cascade_\ : std_logic;
signal \sDAC_mem_32Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_27Z0Z_6\ : std_logic;
signal \sDAC_mem_1Z0Z_3\ : std_logic;
signal \sDAC_mem_33Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_26Z0Z_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_7\ : std_logic;
signal \sDAC_mem_32Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_27Z0Z_7\ : std_logic;
signal \sDAC_mem_1Z0Z_4\ : std_logic;
signal \sDAC_mem_1_1_sqmuxa\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_4Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_14Z0Z_6\ : std_logic;
signal \sDAC_data_2_14_ns_1_6\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_30Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_21Z0Z_6\ : std_logic;
signal \sDAC_data_2_32_ns_1_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_20Z0Z_6\ : std_logic;
signal \sDAC_mem_pointerZ0Z_3\ : std_logic;
signal \sDAC_data_RNO_10Z0Z_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_11Z0Z_6\ : std_logic;
signal \sDAC_mem_pointerZ0Z_4\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_6\ : std_logic;
signal \sDAC_data_2_41_ns_1_6_cascade_\ : std_logic;
signal \sDAC_data_RNO_1Z0Z_6\ : std_logic;
signal \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\ : std_logic;
signal \sDAC_data_2_6_cascade_\ : std_logic;
signal \sDAC_dataZ0Z_6\ : std_logic;
signal op_eq_scounterdac10_g : std_logic;
signal \sDAC_mem_2Z0Z_3\ : std_logic;
signal \sDAC_mem_34Z0Z_3\ : std_logic;
signal \sDAC_mem_35Z0Z_3\ : std_logic;
signal \sDAC_data_2_6_bm_1_6_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_8_cascade_\ : std_logic;
signal \sDAC_mem_40Z0Z_5\ : std_logic;
signal \sDAC_mem_8Z0Z_5\ : std_logic;
signal \sDAC_data_2_20_am_1_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_8_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_8\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_8\ : std_logic;
signal \sDAC_mem_38Z0Z_6\ : std_logic;
signal \sDAC_mem_39Z0Z_6\ : std_logic;
signal \sDAC_data_2_13_bm_1_9_cascade_\ : std_logic;
signal \sDAC_mem_7Z0Z_6\ : std_logic;
signal \sDAC_data_RNO_5Z0Z_9\ : std_logic;
signal \sDAC_mem_6Z0Z_6\ : std_logic;
signal \sDAC_mem_6_1_sqmuxa\ : std_logic;
signal \sDAC_mem_40Z0Z_0\ : std_logic;
signal \sDAC_mem_8Z0Z_0\ : std_logic;
signal \sDAC_data_2_20_am_1_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_3\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_3\ : std_logic;
signal \sDAC_mem_3_1_sqmuxa\ : std_logic;
signal \sDAC_mem_34Z0Z_7\ : std_logic;
signal \sDAC_mem_2Z0Z_7\ : std_logic;
signal \sDAC_mem_35Z0Z_7\ : std_logic;
signal \sDAC_data_2_6_bm_1_10_cascade_\ : std_logic;
signal \sDAC_mem_3Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_15Z0Z_10\ : std_logic;
signal \sDAC_mem_40Z0Z_1\ : std_logic;
signal \sDAC_mem_8Z0Z_1\ : std_logic;
signal \sDAC_data_2_20_am_1_4_cascade_\ : std_logic;
signal \sDAC_mem_pointerZ0Z_5\ : std_logic;
signal \sDAC_data_RNO_17Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_8Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_RNO_7Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_2Z0Z_4\ : std_logic;
signal \N_284_cascade_\ : std_logic;
signal \N_284\ : std_logic;
signal \N_280\ : std_logic;
signal \sPointerZ0Z_1\ : std_logic;
signal un1_spointer11_0 : std_logic;
signal \sDAC_mem_14Z0Z_2\ : std_logic;
signal \sDAC_mem_14Z0Z_3\ : std_logic;
signal \sDAC_mem_14Z0Z_6\ : std_logic;
signal \sDAC_mem_14_1_sqmuxa\ : std_logic;
signal \sDAC_mem_14Z0Z_4\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_7_cascade_\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_7\ : std_logic;
signal \sDAC_data_2_24_ns_1_7\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_8_cascade_\ : std_logic;
signal \sDAC_data_2_24_ns_1_8\ : std_logic;
signal \sDAC_mem_12Z0Z_4\ : std_logic;
signal \sDAC_mem_14Z0Z_5\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_8\ : std_logic;
signal \sDAC_mem_12Z0Z_5\ : std_logic;
signal \sEEADC_freqZ0Z_1\ : std_logic;
signal \sEEADC_freq_1_sqmuxa\ : std_logic;
signal \sDAC_mem_17Z0Z_0\ : std_logic;
signal \sDAC_mem_16Z0Z_0\ : std_logic;
signal \sDAC_data_RNO_29Z0Z_3\ : std_logic;
signal \sDAC_mem_16Z0Z_3\ : std_logic;
signal \sDAC_mem_20Z0Z_7\ : std_logic;
signal \sDAC_mem_20_1_sqmuxa\ : std_logic;
signal \sDAC_mem_41Z0Z_0\ : std_logic;
signal \sDAC_mem_41Z0Z_1\ : std_logic;
signal \sDAC_mem_41Z0Z_2\ : std_logic;
signal \sDAC_mem_41Z0Z_3\ : std_logic;
signal \sDAC_mem_41Z0Z_4\ : std_logic;
signal \sDAC_mem_41Z0Z_5\ : std_logic;
signal \sDAC_mem_41Z0Z_6\ : std_logic;
signal \sDAC_mem_41Z0Z_7\ : std_logic;
signal \sDAC_mem_42Z0Z_0\ : std_logic;
signal \sDAC_mem_42Z0Z_1\ : std_logic;
signal \sDAC_mem_42Z0Z_2\ : std_logic;
signal \sDAC_mem_42Z0Z_3\ : std_logic;
signal \sDAC_mem_42Z0Z_4\ : std_logic;
signal \sDAC_mem_42Z0Z_5\ : std_logic;
signal \sDAC_mem_42Z0Z_6\ : std_logic;
signal \sDAC_mem_42Z0Z_7\ : std_logic;
signal \sDAC_mem_10Z0Z_0\ : std_logic;
signal \sDAC_mem_10Z0Z_1\ : std_logic;
signal \sDAC_mem_10Z0Z_2\ : std_logic;
signal \sDAC_mem_10Z0Z_3\ : std_logic;
signal \sDAC_mem_10Z0Z_4\ : std_logic;
signal \sDAC_mem_10Z0Z_5\ : std_logic;
signal \sDAC_mem_10Z0Z_6\ : std_logic;
signal \sDAC_mem_10_1_sqmuxa\ : std_logic;
signal \sDAC_mem_42_1_sqmuxa\ : std_logic;
signal \sAddressZ0Z_2\ : std_logic;
signal \sAddressZ0Z_1\ : std_logic;
signal \sDAC_mem_30_1_sqmuxa_0_a2_1_0\ : std_logic;
signal \N_275\ : std_logic;
signal \sAddressZ0Z_4\ : std_logic;
signal \N_286\ : std_logic;
signal \N_278_cascade_\ : std_logic;
signal \N_142\ : std_logic;
signal \sDAC_mem_15Z0Z_2\ : std_logic;
signal \sDAC_mem_15Z0Z_3\ : std_logic;
signal \sDAC_mem_15Z0Z_4\ : std_logic;
signal \sDAC_mem_15Z0Z_5\ : std_logic;
signal \sDAC_mem_15Z0Z_6\ : std_logic;
signal \sDAC_mem_15_1_sqmuxa\ : std_logic;
signal \sDAC_mem_11Z0Z_0\ : std_logic;
signal \sDAC_mem_11Z0Z_1\ : std_logic;
signal \sDAC_mem_11Z0Z_2\ : std_logic;
signal \sDAC_mem_11Z0Z_3\ : std_logic;
signal \sDAC_mem_11Z0Z_4\ : std_logic;
signal \sDAC_mem_11Z0Z_5\ : std_logic;
signal \sDAC_mem_11Z0Z_6\ : std_logic;
signal \sDAC_mem_11Z0Z_7\ : std_logic;
signal \sDAC_mem_11_1_sqmuxa\ : std_logic;
signal \sDAC_mem_15Z0Z_0\ : std_logic;
signal \sDAC_mem_14Z0Z_0\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_3_cascade_\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_3\ : std_logic;
signal \sDAC_data_2_24_ns_1_3\ : std_logic;
signal \sDAC_mem_pointerZ0Z_2\ : std_logic;
signal \sDAC_mem_pointerZ0Z_1\ : std_logic;
signal \sDAC_data_RNO_18Z0Z_4_cascade_\ : std_logic;
signal \sDAC_data_2_24_ns_1_4\ : std_logic;
signal \sDAC_mem_12Z0Z_0\ : std_logic;
signal \sDAC_mem_15Z0Z_1\ : std_logic;
signal \sDAC_mem_14Z0Z_1\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_4\ : std_logic;
signal \sDAC_mem_12Z0Z_1\ : std_logic;
signal \sDAC_mem_27Z0Z_0\ : std_logic;
signal \sDAC_mem_27_1_sqmuxa\ : std_logic;
signal \sDAC_mem_13Z0Z_6\ : std_logic;
signal \sDAC_mem_13Z0Z_5\ : std_logic;
signal \sDAC_mem_16Z0Z_1\ : std_logic;
signal \sDAC_mem_16_1_sqmuxa\ : std_logic;
signal \sEEDACZ0Z_7\ : std_logic;
signal \sAddressZ0Z_5\ : std_logic;
signal \N_139\ : std_logic;
signal \N_278\ : std_logic;
signal \sDAC_mem_41_1_sqmuxa\ : std_logic;
signal \N_285\ : std_logic;
signal \N_1480\ : std_logic;
signal \N_360\ : std_logic;
signal \sEEDACZ0Z_0\ : std_logic;
signal \sEEDACZ0Z_1\ : std_logic;
signal \sEEDACZ0Z_2\ : std_logic;
signal \sEEDACZ0Z_3\ : std_logic;
signal \sEEDACZ0Z_4\ : std_logic;
signal \sEEDACZ0Z_5\ : std_logic;
signal \sEEDACZ0Z_6\ : std_logic;
signal \sEEDAC_1_sqmuxa\ : std_logic;
signal \sDAC_mem_9Z0Z_0\ : std_logic;
signal \sDAC_mem_9Z0Z_1\ : std_logic;
signal \sDAC_mem_9Z0Z_2\ : std_logic;
signal \sDAC_mem_9Z0Z_3\ : std_logic;
signal \sDAC_mem_9Z0Z_4\ : std_logic;
signal spi_data_mosi_5 : std_logic;
signal \sDAC_mem_9Z0Z_5\ : std_logic;
signal \sDAC_mem_9Z0Z_6\ : std_logic;
signal \sDAC_mem_9Z0Z_7\ : std_logic;
signal \sDAC_mem_9_1_sqmuxa\ : std_logic;
signal \N_14_3_cascade_\ : std_logic;
signal \N_8_cascade_\ : std_logic;
signal \sDAC_spi_startZ0\ : std_logic;
signal un1_scounterdac8_i_a2_1_2 : std_logic;
signal un1_scounterdac8_i_a2_0 : std_logic;
signal \sDAC_data_RNO_18Z0Z_10\ : std_logic;
signal \sDAC_mem_pointerZ0Z_0\ : std_logic;
signal \sDAC_mem_15Z0Z_7\ : std_logic;
signal \sDAC_mem_14Z0Z_7\ : std_logic;
signal \sDAC_data_RNO_19Z0Z_10\ : std_logic;
signal spi_data_mosi_0 : std_logic;
signal \sDAC_mem_13Z0Z_0\ : std_logic;
signal spi_data_mosi_1 : std_logic;
signal \sDAC_mem_13Z0Z_1\ : std_logic;
signal spi_data_mosi_2 : std_logic;
signal \sDAC_mem_13Z0Z_2\ : std_logic;
signal spi_data_mosi_3 : std_logic;
signal \sDAC_mem_13Z0Z_3\ : std_logic;
signal spi_data_mosi_4 : std_logic;
signal \sDAC_mem_13Z0Z_4\ : std_logic;
signal \sDAC_mem_13Z0Z_7\ : std_logic;
signal \sDAC_mem_13_1_sqmuxa\ : std_logic;
signal spi_data_mosi_7 : std_logic;
signal \sDAC_mem_12Z0Z_7\ : std_logic;
signal spi_data_mosi_6 : std_logic;
signal \sDAC_mem_12Z0Z_6\ : std_logic;
signal pll_clk128_g : std_logic;
signal \sDAC_mem_12_1_sqmuxa\ : std_logic;
signal \N_14_3\ : std_logic;
signal \bfn_22_10_0_\ : std_logic;
signal un2_scounterdac_cry_1 : std_logic;
signal \sCounterDACZ0Z_3\ : std_logic;
signal un2_scounterdac_cry_2 : std_logic;
signal un2_scounterdac_cry_3 : std_logic;
signal \sCounterDACZ0Z_5\ : std_logic;
signal un2_scounterdac_cry_4 : std_logic;
signal \un2_scounterdac_cry_5_THRU_CO\ : std_logic;
signal un2_scounterdac_cry_5 : std_logic;
signal un2_scounterdac_cry_6 : std_logic;
signal \sCounterDACZ0Z_8\ : std_logic;
signal \un2_scounterdac_cry_7_THRU_CO\ : std_logic;
signal un2_scounterdac_cry_7 : std_logic;
signal un2_scounterdac_cry_8 : std_logic;
signal \bfn_22_11_0_\ : std_logic;
signal pll_clk64_0_g : std_logic;
signal \LED3_c_i_g\ : std_logic;
signal spi_mosi_rpi_c : std_logic;
signal spi_mosi_flash_c : std_logic;
signal \sCounterDACZ0Z_4\ : std_logic;
signal \sCounterDACZ0Z_1\ : std_logic;
signal \sCounterDACZ0Z_7\ : std_logic;
signal \sCounterDACZ0Z_2\ : std_logic;
signal \sCounterDACZ0Z_9\ : std_logic;
signal \sCounterDACZ0Z_6\ : std_logic;
signal spi_cs_rpi_c : std_logic;
signal spi_cs_flash_c : std_logic;
signal spi_sclk_rpi_c : std_logic;
signal cs_rpi2flash_c : std_logic;
signal spi_sclk_flash_c : std_logic;
signal op_eq_scounterdac10_0_a2_0 : std_logic;
signal \N_23\ : std_logic;
signal \sCounterDACZ0Z_0\ : std_logic;
signal \N_22\ : std_logic;
signal op_eq_scounterdac10 : std_logic;
signal \_gnd_net_\ : std_logic;

signal \RAM_ADD_wire\ : std_logic_vector(18 downto 0);
signal spi_mosi_rpi_wire : std_logic;
signal spi_sclk_rpi_wire : std_logic;
signal spi_miso_ft_wire : std_logic;
signal \ADC5_wire\ : std_logic;
signal \LED_ACQ_wire\ : std_logic;
signal reset_rpi_wire : std_logic;
signal trig_rpi_wire : std_logic;
signal \ADC2_wire\ : std_logic;
signal \DAC_mosi_wire\ : std_logic;
signal \RAM_nWE_wire\ : std_logic;
signal \ADC0_wire\ : std_logic;
signal \RAM_nLB_wire\ : std_logic;
signal spi_select_wire : std_logic;
signal \RAM_nCE_wire\ : std_logic;
signal spi_sclk_flash_wire : std_logic;
signal \ADC3_wire\ : std_logic;
signal pon_wire : std_logic;
signal \DAC_sclk_wire\ : std_logic;
signal \ADC1_wire\ : std_logic;
signal spi_cs_flash_wire : std_logic;
signal spi_miso_flash_wire : std_logic;
signal trig_ext_wire : std_logic;
signal top_tour1_wire : std_logic;
signal \LED_MODE_wire\ : std_logic;
signal \RAM_nUB_wire\ : std_logic;
signal \DAC_cs_wire\ : std_logic;
signal \ADC8_wire\ : std_logic;
signal \ADC_clk_wire\ : std_logic;
signal poff_wire : std_logic;
signal \ADC4_wire\ : std_logic;
signal \ADC6_wire\ : std_logic;
signal \ADC7_wire\ : std_logic;
signal button_mode_wire : std_logic;
signal spi_sclk_ft_wire : std_logic;
signal trig_ft_wire : std_logic;
signal \ADC9_wire\ : std_logic;
signal cs_rpi2flash_wire : std_logic;
signal \LED3_wire\ : std_logic;
signal spi_mosi_ft_wire : std_logic;
signal \RAM_nOE_wire\ : std_logic;
signal clk_wire : std_logic;
signal top_tour2_wire : std_logic;
signal spi_cs_rpi_wire : std_logic;
signal spi_miso_rpi_wire : std_logic;
signal spi_cs_ft_wire : std_logic;
signal spi_mosi_flash_wire : std_logic;
signal \pll128M2_inst.pll128M2_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    RAM_ADD <= \RAM_ADD_wire\;
    spi_mosi_rpi_wire <= spi_mosi_rpi;
    spi_sclk_rpi_wire <= spi_sclk_rpi;
    spi_miso_ft <= spi_miso_ft_wire;
    \ADC5_wire\ <= ADC5;
    LED_ACQ <= \LED_ACQ_wire\;
    reset_rpi_wire <= reset_rpi;
    trig_rpi_wire <= trig_rpi;
    \ADC2_wire\ <= ADC2;
    DAC_mosi <= \DAC_mosi_wire\;
    RAM_nWE <= \RAM_nWE_wire\;
    \ADC0_wire\ <= ADC0;
    RAM_nLB <= \RAM_nLB_wire\;
    spi_select_wire <= spi_select;
    RAM_nCE <= \RAM_nCE_wire\;
    spi_sclk_flash <= spi_sclk_flash_wire;
    \ADC3_wire\ <= ADC3;
    pon <= pon_wire;
    DAC_sclk <= \DAC_sclk_wire\;
    \ADC1_wire\ <= ADC1;
    spi_cs_flash <= spi_cs_flash_wire;
    spi_miso_flash_wire <= spi_miso_flash;
    trig_ext_wire <= trig_ext;
    top_tour1_wire <= top_tour1;
    LED_MODE <= \LED_MODE_wire\;
    RAM_nUB <= \RAM_nUB_wire\;
    DAC_cs <= \DAC_cs_wire\;
    \ADC8_wire\ <= ADC8;
    ADC_clk <= \ADC_clk_wire\;
    poff <= poff_wire;
    \ADC4_wire\ <= ADC4;
    \ADC6_wire\ <= ADC6;
    \ADC7_wire\ <= ADC7;
    button_mode_wire <= button_mode;
    spi_sclk_ft_wire <= spi_sclk_ft;
    trig_ft_wire <= trig_ft;
    \ADC9_wire\ <= ADC9;
    cs_rpi2flash_wire <= cs_rpi2flash;
    LED3 <= \LED3_wire\;
    spi_mosi_ft_wire <= spi_mosi_ft;
    RAM_nOE <= \RAM_nOE_wire\;
    clk_wire <= clk;
    top_tour2_wire <= top_tour2;
    spi_cs_rpi_wire <= spi_cs_rpi;
    spi_miso_rpi <= spi_miso_rpi_wire;
    spi_cs_ft_wire <= spi_cs_ft;
    spi_mosi_flash <= spi_mosi_flash_wire;
    \pll128M2_inst.pll128M2_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll128M2_inst.pll128M2_inst\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1010100",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \pll128M2_inst.pll_clk64_0\,
            REFERENCECLK => \N__20538\,
            RESETB => \N__32326\,
            BYPASS => \GNDG0\,
            PLLOUTCOREA => \pll128M2_inst.pll_clk128\,
            SDI => \GNDG0\,
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll128M2_inst.pll128M2_inst_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => \GNDG0\,
            PLLOUTGLOBALA => OPEN,
            SCLK => \GNDG0\
        );

    \RAM_ADD_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54196\,
            DIN => \N__54195\,
            DOUT => \N__54194\,
            PACKAGEPIN => \RAM_ADD_wire\(5)
        );

    \RAM_ADD_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54196\,
            PADOUT => \N__54195\,
            PADIN => \N__54194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28581\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_mosi_rpi_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54187\,
            DIN => \N__54186\,
            DOUT => \N__54185\,
            PACKAGEPIN => spi_mosi_rpi_wire
        );

    \spi_mosi_rpi_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54187\,
            PADOUT => \N__54186\,
            PADIN => \N__54185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_mosi_rpi_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_sclk_rpi_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54178\,
            DIN => \N__54177\,
            DOUT => \N__54176\,
            PACKAGEPIN => spi_sclk_rpi_wire
        );

    \spi_sclk_rpi_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54178\,
            PADOUT => \N__54177\,
            PADIN => \N__54176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_sclk_rpi_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_miso_ft_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54169\,
            DIN => \N__54168\,
            DOUT => \N__54167\,
            PACKAGEPIN => spi_miso_ft_wire
        );

    \spi_miso_ft_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54169\,
            PADOUT => \N__54168\,
            PADIN => \N__54167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__38490\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC5_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54160\,
            DIN => \N__54159\,
            DOUT => \N__54158\,
            PACKAGEPIN => \ADC5_wire\
        );

    \ADC5_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54160\,
            PADOUT => \N__54159\,
            PADIN => \N__54158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC5_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_ACQ_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54151\,
            DIN => \N__54150\,
            DOUT => \N__54149\,
            PACKAGEPIN => \LED_ACQ_wire\
        );

    \LED_ACQ_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54151\,
            PADOUT => \N__54150\,
            PADIN => \N__54149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22260\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \reset_rpi_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54142\,
            DIN => \N__54141\,
            DOUT => \N__54140\,
            PACKAGEPIN => reset_rpi_wire
        );

    \reset_rpi_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54142\,
            PADOUT => \N__54141\,
            PADIN => \N__54140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \LED3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54133\,
            DIN => \N__54132\,
            DOUT => \N__54131\,
            PACKAGEPIN => RAM_DATA(6)
        );

    \RAM_DATA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__54133\,
            PADOUT => \N__54132\,
            PADIN => \N__54131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__30558\,
            DIN0 => \RAM_DATA_in_6\,
            DOUT0 => \N__31539\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54124\,
            DIN => \N__54123\,
            DOUT => \N__54122\,
            PACKAGEPIN => \RAM_ADD_wire\(9)
        );

    \RAM_ADD_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54124\,
            PADOUT => \N__54123\,
            PADIN => \N__54122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28392\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54115\,
            DIN => \N__54114\,
            DOUT => \N__54113\,
            PACKAGEPIN => RAM_DATA(11)
        );

    \RAM_DATA_iobuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__54115\,
            PADOUT => \N__54114\,
            PADIN => \N__54113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__31773\,
            DIN0 => \RAM_DATA_in_11\,
            DOUT0 => \N__31455\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \trig_rpi_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54106\,
            DIN => \N__54105\,
            DOUT => \N__54104\,
            PACKAGEPIN => trig_rpi_wire
        );

    \trig_rpi_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54106\,
            PADOUT => \N__54105\,
            PADIN => \N__54104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => trig_rpi_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54097\,
            DIN => \N__54096\,
            DOUT => \N__54095\,
            PACKAGEPIN => RAM_DATA(0)
        );

    \RAM_DATA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__54097\,
            PADOUT => \N__54096\,
            PADIN => \N__54095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__26865\,
            DIN0 => \RAM_DATA_in_0\,
            DOUT0 => \N__30186\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54088\,
            DIN => \N__54087\,
            DOUT => \N__54086\,
            PACKAGEPIN => \ADC2_wire\
        );

    \ADC2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54088\,
            PADOUT => \N__54087\,
            PADIN => \N__54086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC2_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54079\,
            DIN => \N__54078\,
            DOUT => \N__54077\,
            PACKAGEPIN => \RAM_ADD_wire\(18)
        );

    \RAM_ADD_obuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54079\,
            PADOUT => \N__54078\,
            PADIN => \N__54077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28098\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54070\,
            DIN => \N__54069\,
            DOUT => \N__54068\,
            PACKAGEPIN => \RAM_ADD_wire\(2)
        );

    \RAM_ADD_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54070\,
            PADOUT => \N__54069\,
            PADIN => \N__54068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28056\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DAC_mosi_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54061\,
            DIN => \N__54060\,
            DOUT => \N__54059\,
            PACKAGEPIN => \DAC_mosi_wire\
        );

    \DAC_mosi_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54061\,
            PADOUT => \N__54060\,
            PADIN => \N__54059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21147\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54052\,
            DIN => \N__54051\,
            DOUT => \N__54050\,
            PACKAGEPIN => \RAM_ADD_wire\(13)
        );

    \RAM_ADD_obuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54052\,
            PADOUT => \N__54051\,
            PADIN => \N__54050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__30291\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_nWE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54043\,
            DIN => \N__54042\,
            DOUT => \N__54041\,
            PACKAGEPIN => \RAM_nWE_wire\
        );

    \RAM_nWE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54043\,
            PADOUT => \N__54042\,
            PADIN => \N__54041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27660\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54034\,
            DIN => \N__54033\,
            DOUT => \N__54032\,
            PACKAGEPIN => RAM_DATA(7)
        );

    \RAM_DATA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__54034\,
            PADOUT => \N__54033\,
            PADIN => \N__54032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__30486\,
            DIN0 => \RAM_DATA_in_7\,
            DOUT0 => \N__30579\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC0_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54025\,
            DIN => \N__54024\,
            DOUT => \N__54023\,
            PACKAGEPIN => \ADC0_wire\
        );

    \ADC0_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__54025\,
            PADOUT => \N__54024\,
            PADIN => \N__54023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC0_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_nLB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54016\,
            DIN => \N__54015\,
            DOUT => \N__54014\,
            PACKAGEPIN => \RAM_nLB_wire\
        );

    \RAM_nLB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__54016\,
            PADOUT => \N__54015\,
            PADIN => \N__54014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54007\,
            DIN => \N__54006\,
            DOUT => \N__54005\,
            PACKAGEPIN => RAM_DATA(10)
        );

    \RAM_DATA_iobuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__54007\,
            PADOUT => \N__54006\,
            PADIN => \N__54005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__31746\,
            DIN0 => \RAM_DATA_in_10\,
            DOUT0 => \N__31500\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53998\,
            DIN => \N__53997\,
            DOUT => \N__53996\,
            PACKAGEPIN => RAM_DATA(1)
        );

    \RAM_DATA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53998\,
            PADOUT => \N__53997\,
            PADIN => \N__53996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__28326\,
            DIN0 => \RAM_DATA_in_1\,
            DOUT0 => \N__30105\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_select_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53989\,
            DIN => \N__53988\,
            DOUT => \N__53987\,
            PACKAGEPIN => spi_select_wire
        );

    \spi_select_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53989\,
            PADOUT => \N__53988\,
            PADIN => \N__53987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_select_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_nCE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53980\,
            DIN => \N__53979\,
            DOUT => \N__53978\,
            PACKAGEPIN => \RAM_nCE_wire\
        );

    \RAM_nCE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53980\,
            PADOUT => \N__53979\,
            PADIN => \N__53978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_sclk_flash_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53971\,
            DIN => \N__53970\,
            DOUT => \N__53969\,
            PACKAGEPIN => spi_sclk_flash_wire
        );

    \spi_sclk_flash_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53971\,
            PADOUT => \N__53970\,
            PADIN => \N__53969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__52272\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53962\,
            DIN => \N__53961\,
            DOUT => \N__53960\,
            PACKAGEPIN => \RAM_ADD_wire\(3)
        );

    \RAM_ADD_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53962\,
            PADOUT => \N__53961\,
            PADIN => \N__53960\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28662\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53953\,
            DIN => \N__53952\,
            DOUT => \N__53951\,
            PACKAGEPIN => \RAM_ADD_wire\(12)
        );

    \RAM_ADD_obuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53953\,
            PADOUT => \N__53952\,
            PADIN => \N__53951\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__30327\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53944\,
            DIN => \N__53943\,
            DOUT => \N__53942\,
            PACKAGEPIN => \ADC3_wire\
        );

    \ADC3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53944\,
            PADOUT => \N__53943\,
            PADIN => \N__53942\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53935\,
            DIN => \N__53934\,
            DOUT => \N__53933\,
            PACKAGEPIN => RAM_DATA(15)
        );

    \RAM_DATA_iobuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53935\,
            PADOUT => \N__53934\,
            PADIN => \N__53933\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__32721\,
            DIN0 => \RAM_DATA_in_15\,
            DOUT0 => \N__30600\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pon_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53926\,
            DIN => \N__53925\,
            DOUT => \N__53924\,
            PACKAGEPIN => pon_wire
        );

    \pon_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53926\,
            PADOUT => \N__53925\,
            PADIN => \N__53924\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21918\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DAC_sclk_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53917\,
            DIN => \N__53916\,
            DOUT => \N__53915\,
            PACKAGEPIN => \DAC_sclk_wire\
        );

    \DAC_sclk_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53917\,
            PADOUT => \N__53916\,
            PADIN => \N__53915\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21069\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53908\,
            DIN => \N__53907\,
            DOUT => \N__53906\,
            PACKAGEPIN => RAM_DATA(4)
        );

    \RAM_DATA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53908\,
            PADOUT => \N__53907\,
            PADIN => \N__53906\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__27822\,
            DIN0 => \RAM_DATA_in_4\,
            DOUT0 => \N__31572\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53899\,
            DIN => \N__53898\,
            DOUT => \N__53897\,
            PACKAGEPIN => \ADC1_wire\
        );

    \ADC1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53899\,
            PADOUT => \N__53898\,
            PADIN => \N__53897\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_cs_flash_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53890\,
            DIN => \N__53889\,
            DOUT => \N__53888\,
            PACKAGEPIN => spi_cs_flash_wire
        );

    \spi_cs_flash_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53890\,
            PADOUT => \N__53889\,
            PADIN => \N__53888\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__52362\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_miso_flash_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53881\,
            DIN => \N__53880\,
            DOUT => \N__53879\,
            PACKAGEPIN => spi_miso_flash_wire
        );

    \spi_miso_flash_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53881\,
            PADOUT => \N__53880\,
            PADIN => \N__53879\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_miso_flash_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \trig_ext_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53872\,
            DIN => \N__53871\,
            DOUT => \N__53870\,
            PACKAGEPIN => trig_ext_wire
        );

    \trig_ext_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53872\,
            PADOUT => \N__53871\,
            PADIN => \N__53870\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => trig_ext_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53863\,
            DIN => \N__53862\,
            DOUT => \N__53861\,
            PACKAGEPIN => \RAM_ADD_wire\(6)
        );

    \RAM_ADD_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53863\,
            PADOUT => \N__53862\,
            PADIN => \N__53861\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28536\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \top_tour1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53854\,
            DIN => \N__53853\,
            DOUT => \N__53852\,
            PACKAGEPIN => top_tour1_wire
        );

    \top_tour1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53854\,
            PADOUT => \N__53853\,
            PADIN => \N__53852\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => top_tour1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53845\,
            DIN => \N__53844\,
            DOUT => \N__53843\,
            PACKAGEPIN => \RAM_ADD_wire\(17)
        );

    \RAM_ADD_obuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53845\,
            PADOUT => \N__53844\,
            PADIN => \N__53843\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28140\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53836\,
            DIN => \N__53835\,
            DOUT => \N__53834\,
            PACKAGEPIN => \RAM_ADD_wire\(0)
        );

    \RAM_ADD_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53836\,
            PADOUT => \N__53835\,
            PADIN => \N__53834\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29739\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_MODE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53827\,
            DIN => \N__53826\,
            DOUT => \N__53825\,
            PACKAGEPIN => \LED_MODE_wire\
        );

    \LED_MODE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53827\,
            PADOUT => \N__53826\,
            PADIN => \N__53825\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24321\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_nUB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53818\,
            DIN => \N__53817\,
            DOUT => \N__53816\,
            PACKAGEPIN => \RAM_nUB_wire\
        );

    \RAM_nUB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53818\,
            PADOUT => \N__53817\,
            PADIN => \N__53816\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53809\,
            DIN => \N__53808\,
            DOUT => \N__53807\,
            PACKAGEPIN => \RAM_ADD_wire\(11)
        );

    \RAM_ADD_obuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53809\,
            PADOUT => \N__53808\,
            PADIN => \N__53807\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__30381\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53800\,
            DIN => \N__53799\,
            DOUT => \N__53798\,
            PACKAGEPIN => RAM_DATA(14)
        );

    \RAM_DATA_iobuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53800\,
            PADOUT => \N__53799\,
            PADIN => \N__53798\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__32754\,
            DIN0 => \RAM_DATA_in_14\,
            DOUT0 => \N__31230\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DAC_cs_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53791\,
            DIN => \N__53790\,
            DOUT => \N__53789\,
            PACKAGEPIN => \DAC_cs_wire\
        );

    \DAC_cs_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53791\,
            PADOUT => \N__53790\,
            PADIN => \N__53789\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20574\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC8_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53782\,
            DIN => \N__53781\,
            DOUT => \N__53780\,
            PACKAGEPIN => \ADC8_wire\
        );

    \ADC8_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53782\,
            PADOUT => \N__53781\,
            PADIN => \N__53780\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC8_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53773\,
            DIN => \N__53772\,
            DOUT => \N__53771\,
            PACKAGEPIN => RAM_DATA(5)
        );

    \RAM_DATA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53773\,
            PADOUT => \N__53772\,
            PADIN => \N__53771\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__26931\,
            DIN0 => \RAM_DATA_in_5\,
            DOUT0 => \N__30147\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC_clk_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53764\,
            DIN => \N__53763\,
            DOUT => \N__53762\,
            PACKAGEPIN => \ADC_clk_wire\
        );

    \ADC_clk_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53764\,
            PADOUT => \N__53763\,
            PADIN => \N__53762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27615\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53755\,
            DIN => \N__53754\,
            DOUT => \N__53753\,
            PACKAGEPIN => \RAM_ADD_wire\(7)
        );

    \RAM_ADD_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53755\,
            PADOUT => \N__53754\,
            PADIN => \N__53753\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28488\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \poff_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53746\,
            DIN => \N__53745\,
            DOUT => \N__53744\,
            PACKAGEPIN => poff_wire
        );

    \poff_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53746\,
            PADOUT => \N__53745\,
            PADIN => \N__53744\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25335\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC4_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53737\,
            DIN => \N__53736\,
            DOUT => \N__53735\,
            PACKAGEPIN => \ADC4_wire\
        );

    \ADC4_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53737\,
            PADOUT => \N__53736\,
            PADIN => \N__53735\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC4_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC6_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53728\,
            DIN => \N__53727\,
            DOUT => \N__53726\,
            PACKAGEPIN => \ADC6_wire\
        );

    \ADC6_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53728\,
            PADOUT => \N__53727\,
            PADIN => \N__53726\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC6_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53719\,
            DIN => \N__53718\,
            DOUT => \N__53717\,
            PACKAGEPIN => \RAM_ADD_wire\(16)
        );

    \RAM_ADD_obuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53719\,
            PADOUT => \N__53718\,
            PADIN => \N__53717\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28185\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53710\,
            DIN => \N__53709\,
            DOUT => \N__53708\,
            PACKAGEPIN => \RAM_ADD_wire\(1)
        );

    \RAM_ADD_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53710\,
            PADOUT => \N__53709\,
            PADIN => \N__53708\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29664\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC7_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53701\,
            DIN => \N__53700\,
            DOUT => \N__53699\,
            PACKAGEPIN => \ADC7_wire\
        );

    \ADC7_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53701\,
            PADOUT => \N__53700\,
            PADIN => \N__53699\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC7_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \button_mode_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53692\,
            DIN => \N__53691\,
            DOUT => \N__53690\,
            PACKAGEPIN => button_mode_wire
        );

    \button_mode_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53692\,
            PADOUT => \N__53691\,
            PADIN => \N__53690\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => button_mode_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_sclk_ft_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53683\,
            DIN => \N__53682\,
            DOUT => \N__53681\,
            PACKAGEPIN => spi_sclk_ft_wire
        );

    \spi_sclk_ft_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53683\,
            PADOUT => \N__53682\,
            PADIN => \N__53681\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_sclk_ft_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53674\,
            DIN => \N__53673\,
            DOUT => \N__53672\,
            PACKAGEPIN => RAM_DATA(8)
        );

    \RAM_DATA_iobuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53674\,
            PADOUT => \N__53673\,
            PADIN => \N__53672\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__26646\,
            DIN0 => \RAM_DATA_in_8\,
            DOUT0 => \N__30075\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53665\,
            DIN => \N__53664\,
            DOUT => \N__53663\,
            PACKAGEPIN => \RAM_ADD_wire\(10)
        );

    \RAM_ADD_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53665\,
            PADOUT => \N__53664\,
            PADIN => \N__53663\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29616\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53656\,
            DIN => \N__53655\,
            DOUT => \N__53654\,
            PACKAGEPIN => RAM_DATA(13)
        );

    \RAM_DATA_iobuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53656\,
            PADOUT => \N__53655\,
            PADIN => \N__53654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__30522\,
            DIN0 => \RAM_DATA_in_13\,
            DOUT0 => \N__31317\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \trig_ft_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53647\,
            DIN => \N__53646\,
            DOUT => \N__53645\,
            PACKAGEPIN => trig_ft_wire
        );

    \trig_ft_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53647\,
            PADOUT => \N__53646\,
            PADIN => \N__53645\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => trig_ft_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADC9_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53638\,
            DIN => \N__53637\,
            DOUT => \N__53636\,
            PACKAGEPIN => \ADC9_wire\
        );

    \ADC9_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53638\,
            PADOUT => \N__53637\,
            PADIN => \N__53636\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ADC9_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53629\,
            DIN => \N__53628\,
            DOUT => \N__53627\,
            PACKAGEPIN => RAM_DATA(2)
        );

    \RAM_DATA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53629\,
            PADOUT => \N__53628\,
            PADIN => \N__53627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__30447\,
            DIN0 => \RAM_DATA_in_2\,
            DOUT0 => \N__31197\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \cs_rpi2flash_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53620\,
            DIN => \N__53619\,
            DOUT => \N__53618\,
            PACKAGEPIN => cs_rpi2flash_wire
        );

    \cs_rpi2flash_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53620\,
            PADOUT => \N__53619\,
            PADIN => \N__53618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => cs_rpi2flash_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53611\,
            DIN => \N__53610\,
            DOUT => \N__53609\,
            PACKAGEPIN => \LED3_wire\
        );

    \LED3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53611\,
            PADOUT => \N__53610\,
            PADIN => \N__53609\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32583\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_mosi_ft_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53602\,
            DIN => \N__53601\,
            DOUT => \N__53600\,
            PACKAGEPIN => spi_mosi_ft_wire
        );

    \spi_mosi_ft_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53602\,
            PADOUT => \N__53601\,
            PADIN => \N__53600\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_mosi_ft_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_nOE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53593\,
            DIN => \N__53592\,
            DOUT => \N__53591\,
            PACKAGEPIN => \RAM_nOE_wire\
        );

    \RAM_nOE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53593\,
            PADOUT => \N__53592\,
            PADIN => \N__53591\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53584\,
            DIN => \N__53583\,
            DOUT => \N__53582\,
            PACKAGEPIN => \RAM_ADD_wire\(4)
        );

    \RAM_ADD_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53584\,
            PADOUT => \N__53583\,
            PADIN => \N__53582\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28626\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53575\,
            DIN => \N__53574\,
            DOUT => \N__53573\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53575\,
            PADOUT => \N__53574\,
            PADIN => \N__53573\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \top_tour2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53566\,
            DIN => \N__53565\,
            DOUT => \N__53564\,
            PACKAGEPIN => top_tour2_wire
        );

    \top_tour2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53566\,
            PADOUT => \N__53565\,
            PADIN => \N__53564\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => top_tour2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_cs_rpi_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53557\,
            DIN => \N__53556\,
            DOUT => \N__53555\,
            PACKAGEPIN => spi_cs_rpi_wire
        );

    \spi_cs_rpi_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53557\,
            PADOUT => \N__53556\,
            PADIN => \N__53555\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_cs_rpi_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53548\,
            DIN => \N__53547\,
            DOUT => \N__53546\,
            PACKAGEPIN => \RAM_ADD_wire\(15)
        );

    \RAM_ADD_obuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53548\,
            PADOUT => \N__53547\,
            PADIN => \N__53546\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28230\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_miso_rpi_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53539\,
            DIN => \N__53538\,
            DOUT => \N__53537\,
            PACKAGEPIN => spi_miso_rpi_wire
        );

    \spi_miso_rpi_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53539\,
            PADOUT => \N__53538\,
            PADIN => \N__53537\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33120\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53530\,
            DIN => \N__53529\,
            DOUT => \N__53528\,
            PACKAGEPIN => RAM_DATA(9)
        );

    \RAM_DATA_iobuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53530\,
            PADOUT => \N__53529\,
            PADIN => \N__53528\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__28362\,
            DIN0 => \RAM_DATA_in_9\,
            DOUT0 => \N__30624\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53521\,
            DIN => \N__53520\,
            DOUT => \N__53519\,
            PACKAGEPIN => \RAM_ADD_wire\(8)
        );

    \RAM_ADD_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53521\,
            PADOUT => \N__53520\,
            PADIN => \N__53519\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28440\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53512\,
            DIN => \N__53511\,
            DOUT => \N__53510\,
            PACKAGEPIN => RAM_DATA(12)
        );

    \RAM_DATA_iobuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53512\,
            PADOUT => \N__53511\,
            PADIN => \N__53510\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__26898\,
            DIN0 => \RAM_DATA_in_12\,
            DOUT0 => \N__31413\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_DATA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53503\,
            DIN => \N__53502\,
            DOUT => \N__53501\,
            PACKAGEPIN => RAM_DATA(3)
        );

    \RAM_DATA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__53503\,
            PADOUT => \N__53502\,
            PADIN => \N__53501\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__27792\,
            DIN0 => \RAM_DATA_in_3\,
            DOUT0 => \N__30222\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_cs_ft_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53494\,
            DIN => \N__53493\,
            DOUT => \N__53492\,
            PACKAGEPIN => spi_cs_ft_wire
        );

    \spi_cs_ft_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__53494\,
            PADOUT => \N__53493\,
            PADIN => \N__53492\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => spi_cs_ft_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \spi_mosi_flash_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53485\,
            DIN => \N__53484\,
            DOUT => \N__53483\,
            PACKAGEPIN => spi_mosi_flash_wire
        );

    \spi_mosi_flash_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53485\,
            PADOUT => \N__53484\,
            PADIN => \N__53483\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__52563\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAM_ADD_obuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53476\,
            DIN => \N__53475\,
            DOUT => \N__53474\,
            PACKAGEPIN => \RAM_ADD_wire\(14)
        );

    \RAM_ADD_obuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__53476\,
            PADOUT => \N__53475\,
            PADIN => \N__53474\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__28275\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__12722\ : InMux
    port map (
            O => \N__53457\,
            I => \N__53454\
        );

    \I__12721\ : LocalMux
    port map (
            O => \N__53454\,
            I => op_eq_scounterdac10_0_a2_0
        );

    \I__12720\ : InMux
    port map (
            O => \N__53451\,
            I => \N__53446\
        );

    \I__12719\ : InMux
    port map (
            O => \N__53450\,
            I => \N__53443\
        );

    \I__12718\ : InMux
    port map (
            O => \N__53449\,
            I => \N__53440\
        );

    \I__12717\ : LocalMux
    port map (
            O => \N__53446\,
            I => \N__53437\
        );

    \I__12716\ : LocalMux
    port map (
            O => \N__53443\,
            I => \N__53433\
        );

    \I__12715\ : LocalMux
    port map (
            O => \N__53440\,
            I => \N__53430\
        );

    \I__12714\ : Span4Mux_v
    port map (
            O => \N__53437\,
            I => \N__53427\
        );

    \I__12713\ : InMux
    port map (
            O => \N__53436\,
            I => \N__53424\
        );

    \I__12712\ : Odrv4
    port map (
            O => \N__53433\,
            I => \N_23\
        );

    \I__12711\ : Odrv4
    port map (
            O => \N__53430\,
            I => \N_23\
        );

    \I__12710\ : Odrv4
    port map (
            O => \N__53427\,
            I => \N_23\
        );

    \I__12709\ : LocalMux
    port map (
            O => \N__53424\,
            I => \N_23\
        );

    \I__12708\ : CascadeMux
    port map (
            O => \N__53415\,
            I => \N__53411\
        );

    \I__12707\ : CascadeMux
    port map (
            O => \N__53414\,
            I => \N__53407\
        );

    \I__12706\ : InMux
    port map (
            O => \N__53411\,
            I => \N__53402\
        );

    \I__12705\ : InMux
    port map (
            O => \N__53410\,
            I => \N__53399\
        );

    \I__12704\ : InMux
    port map (
            O => \N__53407\,
            I => \N__53396\
        );

    \I__12703\ : InMux
    port map (
            O => \N__53406\,
            I => \N__53390\
        );

    \I__12702\ : InMux
    port map (
            O => \N__53405\,
            I => \N__53390\
        );

    \I__12701\ : LocalMux
    port map (
            O => \N__53402\,
            I => \N__53387\
        );

    \I__12700\ : LocalMux
    port map (
            O => \N__53399\,
            I => \N__53382\
        );

    \I__12699\ : LocalMux
    port map (
            O => \N__53396\,
            I => \N__53382\
        );

    \I__12698\ : CascadeMux
    port map (
            O => \N__53395\,
            I => \N__53379\
        );

    \I__12697\ : LocalMux
    port map (
            O => \N__53390\,
            I => \N__53372\
        );

    \I__12696\ : Span4Mux_v
    port map (
            O => \N__53387\,
            I => \N__53372\
        );

    \I__12695\ : Span4Mux_v
    port map (
            O => \N__53382\,
            I => \N__53372\
        );

    \I__12694\ : InMux
    port map (
            O => \N__53379\,
            I => \N__53369\
        );

    \I__12693\ : Odrv4
    port map (
            O => \N__53372\,
            I => \sCounterDACZ0Z_0\
        );

    \I__12692\ : LocalMux
    port map (
            O => \N__53369\,
            I => \sCounterDACZ0Z_0\
        );

    \I__12691\ : InMux
    port map (
            O => \N__53364\,
            I => \N__53361\
        );

    \I__12690\ : LocalMux
    port map (
            O => \N__53361\,
            I => \N__53358\
        );

    \I__12689\ : Span4Mux_v
    port map (
            O => \N__53358\,
            I => \N__53354\
        );

    \I__12688\ : InMux
    port map (
            O => \N__53357\,
            I => \N__53351\
        );

    \I__12687\ : Odrv4
    port map (
            O => \N__53354\,
            I => \N_22\
        );

    \I__12686\ : LocalMux
    port map (
            O => \N__53351\,
            I => \N_22\
        );

    \I__12685\ : IoInMux
    port map (
            O => \N__53346\,
            I => \N__53343\
        );

    \I__12684\ : LocalMux
    port map (
            O => \N__53343\,
            I => \N__53340\
        );

    \I__12683\ : Odrv12
    port map (
            O => \N__53340\,
            I => op_eq_scounterdac10
        );

    \I__12682\ : InMux
    port map (
            O => \N__53337\,
            I => \N__53332\
        );

    \I__12681\ : InMux
    port map (
            O => \N__53336\,
            I => \N__53326\
        );

    \I__12680\ : InMux
    port map (
            O => \N__53335\,
            I => \N__53326\
        );

    \I__12679\ : LocalMux
    port map (
            O => \N__53332\,
            I => \N__53323\
        );

    \I__12678\ : InMux
    port map (
            O => \N__53331\,
            I => \N__53319\
        );

    \I__12677\ : LocalMux
    port map (
            O => \N__53326\,
            I => \N__53316\
        );

    \I__12676\ : Span12Mux_h
    port map (
            O => \N__53323\,
            I => \N__53313\
        );

    \I__12675\ : InMux
    port map (
            O => \N__53322\,
            I => \N__53310\
        );

    \I__12674\ : LocalMux
    port map (
            O => \N__53319\,
            I => \N__53305\
        );

    \I__12673\ : Span4Mux_h
    port map (
            O => \N__53316\,
            I => \N__53305\
        );

    \I__12672\ : Odrv12
    port map (
            O => \N__53313\,
            I => \sCounterDACZ0Z_8\
        );

    \I__12671\ : LocalMux
    port map (
            O => \N__53310\,
            I => \sCounterDACZ0Z_8\
        );

    \I__12670\ : Odrv4
    port map (
            O => \N__53305\,
            I => \sCounterDACZ0Z_8\
        );

    \I__12669\ : InMux
    port map (
            O => \N__53298\,
            I => \N__53295\
        );

    \I__12668\ : LocalMux
    port map (
            O => \N__53295\,
            I => \N__53292\
        );

    \I__12667\ : Odrv4
    port map (
            O => \N__53292\,
            I => \un2_scounterdac_cry_7_THRU_CO\
        );

    \I__12666\ : InMux
    port map (
            O => \N__53289\,
            I => un2_scounterdac_cry_7
        );

    \I__12665\ : InMux
    port map (
            O => \N__53286\,
            I => \bfn_22_11_0_\
        );

    \I__12664\ : ClkMux
    port map (
            O => \N__53283\,
            I => \N__53154\
        );

    \I__12663\ : ClkMux
    port map (
            O => \N__53282\,
            I => \N__53154\
        );

    \I__12662\ : ClkMux
    port map (
            O => \N__53281\,
            I => \N__53154\
        );

    \I__12661\ : ClkMux
    port map (
            O => \N__53280\,
            I => \N__53154\
        );

    \I__12660\ : ClkMux
    port map (
            O => \N__53279\,
            I => \N__53154\
        );

    \I__12659\ : ClkMux
    port map (
            O => \N__53278\,
            I => \N__53154\
        );

    \I__12658\ : ClkMux
    port map (
            O => \N__53277\,
            I => \N__53154\
        );

    \I__12657\ : ClkMux
    port map (
            O => \N__53276\,
            I => \N__53154\
        );

    \I__12656\ : ClkMux
    port map (
            O => \N__53275\,
            I => \N__53154\
        );

    \I__12655\ : ClkMux
    port map (
            O => \N__53274\,
            I => \N__53154\
        );

    \I__12654\ : ClkMux
    port map (
            O => \N__53273\,
            I => \N__53154\
        );

    \I__12653\ : ClkMux
    port map (
            O => \N__53272\,
            I => \N__53154\
        );

    \I__12652\ : ClkMux
    port map (
            O => \N__53271\,
            I => \N__53154\
        );

    \I__12651\ : ClkMux
    port map (
            O => \N__53270\,
            I => \N__53154\
        );

    \I__12650\ : ClkMux
    port map (
            O => \N__53269\,
            I => \N__53154\
        );

    \I__12649\ : ClkMux
    port map (
            O => \N__53268\,
            I => \N__53154\
        );

    \I__12648\ : ClkMux
    port map (
            O => \N__53267\,
            I => \N__53154\
        );

    \I__12647\ : ClkMux
    port map (
            O => \N__53266\,
            I => \N__53154\
        );

    \I__12646\ : ClkMux
    port map (
            O => \N__53265\,
            I => \N__53154\
        );

    \I__12645\ : ClkMux
    port map (
            O => \N__53264\,
            I => \N__53154\
        );

    \I__12644\ : ClkMux
    port map (
            O => \N__53263\,
            I => \N__53154\
        );

    \I__12643\ : ClkMux
    port map (
            O => \N__53262\,
            I => \N__53154\
        );

    \I__12642\ : ClkMux
    port map (
            O => \N__53261\,
            I => \N__53154\
        );

    \I__12641\ : ClkMux
    port map (
            O => \N__53260\,
            I => \N__53154\
        );

    \I__12640\ : ClkMux
    port map (
            O => \N__53259\,
            I => \N__53154\
        );

    \I__12639\ : ClkMux
    port map (
            O => \N__53258\,
            I => \N__53154\
        );

    \I__12638\ : ClkMux
    port map (
            O => \N__53257\,
            I => \N__53154\
        );

    \I__12637\ : ClkMux
    port map (
            O => \N__53256\,
            I => \N__53154\
        );

    \I__12636\ : ClkMux
    port map (
            O => \N__53255\,
            I => \N__53154\
        );

    \I__12635\ : ClkMux
    port map (
            O => \N__53254\,
            I => \N__53154\
        );

    \I__12634\ : ClkMux
    port map (
            O => \N__53253\,
            I => \N__53154\
        );

    \I__12633\ : ClkMux
    port map (
            O => \N__53252\,
            I => \N__53154\
        );

    \I__12632\ : ClkMux
    port map (
            O => \N__53251\,
            I => \N__53154\
        );

    \I__12631\ : ClkMux
    port map (
            O => \N__53250\,
            I => \N__53154\
        );

    \I__12630\ : ClkMux
    port map (
            O => \N__53249\,
            I => \N__53154\
        );

    \I__12629\ : ClkMux
    port map (
            O => \N__53248\,
            I => \N__53154\
        );

    \I__12628\ : ClkMux
    port map (
            O => \N__53247\,
            I => \N__53154\
        );

    \I__12627\ : ClkMux
    port map (
            O => \N__53246\,
            I => \N__53154\
        );

    \I__12626\ : ClkMux
    port map (
            O => \N__53245\,
            I => \N__53154\
        );

    \I__12625\ : ClkMux
    port map (
            O => \N__53244\,
            I => \N__53154\
        );

    \I__12624\ : ClkMux
    port map (
            O => \N__53243\,
            I => \N__53154\
        );

    \I__12623\ : ClkMux
    port map (
            O => \N__53242\,
            I => \N__53154\
        );

    \I__12622\ : ClkMux
    port map (
            O => \N__53241\,
            I => \N__53154\
        );

    \I__12621\ : GlobalMux
    port map (
            O => \N__53154\,
            I => \N__53151\
        );

    \I__12620\ : gio2CtrlBuf
    port map (
            O => \N__53151\,
            I => pll_clk64_0_g
        );

    \I__12619\ : SRMux
    port map (
            O => \N__53148\,
            I => \N__52602\
        );

    \I__12618\ : SRMux
    port map (
            O => \N__53147\,
            I => \N__52602\
        );

    \I__12617\ : SRMux
    port map (
            O => \N__53146\,
            I => \N__52602\
        );

    \I__12616\ : SRMux
    port map (
            O => \N__53145\,
            I => \N__52602\
        );

    \I__12615\ : SRMux
    port map (
            O => \N__53144\,
            I => \N__52602\
        );

    \I__12614\ : SRMux
    port map (
            O => \N__53143\,
            I => \N__52602\
        );

    \I__12613\ : SRMux
    port map (
            O => \N__53142\,
            I => \N__52602\
        );

    \I__12612\ : SRMux
    port map (
            O => \N__53141\,
            I => \N__52602\
        );

    \I__12611\ : SRMux
    port map (
            O => \N__53140\,
            I => \N__52602\
        );

    \I__12610\ : SRMux
    port map (
            O => \N__53139\,
            I => \N__52602\
        );

    \I__12609\ : SRMux
    port map (
            O => \N__53138\,
            I => \N__52602\
        );

    \I__12608\ : SRMux
    port map (
            O => \N__53137\,
            I => \N__52602\
        );

    \I__12607\ : SRMux
    port map (
            O => \N__53136\,
            I => \N__52602\
        );

    \I__12606\ : SRMux
    port map (
            O => \N__53135\,
            I => \N__52602\
        );

    \I__12605\ : SRMux
    port map (
            O => \N__53134\,
            I => \N__52602\
        );

    \I__12604\ : SRMux
    port map (
            O => \N__53133\,
            I => \N__52602\
        );

    \I__12603\ : SRMux
    port map (
            O => \N__53132\,
            I => \N__52602\
        );

    \I__12602\ : SRMux
    port map (
            O => \N__53131\,
            I => \N__52602\
        );

    \I__12601\ : SRMux
    port map (
            O => \N__53130\,
            I => \N__52602\
        );

    \I__12600\ : SRMux
    port map (
            O => \N__53129\,
            I => \N__52602\
        );

    \I__12599\ : SRMux
    port map (
            O => \N__53128\,
            I => \N__52602\
        );

    \I__12598\ : SRMux
    port map (
            O => \N__53127\,
            I => \N__52602\
        );

    \I__12597\ : SRMux
    port map (
            O => \N__53126\,
            I => \N__52602\
        );

    \I__12596\ : SRMux
    port map (
            O => \N__53125\,
            I => \N__52602\
        );

    \I__12595\ : SRMux
    port map (
            O => \N__53124\,
            I => \N__52602\
        );

    \I__12594\ : SRMux
    port map (
            O => \N__53123\,
            I => \N__52602\
        );

    \I__12593\ : SRMux
    port map (
            O => \N__53122\,
            I => \N__52602\
        );

    \I__12592\ : SRMux
    port map (
            O => \N__53121\,
            I => \N__52602\
        );

    \I__12591\ : SRMux
    port map (
            O => \N__53120\,
            I => \N__52602\
        );

    \I__12590\ : SRMux
    port map (
            O => \N__53119\,
            I => \N__52602\
        );

    \I__12589\ : SRMux
    port map (
            O => \N__53118\,
            I => \N__52602\
        );

    \I__12588\ : SRMux
    port map (
            O => \N__53117\,
            I => \N__52602\
        );

    \I__12587\ : SRMux
    port map (
            O => \N__53116\,
            I => \N__52602\
        );

    \I__12586\ : SRMux
    port map (
            O => \N__53115\,
            I => \N__52602\
        );

    \I__12585\ : SRMux
    port map (
            O => \N__53114\,
            I => \N__52602\
        );

    \I__12584\ : SRMux
    port map (
            O => \N__53113\,
            I => \N__52602\
        );

    \I__12583\ : SRMux
    port map (
            O => \N__53112\,
            I => \N__52602\
        );

    \I__12582\ : SRMux
    port map (
            O => \N__53111\,
            I => \N__52602\
        );

    \I__12581\ : SRMux
    port map (
            O => \N__53110\,
            I => \N__52602\
        );

    \I__12580\ : SRMux
    port map (
            O => \N__53109\,
            I => \N__52602\
        );

    \I__12579\ : SRMux
    port map (
            O => \N__53108\,
            I => \N__52602\
        );

    \I__12578\ : SRMux
    port map (
            O => \N__53107\,
            I => \N__52602\
        );

    \I__12577\ : SRMux
    port map (
            O => \N__53106\,
            I => \N__52602\
        );

    \I__12576\ : SRMux
    port map (
            O => \N__53105\,
            I => \N__52602\
        );

    \I__12575\ : SRMux
    port map (
            O => \N__53104\,
            I => \N__52602\
        );

    \I__12574\ : SRMux
    port map (
            O => \N__53103\,
            I => \N__52602\
        );

    \I__12573\ : SRMux
    port map (
            O => \N__53102\,
            I => \N__52602\
        );

    \I__12572\ : SRMux
    port map (
            O => \N__53101\,
            I => \N__52602\
        );

    \I__12571\ : SRMux
    port map (
            O => \N__53100\,
            I => \N__52602\
        );

    \I__12570\ : SRMux
    port map (
            O => \N__53099\,
            I => \N__52602\
        );

    \I__12569\ : SRMux
    port map (
            O => \N__53098\,
            I => \N__52602\
        );

    \I__12568\ : SRMux
    port map (
            O => \N__53097\,
            I => \N__52602\
        );

    \I__12567\ : SRMux
    port map (
            O => \N__53096\,
            I => \N__52602\
        );

    \I__12566\ : SRMux
    port map (
            O => \N__53095\,
            I => \N__52602\
        );

    \I__12565\ : SRMux
    port map (
            O => \N__53094\,
            I => \N__52602\
        );

    \I__12564\ : SRMux
    port map (
            O => \N__53093\,
            I => \N__52602\
        );

    \I__12563\ : SRMux
    port map (
            O => \N__53092\,
            I => \N__52602\
        );

    \I__12562\ : SRMux
    port map (
            O => \N__53091\,
            I => \N__52602\
        );

    \I__12561\ : SRMux
    port map (
            O => \N__53090\,
            I => \N__52602\
        );

    \I__12560\ : SRMux
    port map (
            O => \N__53089\,
            I => \N__52602\
        );

    \I__12559\ : SRMux
    port map (
            O => \N__53088\,
            I => \N__52602\
        );

    \I__12558\ : SRMux
    port map (
            O => \N__53087\,
            I => \N__52602\
        );

    \I__12557\ : SRMux
    port map (
            O => \N__53086\,
            I => \N__52602\
        );

    \I__12556\ : SRMux
    port map (
            O => \N__53085\,
            I => \N__52602\
        );

    \I__12555\ : SRMux
    port map (
            O => \N__53084\,
            I => \N__52602\
        );

    \I__12554\ : SRMux
    port map (
            O => \N__53083\,
            I => \N__52602\
        );

    \I__12553\ : SRMux
    port map (
            O => \N__53082\,
            I => \N__52602\
        );

    \I__12552\ : SRMux
    port map (
            O => \N__53081\,
            I => \N__52602\
        );

    \I__12551\ : SRMux
    port map (
            O => \N__53080\,
            I => \N__52602\
        );

    \I__12550\ : SRMux
    port map (
            O => \N__53079\,
            I => \N__52602\
        );

    \I__12549\ : SRMux
    port map (
            O => \N__53078\,
            I => \N__52602\
        );

    \I__12548\ : SRMux
    port map (
            O => \N__53077\,
            I => \N__52602\
        );

    \I__12547\ : SRMux
    port map (
            O => \N__53076\,
            I => \N__52602\
        );

    \I__12546\ : SRMux
    port map (
            O => \N__53075\,
            I => \N__52602\
        );

    \I__12545\ : SRMux
    port map (
            O => \N__53074\,
            I => \N__52602\
        );

    \I__12544\ : SRMux
    port map (
            O => \N__53073\,
            I => \N__52602\
        );

    \I__12543\ : SRMux
    port map (
            O => \N__53072\,
            I => \N__52602\
        );

    \I__12542\ : SRMux
    port map (
            O => \N__53071\,
            I => \N__52602\
        );

    \I__12541\ : SRMux
    port map (
            O => \N__53070\,
            I => \N__52602\
        );

    \I__12540\ : SRMux
    port map (
            O => \N__53069\,
            I => \N__52602\
        );

    \I__12539\ : SRMux
    port map (
            O => \N__53068\,
            I => \N__52602\
        );

    \I__12538\ : SRMux
    port map (
            O => \N__53067\,
            I => \N__52602\
        );

    \I__12537\ : SRMux
    port map (
            O => \N__53066\,
            I => \N__52602\
        );

    \I__12536\ : SRMux
    port map (
            O => \N__53065\,
            I => \N__52602\
        );

    \I__12535\ : SRMux
    port map (
            O => \N__53064\,
            I => \N__52602\
        );

    \I__12534\ : SRMux
    port map (
            O => \N__53063\,
            I => \N__52602\
        );

    \I__12533\ : SRMux
    port map (
            O => \N__53062\,
            I => \N__52602\
        );

    \I__12532\ : SRMux
    port map (
            O => \N__53061\,
            I => \N__52602\
        );

    \I__12531\ : SRMux
    port map (
            O => \N__53060\,
            I => \N__52602\
        );

    \I__12530\ : SRMux
    port map (
            O => \N__53059\,
            I => \N__52602\
        );

    \I__12529\ : SRMux
    port map (
            O => \N__53058\,
            I => \N__52602\
        );

    \I__12528\ : SRMux
    port map (
            O => \N__53057\,
            I => \N__52602\
        );

    \I__12527\ : SRMux
    port map (
            O => \N__53056\,
            I => \N__52602\
        );

    \I__12526\ : SRMux
    port map (
            O => \N__53055\,
            I => \N__52602\
        );

    \I__12525\ : SRMux
    port map (
            O => \N__53054\,
            I => \N__52602\
        );

    \I__12524\ : SRMux
    port map (
            O => \N__53053\,
            I => \N__52602\
        );

    \I__12523\ : SRMux
    port map (
            O => \N__53052\,
            I => \N__52602\
        );

    \I__12522\ : SRMux
    port map (
            O => \N__53051\,
            I => \N__52602\
        );

    \I__12521\ : SRMux
    port map (
            O => \N__53050\,
            I => \N__52602\
        );

    \I__12520\ : SRMux
    port map (
            O => \N__53049\,
            I => \N__52602\
        );

    \I__12519\ : SRMux
    port map (
            O => \N__53048\,
            I => \N__52602\
        );

    \I__12518\ : SRMux
    port map (
            O => \N__53047\,
            I => \N__52602\
        );

    \I__12517\ : SRMux
    port map (
            O => \N__53046\,
            I => \N__52602\
        );

    \I__12516\ : SRMux
    port map (
            O => \N__53045\,
            I => \N__52602\
        );

    \I__12515\ : SRMux
    port map (
            O => \N__53044\,
            I => \N__52602\
        );

    \I__12514\ : SRMux
    port map (
            O => \N__53043\,
            I => \N__52602\
        );

    \I__12513\ : SRMux
    port map (
            O => \N__53042\,
            I => \N__52602\
        );

    \I__12512\ : SRMux
    port map (
            O => \N__53041\,
            I => \N__52602\
        );

    \I__12511\ : SRMux
    port map (
            O => \N__53040\,
            I => \N__52602\
        );

    \I__12510\ : SRMux
    port map (
            O => \N__53039\,
            I => \N__52602\
        );

    \I__12509\ : SRMux
    port map (
            O => \N__53038\,
            I => \N__52602\
        );

    \I__12508\ : SRMux
    port map (
            O => \N__53037\,
            I => \N__52602\
        );

    \I__12507\ : SRMux
    port map (
            O => \N__53036\,
            I => \N__52602\
        );

    \I__12506\ : SRMux
    port map (
            O => \N__53035\,
            I => \N__52602\
        );

    \I__12505\ : SRMux
    port map (
            O => \N__53034\,
            I => \N__52602\
        );

    \I__12504\ : SRMux
    port map (
            O => \N__53033\,
            I => \N__52602\
        );

    \I__12503\ : SRMux
    port map (
            O => \N__53032\,
            I => \N__52602\
        );

    \I__12502\ : SRMux
    port map (
            O => \N__53031\,
            I => \N__52602\
        );

    \I__12501\ : SRMux
    port map (
            O => \N__53030\,
            I => \N__52602\
        );

    \I__12500\ : SRMux
    port map (
            O => \N__53029\,
            I => \N__52602\
        );

    \I__12499\ : SRMux
    port map (
            O => \N__53028\,
            I => \N__52602\
        );

    \I__12498\ : SRMux
    port map (
            O => \N__53027\,
            I => \N__52602\
        );

    \I__12497\ : SRMux
    port map (
            O => \N__53026\,
            I => \N__52602\
        );

    \I__12496\ : SRMux
    port map (
            O => \N__53025\,
            I => \N__52602\
        );

    \I__12495\ : SRMux
    port map (
            O => \N__53024\,
            I => \N__52602\
        );

    \I__12494\ : SRMux
    port map (
            O => \N__53023\,
            I => \N__52602\
        );

    \I__12493\ : SRMux
    port map (
            O => \N__53022\,
            I => \N__52602\
        );

    \I__12492\ : SRMux
    port map (
            O => \N__53021\,
            I => \N__52602\
        );

    \I__12491\ : SRMux
    port map (
            O => \N__53020\,
            I => \N__52602\
        );

    \I__12490\ : SRMux
    port map (
            O => \N__53019\,
            I => \N__52602\
        );

    \I__12489\ : SRMux
    port map (
            O => \N__53018\,
            I => \N__52602\
        );

    \I__12488\ : SRMux
    port map (
            O => \N__53017\,
            I => \N__52602\
        );

    \I__12487\ : SRMux
    port map (
            O => \N__53016\,
            I => \N__52602\
        );

    \I__12486\ : SRMux
    port map (
            O => \N__53015\,
            I => \N__52602\
        );

    \I__12485\ : SRMux
    port map (
            O => \N__53014\,
            I => \N__52602\
        );

    \I__12484\ : SRMux
    port map (
            O => \N__53013\,
            I => \N__52602\
        );

    \I__12483\ : SRMux
    port map (
            O => \N__53012\,
            I => \N__52602\
        );

    \I__12482\ : SRMux
    port map (
            O => \N__53011\,
            I => \N__52602\
        );

    \I__12481\ : SRMux
    port map (
            O => \N__53010\,
            I => \N__52602\
        );

    \I__12480\ : SRMux
    port map (
            O => \N__53009\,
            I => \N__52602\
        );

    \I__12479\ : SRMux
    port map (
            O => \N__53008\,
            I => \N__52602\
        );

    \I__12478\ : SRMux
    port map (
            O => \N__53007\,
            I => \N__52602\
        );

    \I__12477\ : SRMux
    port map (
            O => \N__53006\,
            I => \N__52602\
        );

    \I__12476\ : SRMux
    port map (
            O => \N__53005\,
            I => \N__52602\
        );

    \I__12475\ : SRMux
    port map (
            O => \N__53004\,
            I => \N__52602\
        );

    \I__12474\ : SRMux
    port map (
            O => \N__53003\,
            I => \N__52602\
        );

    \I__12473\ : SRMux
    port map (
            O => \N__53002\,
            I => \N__52602\
        );

    \I__12472\ : SRMux
    port map (
            O => \N__53001\,
            I => \N__52602\
        );

    \I__12471\ : SRMux
    port map (
            O => \N__53000\,
            I => \N__52602\
        );

    \I__12470\ : SRMux
    port map (
            O => \N__52999\,
            I => \N__52602\
        );

    \I__12469\ : SRMux
    port map (
            O => \N__52998\,
            I => \N__52602\
        );

    \I__12468\ : SRMux
    port map (
            O => \N__52997\,
            I => \N__52602\
        );

    \I__12467\ : SRMux
    port map (
            O => \N__52996\,
            I => \N__52602\
        );

    \I__12466\ : SRMux
    port map (
            O => \N__52995\,
            I => \N__52602\
        );

    \I__12465\ : SRMux
    port map (
            O => \N__52994\,
            I => \N__52602\
        );

    \I__12464\ : SRMux
    port map (
            O => \N__52993\,
            I => \N__52602\
        );

    \I__12463\ : SRMux
    port map (
            O => \N__52992\,
            I => \N__52602\
        );

    \I__12462\ : SRMux
    port map (
            O => \N__52991\,
            I => \N__52602\
        );

    \I__12461\ : SRMux
    port map (
            O => \N__52990\,
            I => \N__52602\
        );

    \I__12460\ : SRMux
    port map (
            O => \N__52989\,
            I => \N__52602\
        );

    \I__12459\ : SRMux
    port map (
            O => \N__52988\,
            I => \N__52602\
        );

    \I__12458\ : SRMux
    port map (
            O => \N__52987\,
            I => \N__52602\
        );

    \I__12457\ : SRMux
    port map (
            O => \N__52986\,
            I => \N__52602\
        );

    \I__12456\ : SRMux
    port map (
            O => \N__52985\,
            I => \N__52602\
        );

    \I__12455\ : SRMux
    port map (
            O => \N__52984\,
            I => \N__52602\
        );

    \I__12454\ : SRMux
    port map (
            O => \N__52983\,
            I => \N__52602\
        );

    \I__12453\ : SRMux
    port map (
            O => \N__52982\,
            I => \N__52602\
        );

    \I__12452\ : SRMux
    port map (
            O => \N__52981\,
            I => \N__52602\
        );

    \I__12451\ : SRMux
    port map (
            O => \N__52980\,
            I => \N__52602\
        );

    \I__12450\ : SRMux
    port map (
            O => \N__52979\,
            I => \N__52602\
        );

    \I__12449\ : SRMux
    port map (
            O => \N__52978\,
            I => \N__52602\
        );

    \I__12448\ : SRMux
    port map (
            O => \N__52977\,
            I => \N__52602\
        );

    \I__12447\ : SRMux
    port map (
            O => \N__52976\,
            I => \N__52602\
        );

    \I__12446\ : SRMux
    port map (
            O => \N__52975\,
            I => \N__52602\
        );

    \I__12445\ : SRMux
    port map (
            O => \N__52974\,
            I => \N__52602\
        );

    \I__12444\ : SRMux
    port map (
            O => \N__52973\,
            I => \N__52602\
        );

    \I__12443\ : SRMux
    port map (
            O => \N__52972\,
            I => \N__52602\
        );

    \I__12442\ : SRMux
    port map (
            O => \N__52971\,
            I => \N__52602\
        );

    \I__12441\ : SRMux
    port map (
            O => \N__52970\,
            I => \N__52602\
        );

    \I__12440\ : SRMux
    port map (
            O => \N__52969\,
            I => \N__52602\
        );

    \I__12439\ : SRMux
    port map (
            O => \N__52968\,
            I => \N__52602\
        );

    \I__12438\ : SRMux
    port map (
            O => \N__52967\,
            I => \N__52602\
        );

    \I__12437\ : GlobalMux
    port map (
            O => \N__52602\,
            I => \N__52599\
        );

    \I__12436\ : gio2CtrlBuf
    port map (
            O => \N__52599\,
            I => \LED3_c_i_g\
        );

    \I__12435\ : InMux
    port map (
            O => \N__52596\,
            I => \N__52593\
        );

    \I__12434\ : LocalMux
    port map (
            O => \N__52593\,
            I => \N__52589\
        );

    \I__12433\ : InMux
    port map (
            O => \N__52592\,
            I => \N__52586\
        );

    \I__12432\ : Span4Mux_v
    port map (
            O => \N__52589\,
            I => \N__52583\
        );

    \I__12431\ : LocalMux
    port map (
            O => \N__52586\,
            I => \N__52580\
        );

    \I__12430\ : Sp12to4
    port map (
            O => \N__52583\,
            I => \N__52577\
        );

    \I__12429\ : Span4Mux_v
    port map (
            O => \N__52580\,
            I => \N__52574\
        );

    \I__12428\ : Span12Mux_h
    port map (
            O => \N__52577\,
            I => \N__52569\
        );

    \I__12427\ : Sp12to4
    port map (
            O => \N__52574\,
            I => \N__52569\
        );

    \I__12426\ : Span12Mux_h
    port map (
            O => \N__52569\,
            I => \N__52566\
        );

    \I__12425\ : Odrv12
    port map (
            O => \N__52566\,
            I => spi_mosi_rpi_c
        );

    \I__12424\ : IoInMux
    port map (
            O => \N__52563\,
            I => \N__52560\
        );

    \I__12423\ : LocalMux
    port map (
            O => \N__52560\,
            I => \N__52557\
        );

    \I__12422\ : Span4Mux_s2_v
    port map (
            O => \N__52557\,
            I => \N__52554\
        );

    \I__12421\ : Span4Mux_v
    port map (
            O => \N__52554\,
            I => \N__52551\
        );

    \I__12420\ : Odrv4
    port map (
            O => \N__52551\,
            I => spi_mosi_flash_c
        );

    \I__12419\ : InMux
    port map (
            O => \N__52548\,
            I => \N__52542\
        );

    \I__12418\ : InMux
    port map (
            O => \N__52547\,
            I => \N__52542\
        );

    \I__12417\ : LocalMux
    port map (
            O => \N__52542\,
            I => \N__52537\
        );

    \I__12416\ : InMux
    port map (
            O => \N__52541\,
            I => \N__52534\
        );

    \I__12415\ : InMux
    port map (
            O => \N__52540\,
            I => \N__52531\
        );

    \I__12414\ : Odrv4
    port map (
            O => \N__52537\,
            I => \sCounterDACZ0Z_4\
        );

    \I__12413\ : LocalMux
    port map (
            O => \N__52534\,
            I => \sCounterDACZ0Z_4\
        );

    \I__12412\ : LocalMux
    port map (
            O => \N__52531\,
            I => \sCounterDACZ0Z_4\
        );

    \I__12411\ : InMux
    port map (
            O => \N__52524\,
            I => \N__52521\
        );

    \I__12410\ : LocalMux
    port map (
            O => \N__52521\,
            I => \N__52516\
        );

    \I__12409\ : InMux
    port map (
            O => \N__52520\,
            I => \N__52513\
        );

    \I__12408\ : InMux
    port map (
            O => \N__52519\,
            I => \N__52508\
        );

    \I__12407\ : Span4Mux_v
    port map (
            O => \N__52516\,
            I => \N__52503\
        );

    \I__12406\ : LocalMux
    port map (
            O => \N__52513\,
            I => \N__52503\
        );

    \I__12405\ : InMux
    port map (
            O => \N__52512\,
            I => \N__52500\
        );

    \I__12404\ : InMux
    port map (
            O => \N__52511\,
            I => \N__52497\
        );

    \I__12403\ : LocalMux
    port map (
            O => \N__52508\,
            I => \sCounterDACZ0Z_1\
        );

    \I__12402\ : Odrv4
    port map (
            O => \N__52503\,
            I => \sCounterDACZ0Z_1\
        );

    \I__12401\ : LocalMux
    port map (
            O => \N__52500\,
            I => \sCounterDACZ0Z_1\
        );

    \I__12400\ : LocalMux
    port map (
            O => \N__52497\,
            I => \sCounterDACZ0Z_1\
        );

    \I__12399\ : InMux
    port map (
            O => \N__52488\,
            I => \N__52484\
        );

    \I__12398\ : InMux
    port map (
            O => \N__52487\,
            I => \N__52481\
        );

    \I__12397\ : LocalMux
    port map (
            O => \N__52484\,
            I => \sCounterDACZ0Z_7\
        );

    \I__12396\ : LocalMux
    port map (
            O => \N__52481\,
            I => \sCounterDACZ0Z_7\
        );

    \I__12395\ : InMux
    port map (
            O => \N__52476\,
            I => \N__52472\
        );

    \I__12394\ : InMux
    port map (
            O => \N__52475\,
            I => \N__52469\
        );

    \I__12393\ : LocalMux
    port map (
            O => \N__52472\,
            I => \sCounterDACZ0Z_2\
        );

    \I__12392\ : LocalMux
    port map (
            O => \N__52469\,
            I => \sCounterDACZ0Z_2\
        );

    \I__12391\ : CascadeMux
    port map (
            O => \N__52464\,
            I => \N__52460\
        );

    \I__12390\ : InMux
    port map (
            O => \N__52463\,
            I => \N__52457\
        );

    \I__12389\ : InMux
    port map (
            O => \N__52460\,
            I => \N__52454\
        );

    \I__12388\ : LocalMux
    port map (
            O => \N__52457\,
            I => \sCounterDACZ0Z_9\
        );

    \I__12387\ : LocalMux
    port map (
            O => \N__52454\,
            I => \sCounterDACZ0Z_9\
        );

    \I__12386\ : CascadeMux
    port map (
            O => \N__52449\,
            I => \N__52446\
        );

    \I__12385\ : InMux
    port map (
            O => \N__52446\,
            I => \N__52441\
        );

    \I__12384\ : InMux
    port map (
            O => \N__52445\,
            I => \N__52438\
        );

    \I__12383\ : InMux
    port map (
            O => \N__52444\,
            I => \N__52435\
        );

    \I__12382\ : LocalMux
    port map (
            O => \N__52441\,
            I => \N__52430\
        );

    \I__12381\ : LocalMux
    port map (
            O => \N__52438\,
            I => \N__52430\
        );

    \I__12380\ : LocalMux
    port map (
            O => \N__52435\,
            I => \sCounterDACZ0Z_6\
        );

    \I__12379\ : Odrv12
    port map (
            O => \N__52430\,
            I => \sCounterDACZ0Z_6\
        );

    \I__12378\ : InMux
    port map (
            O => \N__52425\,
            I => \N__52422\
        );

    \I__12377\ : LocalMux
    port map (
            O => \N__52422\,
            I => \N__52416\
        );

    \I__12376\ : InMux
    port map (
            O => \N__52421\,
            I => \N__52407\
        );

    \I__12375\ : InMux
    port map (
            O => \N__52420\,
            I => \N__52407\
        );

    \I__12374\ : InMux
    port map (
            O => \N__52419\,
            I => \N__52407\
        );

    \I__12373\ : Span4Mux_h
    port map (
            O => \N__52416\,
            I => \N__52404\
        );

    \I__12372\ : InMux
    port map (
            O => \N__52415\,
            I => \N__52401\
        );

    \I__12371\ : InMux
    port map (
            O => \N__52414\,
            I => \N__52398\
        );

    \I__12370\ : LocalMux
    port map (
            O => \N__52407\,
            I => \N__52395\
        );

    \I__12369\ : Sp12to4
    port map (
            O => \N__52404\,
            I => \N__52390\
        );

    \I__12368\ : LocalMux
    port map (
            O => \N__52401\,
            I => \N__52390\
        );

    \I__12367\ : LocalMux
    port map (
            O => \N__52398\,
            I => \N__52387\
        );

    \I__12366\ : Span12Mux_v
    port map (
            O => \N__52395\,
            I => \N__52384\
        );

    \I__12365\ : Span12Mux_v
    port map (
            O => \N__52390\,
            I => \N__52381\
        );

    \I__12364\ : Span4Mux_v
    port map (
            O => \N__52387\,
            I => \N__52378\
        );

    \I__12363\ : Span12Mux_h
    port map (
            O => \N__52384\,
            I => \N__52375\
        );

    \I__12362\ : Span12Mux_h
    port map (
            O => \N__52381\,
            I => \N__52372\
        );

    \I__12361\ : Span4Mux_v
    port map (
            O => \N__52378\,
            I => \N__52369\
        );

    \I__12360\ : Odrv12
    port map (
            O => \N__52375\,
            I => spi_cs_rpi_c
        );

    \I__12359\ : Odrv12
    port map (
            O => \N__52372\,
            I => spi_cs_rpi_c
        );

    \I__12358\ : Odrv4
    port map (
            O => \N__52369\,
            I => spi_cs_rpi_c
        );

    \I__12357\ : IoInMux
    port map (
            O => \N__52362\,
            I => \N__52359\
        );

    \I__12356\ : LocalMux
    port map (
            O => \N__52359\,
            I => \N__52356\
        );

    \I__12355\ : Span4Mux_s2_v
    port map (
            O => \N__52356\,
            I => \N__52353\
        );

    \I__12354\ : Span4Mux_v
    port map (
            O => \N__52353\,
            I => \N__52350\
        );

    \I__12353\ : Odrv4
    port map (
            O => \N__52350\,
            I => spi_cs_flash_c
        );

    \I__12352\ : InMux
    port map (
            O => \N__52347\,
            I => \N__52344\
        );

    \I__12351\ : LocalMux
    port map (
            O => \N__52344\,
            I => \N__52340\
        );

    \I__12350\ : InMux
    port map (
            O => \N__52343\,
            I => \N__52337\
        );

    \I__12349\ : Span4Mux_v
    port map (
            O => \N__52340\,
            I => \N__52334\
        );

    \I__12348\ : LocalMux
    port map (
            O => \N__52337\,
            I => \N__52331\
        );

    \I__12347\ : Sp12to4
    port map (
            O => \N__52334\,
            I => \N__52328\
        );

    \I__12346\ : Span4Mux_v
    port map (
            O => \N__52331\,
            I => \N__52325\
        );

    \I__12345\ : Span12Mux_h
    port map (
            O => \N__52328\,
            I => \N__52320\
        );

    \I__12344\ : Sp12to4
    port map (
            O => \N__52325\,
            I => \N__52320\
        );

    \I__12343\ : Span12Mux_h
    port map (
            O => \N__52320\,
            I => \N__52317\
        );

    \I__12342\ : Odrv12
    port map (
            O => \N__52317\,
            I => spi_sclk_rpi_c
        );

    \I__12341\ : InMux
    port map (
            O => \N__52314\,
            I => \N__52311\
        );

    \I__12340\ : LocalMux
    port map (
            O => \N__52311\,
            I => \N__52308\
        );

    \I__12339\ : Span4Mux_h
    port map (
            O => \N__52308\,
            I => \N__52305\
        );

    \I__12338\ : Span4Mux_h
    port map (
            O => \N__52305\,
            I => \N__52301\
        );

    \I__12337\ : InMux
    port map (
            O => \N__52304\,
            I => \N__52298\
        );

    \I__12336\ : Span4Mux_h
    port map (
            O => \N__52301\,
            I => \N__52291\
        );

    \I__12335\ : LocalMux
    port map (
            O => \N__52298\,
            I => \N__52291\
        );

    \I__12334\ : InMux
    port map (
            O => \N__52297\,
            I => \N__52288\
        );

    \I__12333\ : InMux
    port map (
            O => \N__52296\,
            I => \N__52285\
        );

    \I__12332\ : Sp12to4
    port map (
            O => \N__52291\,
            I => \N__52278\
        );

    \I__12331\ : LocalMux
    port map (
            O => \N__52288\,
            I => \N__52278\
        );

    \I__12330\ : LocalMux
    port map (
            O => \N__52285\,
            I => \N__52278\
        );

    \I__12329\ : Span12Mux_v
    port map (
            O => \N__52278\,
            I => \N__52275\
        );

    \I__12328\ : Odrv12
    port map (
            O => \N__52275\,
            I => cs_rpi2flash_c
        );

    \I__12327\ : IoInMux
    port map (
            O => \N__52272\,
            I => \N__52269\
        );

    \I__12326\ : LocalMux
    port map (
            O => \N__52269\,
            I => \N__52266\
        );

    \I__12325\ : Span12Mux_s6_v
    port map (
            O => \N__52266\,
            I => \N__52263\
        );

    \I__12324\ : Odrv12
    port map (
            O => \N__52263\,
            I => spi_sclk_flash_c
        );

    \I__12323\ : CascadeMux
    port map (
            O => \N__52260\,
            I => \N__52257\
        );

    \I__12322\ : InMux
    port map (
            O => \N__52257\,
            I => \N__52254\
        );

    \I__12321\ : LocalMux
    port map (
            O => \N__52254\,
            I => \N__52250\
        );

    \I__12320\ : CascadeMux
    port map (
            O => \N__52253\,
            I => \N__52247\
        );

    \I__12319\ : Span4Mux_v
    port map (
            O => \N__52250\,
            I => \N__52244\
        );

    \I__12318\ : InMux
    port map (
            O => \N__52247\,
            I => \N__52241\
        );

    \I__12317\ : Odrv4
    port map (
            O => \N__52244\,
            I => \N_14_3\
        );

    \I__12316\ : LocalMux
    port map (
            O => \N__52241\,
            I => \N_14_3\
        );

    \I__12315\ : InMux
    port map (
            O => \N__52236\,
            I => un2_scounterdac_cry_1
        );

    \I__12314\ : InMux
    port map (
            O => \N__52233\,
            I => \N__52229\
        );

    \I__12313\ : InMux
    port map (
            O => \N__52232\,
            I => \N__52226\
        );

    \I__12312\ : LocalMux
    port map (
            O => \N__52229\,
            I => \N__52222\
        );

    \I__12311\ : LocalMux
    port map (
            O => \N__52226\,
            I => \N__52219\
        );

    \I__12310\ : InMux
    port map (
            O => \N__52225\,
            I => \N__52216\
        );

    \I__12309\ : Span4Mux_h
    port map (
            O => \N__52222\,
            I => \N__52213\
        );

    \I__12308\ : Odrv4
    port map (
            O => \N__52219\,
            I => \sCounterDACZ0Z_3\
        );

    \I__12307\ : LocalMux
    port map (
            O => \N__52216\,
            I => \sCounterDACZ0Z_3\
        );

    \I__12306\ : Odrv4
    port map (
            O => \N__52213\,
            I => \sCounterDACZ0Z_3\
        );

    \I__12305\ : InMux
    port map (
            O => \N__52206\,
            I => un2_scounterdac_cry_2
        );

    \I__12304\ : InMux
    port map (
            O => \N__52203\,
            I => un2_scounterdac_cry_3
        );

    \I__12303\ : InMux
    port map (
            O => \N__52200\,
            I => \N__52194\
        );

    \I__12302\ : InMux
    port map (
            O => \N__52199\,
            I => \N__52194\
        );

    \I__12301\ : LocalMux
    port map (
            O => \N__52194\,
            I => \N__52190\
        );

    \I__12300\ : InMux
    port map (
            O => \N__52193\,
            I => \N__52187\
        );

    \I__12299\ : Span4Mux_v
    port map (
            O => \N__52190\,
            I => \N__52184\
        );

    \I__12298\ : LocalMux
    port map (
            O => \N__52187\,
            I => \sCounterDACZ0Z_5\
        );

    \I__12297\ : Odrv4
    port map (
            O => \N__52184\,
            I => \sCounterDACZ0Z_5\
        );

    \I__12296\ : InMux
    port map (
            O => \N__52179\,
            I => un2_scounterdac_cry_4
        );

    \I__12295\ : InMux
    port map (
            O => \N__52176\,
            I => \N__52173\
        );

    \I__12294\ : LocalMux
    port map (
            O => \N__52173\,
            I => \N__52170\
        );

    \I__12293\ : Odrv4
    port map (
            O => \N__52170\,
            I => \un2_scounterdac_cry_5_THRU_CO\
        );

    \I__12292\ : InMux
    port map (
            O => \N__52167\,
            I => un2_scounterdac_cry_5
        );

    \I__12291\ : InMux
    port map (
            O => \N__52164\,
            I => un2_scounterdac_cry_6
        );

    \I__12290\ : InMux
    port map (
            O => \N__52161\,
            I => \N__52132\
        );

    \I__12289\ : InMux
    port map (
            O => \N__52160\,
            I => \N__52132\
        );

    \I__12288\ : InMux
    port map (
            O => \N__52159\,
            I => \N__52123\
        );

    \I__12287\ : InMux
    port map (
            O => \N__52158\,
            I => \N__52123\
        );

    \I__12286\ : InMux
    port map (
            O => \N__52157\,
            I => \N__52123\
        );

    \I__12285\ : InMux
    port map (
            O => \N__52156\,
            I => \N__52123\
        );

    \I__12284\ : InMux
    port map (
            O => \N__52155\,
            I => \N__52099\
        );

    \I__12283\ : InMux
    port map (
            O => \N__52154\,
            I => \N__52099\
        );

    \I__12282\ : InMux
    port map (
            O => \N__52153\,
            I => \N__52096\
        );

    \I__12281\ : InMux
    port map (
            O => \N__52152\,
            I => \N__52084\
        );

    \I__12280\ : InMux
    port map (
            O => \N__52151\,
            I => \N__52084\
        );

    \I__12279\ : InMux
    port map (
            O => \N__52150\,
            I => \N__52084\
        );

    \I__12278\ : InMux
    port map (
            O => \N__52149\,
            I => \N__52068\
        );

    \I__12277\ : InMux
    port map (
            O => \N__52148\,
            I => \N__52068\
        );

    \I__12276\ : InMux
    port map (
            O => \N__52147\,
            I => \N__52059\
        );

    \I__12275\ : InMux
    port map (
            O => \N__52146\,
            I => \N__52059\
        );

    \I__12274\ : InMux
    port map (
            O => \N__52145\,
            I => \N__52054\
        );

    \I__12273\ : InMux
    port map (
            O => \N__52144\,
            I => \N__52054\
        );

    \I__12272\ : InMux
    port map (
            O => \N__52143\,
            I => \N__52047\
        );

    \I__12271\ : InMux
    port map (
            O => \N__52142\,
            I => \N__52047\
        );

    \I__12270\ : InMux
    port map (
            O => \N__52141\,
            I => \N__52047\
        );

    \I__12269\ : InMux
    port map (
            O => \N__52140\,
            I => \N__52042\
        );

    \I__12268\ : InMux
    port map (
            O => \N__52139\,
            I => \N__52042\
        );

    \I__12267\ : InMux
    port map (
            O => \N__52138\,
            I => \N__52036\
        );

    \I__12266\ : InMux
    port map (
            O => \N__52137\,
            I => \N__52036\
        );

    \I__12265\ : LocalMux
    port map (
            O => \N__52132\,
            I => \N__52031\
        );

    \I__12264\ : LocalMux
    port map (
            O => \N__52123\,
            I => \N__52031\
        );

    \I__12263\ : InMux
    port map (
            O => \N__52122\,
            I => \N__52028\
        );

    \I__12262\ : InMux
    port map (
            O => \N__52121\,
            I => \N__52023\
        );

    \I__12261\ : InMux
    port map (
            O => \N__52120\,
            I => \N__52023\
        );

    \I__12260\ : InMux
    port map (
            O => \N__52119\,
            I => \N__52020\
        );

    \I__12259\ : CascadeMux
    port map (
            O => \N__52118\,
            I => \N__52009\
        );

    \I__12258\ : InMux
    port map (
            O => \N__52117\,
            I => \N__51986\
        );

    \I__12257\ : InMux
    port map (
            O => \N__52116\,
            I => \N__51986\
        );

    \I__12256\ : InMux
    port map (
            O => \N__52115\,
            I => \N__51986\
        );

    \I__12255\ : InMux
    port map (
            O => \N__52114\,
            I => \N__51980\
        );

    \I__12254\ : InMux
    port map (
            O => \N__52113\,
            I => \N__51975\
        );

    \I__12253\ : InMux
    port map (
            O => \N__52112\,
            I => \N__51975\
        );

    \I__12252\ : InMux
    port map (
            O => \N__52111\,
            I => \N__51963\
        );

    \I__12251\ : InMux
    port map (
            O => \N__52110\,
            I => \N__51963\
        );

    \I__12250\ : InMux
    port map (
            O => \N__52109\,
            I => \N__51963\
        );

    \I__12249\ : InMux
    port map (
            O => \N__52108\,
            I => \N__51958\
        );

    \I__12248\ : InMux
    port map (
            O => \N__52107\,
            I => \N__51958\
        );

    \I__12247\ : InMux
    port map (
            O => \N__52106\,
            I => \N__51951\
        );

    \I__12246\ : InMux
    port map (
            O => \N__52105\,
            I => \N__51951\
        );

    \I__12245\ : InMux
    port map (
            O => \N__52104\,
            I => \N__51951\
        );

    \I__12244\ : LocalMux
    port map (
            O => \N__52099\,
            I => \N__51948\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__52096\,
            I => \N__51945\
        );

    \I__12242\ : InMux
    port map (
            O => \N__52095\,
            I => \N__51934\
        );

    \I__12241\ : InMux
    port map (
            O => \N__52094\,
            I => \N__51934\
        );

    \I__12240\ : InMux
    port map (
            O => \N__52093\,
            I => \N__51934\
        );

    \I__12239\ : InMux
    port map (
            O => \N__52092\,
            I => \N__51934\
        );

    \I__12238\ : InMux
    port map (
            O => \N__52091\,
            I => \N__51934\
        );

    \I__12237\ : LocalMux
    port map (
            O => \N__52084\,
            I => \N__51931\
        );

    \I__12236\ : InMux
    port map (
            O => \N__52083\,
            I => \N__51924\
        );

    \I__12235\ : InMux
    port map (
            O => \N__52082\,
            I => \N__51924\
        );

    \I__12234\ : InMux
    port map (
            O => \N__52081\,
            I => \N__51924\
        );

    \I__12233\ : InMux
    port map (
            O => \N__52080\,
            I => \N__51917\
        );

    \I__12232\ : InMux
    port map (
            O => \N__52079\,
            I => \N__51917\
        );

    \I__12231\ : InMux
    port map (
            O => \N__52078\,
            I => \N__51917\
        );

    \I__12230\ : InMux
    port map (
            O => \N__52077\,
            I => \N__51914\
        );

    \I__12229\ : InMux
    port map (
            O => \N__52076\,
            I => \N__51911\
        );

    \I__12228\ : InMux
    port map (
            O => \N__52075\,
            I => \N__51897\
        );

    \I__12227\ : InMux
    port map (
            O => \N__52074\,
            I => \N__51897\
        );

    \I__12226\ : InMux
    port map (
            O => \N__52073\,
            I => \N__51882\
        );

    \I__12225\ : LocalMux
    port map (
            O => \N__52068\,
            I => \N__51875\
        );

    \I__12224\ : InMux
    port map (
            O => \N__52067\,
            I => \N__51868\
        );

    \I__12223\ : InMux
    port map (
            O => \N__52066\,
            I => \N__51868\
        );

    \I__12222\ : InMux
    port map (
            O => \N__52065\,
            I => \N__51868\
        );

    \I__12221\ : InMux
    port map (
            O => \N__52064\,
            I => \N__51861\
        );

    \I__12220\ : LocalMux
    port map (
            O => \N__52059\,
            I => \N__51858\
        );

    \I__12219\ : LocalMux
    port map (
            O => \N__52054\,
            I => \N__51851\
        );

    \I__12218\ : LocalMux
    port map (
            O => \N__52047\,
            I => \N__51851\
        );

    \I__12217\ : LocalMux
    port map (
            O => \N__52042\,
            I => \N__51851\
        );

    \I__12216\ : InMux
    port map (
            O => \N__52041\,
            I => \N__51848\
        );

    \I__12215\ : LocalMux
    port map (
            O => \N__52036\,
            I => \N__51843\
        );

    \I__12214\ : Span4Mux_h
    port map (
            O => \N__52031\,
            I => \N__51843\
        );

    \I__12213\ : LocalMux
    port map (
            O => \N__52028\,
            I => \N__51836\
        );

    \I__12212\ : LocalMux
    port map (
            O => \N__52023\,
            I => \N__51836\
        );

    \I__12211\ : LocalMux
    port map (
            O => \N__52020\,
            I => \N__51836\
        );

    \I__12210\ : InMux
    port map (
            O => \N__52019\,
            I => \N__51831\
        );

    \I__12209\ : InMux
    port map (
            O => \N__52018\,
            I => \N__51831\
        );

    \I__12208\ : InMux
    port map (
            O => \N__52017\,
            I => \N__51826\
        );

    \I__12207\ : InMux
    port map (
            O => \N__52016\,
            I => \N__51826\
        );

    \I__12206\ : InMux
    port map (
            O => \N__52015\,
            I => \N__51819\
        );

    \I__12205\ : InMux
    port map (
            O => \N__52014\,
            I => \N__51819\
        );

    \I__12204\ : InMux
    port map (
            O => \N__52013\,
            I => \N__51819\
        );

    \I__12203\ : CascadeMux
    port map (
            O => \N__52012\,
            I => \N__51805\
        );

    \I__12202\ : InMux
    port map (
            O => \N__52009\,
            I => \N__51794\
        );

    \I__12201\ : InMux
    port map (
            O => \N__52008\,
            I => \N__51794\
        );

    \I__12200\ : InMux
    port map (
            O => \N__52007\,
            I => \N__51794\
        );

    \I__12199\ : InMux
    port map (
            O => \N__52006\,
            I => \N__51785\
        );

    \I__12198\ : InMux
    port map (
            O => \N__52005\,
            I => \N__51785\
        );

    \I__12197\ : InMux
    port map (
            O => \N__52004\,
            I => \N__51785\
        );

    \I__12196\ : InMux
    port map (
            O => \N__52003\,
            I => \N__51785\
        );

    \I__12195\ : InMux
    port map (
            O => \N__52002\,
            I => \N__51778\
        );

    \I__12194\ : InMux
    port map (
            O => \N__52001\,
            I => \N__51778\
        );

    \I__12193\ : InMux
    port map (
            O => \N__52000\,
            I => \N__51778\
        );

    \I__12192\ : InMux
    port map (
            O => \N__51999\,
            I => \N__51773\
        );

    \I__12191\ : InMux
    port map (
            O => \N__51998\,
            I => \N__51773\
        );

    \I__12190\ : InMux
    port map (
            O => \N__51997\,
            I => \N__51763\
        );

    \I__12189\ : InMux
    port map (
            O => \N__51996\,
            I => \N__51763\
        );

    \I__12188\ : InMux
    port map (
            O => \N__51995\,
            I => \N__51763\
        );

    \I__12187\ : InMux
    port map (
            O => \N__51994\,
            I => \N__51758\
        );

    \I__12186\ : InMux
    port map (
            O => \N__51993\,
            I => \N__51758\
        );

    \I__12185\ : LocalMux
    port map (
            O => \N__51986\,
            I => \N__51755\
        );

    \I__12184\ : InMux
    port map (
            O => \N__51985\,
            I => \N__51752\
        );

    \I__12183\ : InMux
    port map (
            O => \N__51984\,
            I => \N__51747\
        );

    \I__12182\ : InMux
    port map (
            O => \N__51983\,
            I => \N__51747\
        );

    \I__12181\ : LocalMux
    port map (
            O => \N__51980\,
            I => \N__51742\
        );

    \I__12180\ : LocalMux
    port map (
            O => \N__51975\,
            I => \N__51742\
        );

    \I__12179\ : InMux
    port map (
            O => \N__51974\,
            I => \N__51737\
        );

    \I__12178\ : InMux
    port map (
            O => \N__51973\,
            I => \N__51737\
        );

    \I__12177\ : InMux
    port map (
            O => \N__51972\,
            I => \N__51730\
        );

    \I__12176\ : InMux
    port map (
            O => \N__51971\,
            I => \N__51730\
        );

    \I__12175\ : InMux
    port map (
            O => \N__51970\,
            I => \N__51730\
        );

    \I__12174\ : LocalMux
    port map (
            O => \N__51963\,
            I => \N__51727\
        );

    \I__12173\ : LocalMux
    port map (
            O => \N__51958\,
            I => \N__51722\
        );

    \I__12172\ : LocalMux
    port map (
            O => \N__51951\,
            I => \N__51722\
        );

    \I__12171\ : Span4Mux_h
    port map (
            O => \N__51948\,
            I => \N__51711\
        );

    \I__12170\ : Span4Mux_v
    port map (
            O => \N__51945\,
            I => \N__51711\
        );

    \I__12169\ : LocalMux
    port map (
            O => \N__51934\,
            I => \N__51711\
        );

    \I__12168\ : Span4Mux_v
    port map (
            O => \N__51931\,
            I => \N__51711\
        );

    \I__12167\ : LocalMux
    port map (
            O => \N__51924\,
            I => \N__51711\
        );

    \I__12166\ : LocalMux
    port map (
            O => \N__51917\,
            I => \N__51704\
        );

    \I__12165\ : LocalMux
    port map (
            O => \N__51914\,
            I => \N__51704\
        );

    \I__12164\ : LocalMux
    port map (
            O => \N__51911\,
            I => \N__51704\
        );

    \I__12163\ : InMux
    port map (
            O => \N__51910\,
            I => \N__51695\
        );

    \I__12162\ : InMux
    port map (
            O => \N__51909\,
            I => \N__51695\
        );

    \I__12161\ : InMux
    port map (
            O => \N__51908\,
            I => \N__51695\
        );

    \I__12160\ : InMux
    port map (
            O => \N__51907\,
            I => \N__51695\
        );

    \I__12159\ : InMux
    port map (
            O => \N__51906\,
            I => \N__51684\
        );

    \I__12158\ : InMux
    port map (
            O => \N__51905\,
            I => \N__51684\
        );

    \I__12157\ : InMux
    port map (
            O => \N__51904\,
            I => \N__51684\
        );

    \I__12156\ : InMux
    port map (
            O => \N__51903\,
            I => \N__51684\
        );

    \I__12155\ : InMux
    port map (
            O => \N__51902\,
            I => \N__51684\
        );

    \I__12154\ : LocalMux
    port map (
            O => \N__51897\,
            I => \N__51681\
        );

    \I__12153\ : InMux
    port map (
            O => \N__51896\,
            I => \N__51678\
        );

    \I__12152\ : InMux
    port map (
            O => \N__51895\,
            I => \N__51671\
        );

    \I__12151\ : InMux
    port map (
            O => \N__51894\,
            I => \N__51671\
        );

    \I__12150\ : InMux
    port map (
            O => \N__51893\,
            I => \N__51671\
        );

    \I__12149\ : InMux
    port map (
            O => \N__51892\,
            I => \N__51666\
        );

    \I__12148\ : InMux
    port map (
            O => \N__51891\,
            I => \N__51666\
        );

    \I__12147\ : InMux
    port map (
            O => \N__51890\,
            I => \N__51663\
        );

    \I__12146\ : InMux
    port map (
            O => \N__51889\,
            I => \N__51656\
        );

    \I__12145\ : InMux
    port map (
            O => \N__51888\,
            I => \N__51656\
        );

    \I__12144\ : InMux
    port map (
            O => \N__51887\,
            I => \N__51656\
        );

    \I__12143\ : InMux
    port map (
            O => \N__51886\,
            I => \N__51651\
        );

    \I__12142\ : InMux
    port map (
            O => \N__51885\,
            I => \N__51651\
        );

    \I__12141\ : LocalMux
    port map (
            O => \N__51882\,
            I => \N__51648\
        );

    \I__12140\ : InMux
    port map (
            O => \N__51881\,
            I => \N__51645\
        );

    \I__12139\ : InMux
    port map (
            O => \N__51880\,
            I => \N__51638\
        );

    \I__12138\ : InMux
    port map (
            O => \N__51879\,
            I => \N__51638\
        );

    \I__12137\ : InMux
    port map (
            O => \N__51878\,
            I => \N__51638\
        );

    \I__12136\ : Span4Mux_v
    port map (
            O => \N__51875\,
            I => \N__51633\
        );

    \I__12135\ : LocalMux
    port map (
            O => \N__51868\,
            I => \N__51633\
        );

    \I__12134\ : InMux
    port map (
            O => \N__51867\,
            I => \N__51624\
        );

    \I__12133\ : InMux
    port map (
            O => \N__51866\,
            I => \N__51624\
        );

    \I__12132\ : InMux
    port map (
            O => \N__51865\,
            I => \N__51624\
        );

    \I__12131\ : InMux
    port map (
            O => \N__51864\,
            I => \N__51624\
        );

    \I__12130\ : LocalMux
    port map (
            O => \N__51861\,
            I => \N__51617\
        );

    \I__12129\ : Span4Mux_v
    port map (
            O => \N__51858\,
            I => \N__51617\
        );

    \I__12128\ : Span4Mux_v
    port map (
            O => \N__51851\,
            I => \N__51617\
        );

    \I__12127\ : LocalMux
    port map (
            O => \N__51848\,
            I => \N__51610\
        );

    \I__12126\ : Span4Mux_v
    port map (
            O => \N__51843\,
            I => \N__51610\
        );

    \I__12125\ : Span4Mux_h
    port map (
            O => \N__51836\,
            I => \N__51610\
        );

    \I__12124\ : LocalMux
    port map (
            O => \N__51831\,
            I => \N__51603\
        );

    \I__12123\ : LocalMux
    port map (
            O => \N__51826\,
            I => \N__51603\
        );

    \I__12122\ : LocalMux
    port map (
            O => \N__51819\,
            I => \N__51603\
        );

    \I__12121\ : InMux
    port map (
            O => \N__51818\,
            I => \N__51589\
        );

    \I__12120\ : InMux
    port map (
            O => \N__51817\,
            I => \N__51589\
        );

    \I__12119\ : InMux
    port map (
            O => \N__51816\,
            I => \N__51582\
        );

    \I__12118\ : InMux
    port map (
            O => \N__51815\,
            I => \N__51582\
        );

    \I__12117\ : InMux
    port map (
            O => \N__51814\,
            I => \N__51582\
        );

    \I__12116\ : InMux
    port map (
            O => \N__51813\,
            I => \N__51577\
        );

    \I__12115\ : InMux
    port map (
            O => \N__51812\,
            I => \N__51577\
        );

    \I__12114\ : InMux
    port map (
            O => \N__51811\,
            I => \N__51570\
        );

    \I__12113\ : InMux
    port map (
            O => \N__51810\,
            I => \N__51570\
        );

    \I__12112\ : InMux
    port map (
            O => \N__51809\,
            I => \N__51570\
        );

    \I__12111\ : InMux
    port map (
            O => \N__51808\,
            I => \N__51565\
        );

    \I__12110\ : InMux
    port map (
            O => \N__51805\,
            I => \N__51565\
        );

    \I__12109\ : InMux
    port map (
            O => \N__51804\,
            I => \N__51556\
        );

    \I__12108\ : InMux
    port map (
            O => \N__51803\,
            I => \N__51556\
        );

    \I__12107\ : InMux
    port map (
            O => \N__51802\,
            I => \N__51556\
        );

    \I__12106\ : InMux
    port map (
            O => \N__51801\,
            I => \N__51556\
        );

    \I__12105\ : LocalMux
    port map (
            O => \N__51794\,
            I => \N__51542\
        );

    \I__12104\ : LocalMux
    port map (
            O => \N__51785\,
            I => \N__51542\
        );

    \I__12103\ : LocalMux
    port map (
            O => \N__51778\,
            I => \N__51542\
        );

    \I__12102\ : LocalMux
    port map (
            O => \N__51773\,
            I => \N__51542\
        );

    \I__12101\ : InMux
    port map (
            O => \N__51772\,
            I => \N__51530\
        );

    \I__12100\ : InMux
    port map (
            O => \N__51771\,
            I => \N__51530\
        );

    \I__12099\ : InMux
    port map (
            O => \N__51770\,
            I => \N__51530\
        );

    \I__12098\ : LocalMux
    port map (
            O => \N__51763\,
            I => \N__51521\
        );

    \I__12097\ : LocalMux
    port map (
            O => \N__51758\,
            I => \N__51521\
        );

    \I__12096\ : Span4Mux_v
    port map (
            O => \N__51755\,
            I => \N__51521\
        );

    \I__12095\ : LocalMux
    port map (
            O => \N__51752\,
            I => \N__51521\
        );

    \I__12094\ : LocalMux
    port map (
            O => \N__51747\,
            I => \N__51514\
        );

    \I__12093\ : Span4Mux_h
    port map (
            O => \N__51742\,
            I => \N__51514\
        );

    \I__12092\ : LocalMux
    port map (
            O => \N__51737\,
            I => \N__51514\
        );

    \I__12091\ : LocalMux
    port map (
            O => \N__51730\,
            I => \N__51503\
        );

    \I__12090\ : Span4Mux_v
    port map (
            O => \N__51727\,
            I => \N__51503\
        );

    \I__12089\ : Span4Mux_v
    port map (
            O => \N__51722\,
            I => \N__51503\
        );

    \I__12088\ : Span4Mux_h
    port map (
            O => \N__51711\,
            I => \N__51503\
        );

    \I__12087\ : Span4Mux_h
    port map (
            O => \N__51704\,
            I => \N__51503\
        );

    \I__12086\ : LocalMux
    port map (
            O => \N__51695\,
            I => \N__51496\
        );

    \I__12085\ : LocalMux
    port map (
            O => \N__51684\,
            I => \N__51496\
        );

    \I__12084\ : Span4Mux_h
    port map (
            O => \N__51681\,
            I => \N__51490\
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__51678\,
            I => \N__51481\
        );

    \I__12082\ : LocalMux
    port map (
            O => \N__51671\,
            I => \N__51481\
        );

    \I__12081\ : LocalMux
    port map (
            O => \N__51666\,
            I => \N__51481\
        );

    \I__12080\ : LocalMux
    port map (
            O => \N__51663\,
            I => \N__51481\
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__51656\,
            I => \N__51472\
        );

    \I__12078\ : LocalMux
    port map (
            O => \N__51651\,
            I => \N__51472\
        );

    \I__12077\ : Span4Mux_h
    port map (
            O => \N__51648\,
            I => \N__51461\
        );

    \I__12076\ : LocalMux
    port map (
            O => \N__51645\,
            I => \N__51461\
        );

    \I__12075\ : LocalMux
    port map (
            O => \N__51638\,
            I => \N__51461\
        );

    \I__12074\ : Span4Mux_h
    port map (
            O => \N__51633\,
            I => \N__51461\
        );

    \I__12073\ : LocalMux
    port map (
            O => \N__51624\,
            I => \N__51461\
        );

    \I__12072\ : Span4Mux_h
    port map (
            O => \N__51617\,
            I => \N__51454\
        );

    \I__12071\ : Span4Mux_v
    port map (
            O => \N__51610\,
            I => \N__51454\
        );

    \I__12070\ : Span4Mux_v
    port map (
            O => \N__51603\,
            I => \N__51454\
        );

    \I__12069\ : InMux
    port map (
            O => \N__51602\,
            I => \N__51443\
        );

    \I__12068\ : InMux
    port map (
            O => \N__51601\,
            I => \N__51443\
        );

    \I__12067\ : InMux
    port map (
            O => \N__51600\,
            I => \N__51443\
        );

    \I__12066\ : InMux
    port map (
            O => \N__51599\,
            I => \N__51443\
        );

    \I__12065\ : InMux
    port map (
            O => \N__51598\,
            I => \N__51443\
        );

    \I__12064\ : InMux
    port map (
            O => \N__51597\,
            I => \N__51434\
        );

    \I__12063\ : InMux
    port map (
            O => \N__51596\,
            I => \N__51434\
        );

    \I__12062\ : InMux
    port map (
            O => \N__51595\,
            I => \N__51434\
        );

    \I__12061\ : InMux
    port map (
            O => \N__51594\,
            I => \N__51434\
        );

    \I__12060\ : LocalMux
    port map (
            O => \N__51589\,
            I => \N__51421\
        );

    \I__12059\ : LocalMux
    port map (
            O => \N__51582\,
            I => \N__51421\
        );

    \I__12058\ : LocalMux
    port map (
            O => \N__51577\,
            I => \N__51421\
        );

    \I__12057\ : LocalMux
    port map (
            O => \N__51570\,
            I => \N__51421\
        );

    \I__12056\ : LocalMux
    port map (
            O => \N__51565\,
            I => \N__51421\
        );

    \I__12055\ : LocalMux
    port map (
            O => \N__51556\,
            I => \N__51421\
        );

    \I__12054\ : InMux
    port map (
            O => \N__51555\,
            I => \N__51412\
        );

    \I__12053\ : InMux
    port map (
            O => \N__51554\,
            I => \N__51412\
        );

    \I__12052\ : InMux
    port map (
            O => \N__51553\,
            I => \N__51412\
        );

    \I__12051\ : InMux
    port map (
            O => \N__51552\,
            I => \N__51412\
        );

    \I__12050\ : InMux
    port map (
            O => \N__51551\,
            I => \N__51409\
        );

    \I__12049\ : Span12Mux_h
    port map (
            O => \N__51542\,
            I => \N__51406\
        );

    \I__12048\ : InMux
    port map (
            O => \N__51541\,
            I => \N__51395\
        );

    \I__12047\ : InMux
    port map (
            O => \N__51540\,
            I => \N__51395\
        );

    \I__12046\ : InMux
    port map (
            O => \N__51539\,
            I => \N__51395\
        );

    \I__12045\ : InMux
    port map (
            O => \N__51538\,
            I => \N__51395\
        );

    \I__12044\ : InMux
    port map (
            O => \N__51537\,
            I => \N__51395\
        );

    \I__12043\ : LocalMux
    port map (
            O => \N__51530\,
            I => \N__51386\
        );

    \I__12042\ : Span4Mux_v
    port map (
            O => \N__51521\,
            I => \N__51386\
        );

    \I__12041\ : Span4Mux_h
    port map (
            O => \N__51514\,
            I => \N__51386\
        );

    \I__12040\ : Span4Mux_v
    port map (
            O => \N__51503\,
            I => \N__51386\
        );

    \I__12039\ : InMux
    port map (
            O => \N__51502\,
            I => \N__51383\
        );

    \I__12038\ : InMux
    port map (
            O => \N__51501\,
            I => \N__51380\
        );

    \I__12037\ : Span12Mux_v
    port map (
            O => \N__51496\,
            I => \N__51377\
        );

    \I__12036\ : InMux
    port map (
            O => \N__51495\,
            I => \N__51370\
        );

    \I__12035\ : InMux
    port map (
            O => \N__51494\,
            I => \N__51370\
        );

    \I__12034\ : InMux
    port map (
            O => \N__51493\,
            I => \N__51370\
        );

    \I__12033\ : Span4Mux_h
    port map (
            O => \N__51490\,
            I => \N__51365\
        );

    \I__12032\ : Span4Mux_h
    port map (
            O => \N__51481\,
            I => \N__51365\
        );

    \I__12031\ : InMux
    port map (
            O => \N__51480\,
            I => \N__51362\
        );

    \I__12030\ : InMux
    port map (
            O => \N__51479\,
            I => \N__51355\
        );

    \I__12029\ : InMux
    port map (
            O => \N__51478\,
            I => \N__51355\
        );

    \I__12028\ : InMux
    port map (
            O => \N__51477\,
            I => \N__51355\
        );

    \I__12027\ : Span4Mux_h
    port map (
            O => \N__51472\,
            I => \N__51348\
        );

    \I__12026\ : Span4Mux_v
    port map (
            O => \N__51461\,
            I => \N__51348\
        );

    \I__12025\ : Span4Mux_v
    port map (
            O => \N__51454\,
            I => \N__51348\
        );

    \I__12024\ : LocalMux
    port map (
            O => \N__51443\,
            I => \N__51339\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__51434\,
            I => \N__51339\
        );

    \I__12022\ : Span12Mux_h
    port map (
            O => \N__51421\,
            I => \N__51339\
        );

    \I__12021\ : LocalMux
    port map (
            O => \N__51412\,
            I => \N__51339\
        );

    \I__12020\ : LocalMux
    port map (
            O => \N__51409\,
            I => \N__51334\
        );

    \I__12019\ : Span12Mux_v
    port map (
            O => \N__51406\,
            I => \N__51334\
        );

    \I__12018\ : LocalMux
    port map (
            O => \N__51395\,
            I => \N__51329\
        );

    \I__12017\ : Span4Mux_v
    port map (
            O => \N__51386\,
            I => \N__51329\
        );

    \I__12016\ : LocalMux
    port map (
            O => \N__51383\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__12015\ : LocalMux
    port map (
            O => \N__51380\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__12014\ : Odrv12
    port map (
            O => \N__51377\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__12013\ : LocalMux
    port map (
            O => \N__51370\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__12012\ : Odrv4
    port map (
            O => \N__51365\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__12011\ : LocalMux
    port map (
            O => \N__51362\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__12010\ : LocalMux
    port map (
            O => \N__51355\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__12009\ : Odrv4
    port map (
            O => \N__51348\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__12008\ : Odrv12
    port map (
            O => \N__51339\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__12007\ : Odrv12
    port map (
            O => \N__51334\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__12006\ : Odrv4
    port map (
            O => \N__51329\,
            I => \sDAC_mem_pointerZ0Z_0\
        );

    \I__12005\ : InMux
    port map (
            O => \N__51306\,
            I => \N__51303\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__51303\,
            I => \sDAC_mem_15Z0Z_7\
        );

    \I__12003\ : InMux
    port map (
            O => \N__51300\,
            I => \N__51297\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__51297\,
            I => \N__51294\
        );

    \I__12001\ : Span4Mux_h
    port map (
            O => \N__51294\,
            I => \N__51291\
        );

    \I__12000\ : Odrv4
    port map (
            O => \N__51291\,
            I => \sDAC_mem_14Z0Z_7\
        );

    \I__11999\ : InMux
    port map (
            O => \N__51288\,
            I => \N__51285\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__51285\,
            I => \N__51282\
        );

    \I__11997\ : Span4Mux_h
    port map (
            O => \N__51282\,
            I => \N__51279\
        );

    \I__11996\ : Odrv4
    port map (
            O => \N__51279\,
            I => \sDAC_data_RNO_19Z0Z_10\
        );

    \I__11995\ : InMux
    port map (
            O => \N__51276\,
            I => \N__51273\
        );

    \I__11994\ : LocalMux
    port map (
            O => \N__51273\,
            I => \N__51263\
        );

    \I__11993\ : InMux
    port map (
            O => \N__51272\,
            I => \N__51254\
        );

    \I__11992\ : InMux
    port map (
            O => \N__51271\,
            I => \N__51249\
        );

    \I__11991\ : InMux
    port map (
            O => \N__51270\,
            I => \N__51243\
        );

    \I__11990\ : InMux
    port map (
            O => \N__51269\,
            I => \N__51236\
        );

    \I__11989\ : InMux
    port map (
            O => \N__51268\,
            I => \N__51233\
        );

    \I__11988\ : InMux
    port map (
            O => \N__51267\,
            I => \N__51229\
        );

    \I__11987\ : InMux
    port map (
            O => \N__51266\,
            I => \N__51226\
        );

    \I__11986\ : Span4Mux_v
    port map (
            O => \N__51263\,
            I => \N__51223\
        );

    \I__11985\ : InMux
    port map (
            O => \N__51262\,
            I => \N__51220\
        );

    \I__11984\ : InMux
    port map (
            O => \N__51261\,
            I => \N__51217\
        );

    \I__11983\ : InMux
    port map (
            O => \N__51260\,
            I => \N__51213\
        );

    \I__11982\ : InMux
    port map (
            O => \N__51259\,
            I => \N__51210\
        );

    \I__11981\ : InMux
    port map (
            O => \N__51258\,
            I => \N__51207\
        );

    \I__11980\ : InMux
    port map (
            O => \N__51257\,
            I => \N__51204\
        );

    \I__11979\ : LocalMux
    port map (
            O => \N__51254\,
            I => \N__51200\
        );

    \I__11978\ : InMux
    port map (
            O => \N__51253\,
            I => \N__51197\
        );

    \I__11977\ : InMux
    port map (
            O => \N__51252\,
            I => \N__51194\
        );

    \I__11976\ : LocalMux
    port map (
            O => \N__51249\,
            I => \N__51191\
        );

    \I__11975\ : InMux
    port map (
            O => \N__51248\,
            I => \N__51188\
        );

    \I__11974\ : InMux
    port map (
            O => \N__51247\,
            I => \N__51185\
        );

    \I__11973\ : InMux
    port map (
            O => \N__51246\,
            I => \N__51182\
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__51243\,
            I => \N__51178\
        );

    \I__11971\ : InMux
    port map (
            O => \N__51242\,
            I => \N__51175\
        );

    \I__11970\ : InMux
    port map (
            O => \N__51241\,
            I => \N__51172\
        );

    \I__11969\ : InMux
    port map (
            O => \N__51240\,
            I => \N__51169\
        );

    \I__11968\ : InMux
    port map (
            O => \N__51239\,
            I => \N__51165\
        );

    \I__11967\ : LocalMux
    port map (
            O => \N__51236\,
            I => \N__51159\
        );

    \I__11966\ : LocalMux
    port map (
            O => \N__51233\,
            I => \N__51159\
        );

    \I__11965\ : InMux
    port map (
            O => \N__51232\,
            I => \N__51152\
        );

    \I__11964\ : LocalMux
    port map (
            O => \N__51229\,
            I => \N__51147\
        );

    \I__11963\ : LocalMux
    port map (
            O => \N__51226\,
            I => \N__51147\
        );

    \I__11962\ : Span4Mux_v
    port map (
            O => \N__51223\,
            I => \N__51140\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__51220\,
            I => \N__51140\
        );

    \I__11960\ : LocalMux
    port map (
            O => \N__51217\,
            I => \N__51140\
        );

    \I__11959\ : InMux
    port map (
            O => \N__51216\,
            I => \N__51135\
        );

    \I__11958\ : LocalMux
    port map (
            O => \N__51213\,
            I => \N__51127\
        );

    \I__11957\ : LocalMux
    port map (
            O => \N__51210\,
            I => \N__51127\
        );

    \I__11956\ : LocalMux
    port map (
            O => \N__51207\,
            I => \N__51122\
        );

    \I__11955\ : LocalMux
    port map (
            O => \N__51204\,
            I => \N__51122\
        );

    \I__11954\ : InMux
    port map (
            O => \N__51203\,
            I => \N__51119\
        );

    \I__11953\ : Span4Mux_h
    port map (
            O => \N__51200\,
            I => \N__51112\
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__51197\,
            I => \N__51112\
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__51194\,
            I => \N__51112\
        );

    \I__11950\ : Span4Mux_v
    port map (
            O => \N__51191\,
            I => \N__51105\
        );

    \I__11949\ : LocalMux
    port map (
            O => \N__51188\,
            I => \N__51105\
        );

    \I__11948\ : LocalMux
    port map (
            O => \N__51185\,
            I => \N__51105\
        );

    \I__11947\ : LocalMux
    port map (
            O => \N__51182\,
            I => \N__51102\
        );

    \I__11946\ : InMux
    port map (
            O => \N__51181\,
            I => \N__51096\
        );

    \I__11945\ : Span4Mux_v
    port map (
            O => \N__51178\,
            I => \N__51087\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__51175\,
            I => \N__51087\
        );

    \I__11943\ : LocalMux
    port map (
            O => \N__51172\,
            I => \N__51087\
        );

    \I__11942\ : LocalMux
    port map (
            O => \N__51169\,
            I => \N__51087\
        );

    \I__11941\ : InMux
    port map (
            O => \N__51168\,
            I => \N__51084\
        );

    \I__11940\ : LocalMux
    port map (
            O => \N__51165\,
            I => \N__51075\
        );

    \I__11939\ : InMux
    port map (
            O => \N__51164\,
            I => \N__51072\
        );

    \I__11938\ : Span4Mux_v
    port map (
            O => \N__51159\,
            I => \N__51069\
        );

    \I__11937\ : InMux
    port map (
            O => \N__51158\,
            I => \N__51066\
        );

    \I__11936\ : InMux
    port map (
            O => \N__51157\,
            I => \N__51063\
        );

    \I__11935\ : InMux
    port map (
            O => \N__51156\,
            I => \N__51060\
        );

    \I__11934\ : InMux
    port map (
            O => \N__51155\,
            I => \N__51057\
        );

    \I__11933\ : LocalMux
    port map (
            O => \N__51152\,
            I => \N__51054\
        );

    \I__11932\ : Span4Mux_v
    port map (
            O => \N__51147\,
            I => \N__51051\
        );

    \I__11931\ : Span4Mux_v
    port map (
            O => \N__51140\,
            I => \N__51048\
        );

    \I__11930\ : InMux
    port map (
            O => \N__51139\,
            I => \N__51045\
        );

    \I__11929\ : InMux
    port map (
            O => \N__51138\,
            I => \N__51042\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__51135\,
            I => \N__51037\
        );

    \I__11927\ : InMux
    port map (
            O => \N__51134\,
            I => \N__51034\
        );

    \I__11926\ : InMux
    port map (
            O => \N__51133\,
            I => \N__51031\
        );

    \I__11925\ : InMux
    port map (
            O => \N__51132\,
            I => \N__51028\
        );

    \I__11924\ : Span4Mux_v
    port map (
            O => \N__51127\,
            I => \N__51017\
        );

    \I__11923\ : Span4Mux_h
    port map (
            O => \N__51122\,
            I => \N__51017\
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__51119\,
            I => \N__51017\
        );

    \I__11921\ : Span4Mux_v
    port map (
            O => \N__51112\,
            I => \N__51010\
        );

    \I__11920\ : Span4Mux_v
    port map (
            O => \N__51105\,
            I => \N__51010\
        );

    \I__11919\ : Span4Mux_h
    port map (
            O => \N__51102\,
            I => \N__51010\
        );

    \I__11918\ : InMux
    port map (
            O => \N__51101\,
            I => \N__51007\
        );

    \I__11917\ : InMux
    port map (
            O => \N__51100\,
            I => \N__51004\
        );

    \I__11916\ : InMux
    port map (
            O => \N__51099\,
            I => \N__51001\
        );

    \I__11915\ : LocalMux
    port map (
            O => \N__51096\,
            I => \N__50994\
        );

    \I__11914\ : Span4Mux_v
    port map (
            O => \N__51087\,
            I => \N__50994\
        );

    \I__11913\ : LocalMux
    port map (
            O => \N__51084\,
            I => \N__50994\
        );

    \I__11912\ : InMux
    port map (
            O => \N__51083\,
            I => \N__50991\
        );

    \I__11911\ : InMux
    port map (
            O => \N__51082\,
            I => \N__50988\
        );

    \I__11910\ : InMux
    port map (
            O => \N__51081\,
            I => \N__50983\
        );

    \I__11909\ : InMux
    port map (
            O => \N__51080\,
            I => \N__50978\
        );

    \I__11908\ : InMux
    port map (
            O => \N__51079\,
            I => \N__50975\
        );

    \I__11907\ : InMux
    port map (
            O => \N__51078\,
            I => \N__50972\
        );

    \I__11906\ : Span4Mux_h
    port map (
            O => \N__51075\,
            I => \N__50967\
        );

    \I__11905\ : LocalMux
    port map (
            O => \N__51072\,
            I => \N__50967\
        );

    \I__11904\ : Span4Mux_v
    port map (
            O => \N__51069\,
            I => \N__50956\
        );

    \I__11903\ : LocalMux
    port map (
            O => \N__51066\,
            I => \N__50956\
        );

    \I__11902\ : LocalMux
    port map (
            O => \N__51063\,
            I => \N__50956\
        );

    \I__11901\ : LocalMux
    port map (
            O => \N__51060\,
            I => \N__50956\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__51057\,
            I => \N__50956\
        );

    \I__11899\ : Span4Mux_v
    port map (
            O => \N__51054\,
            I => \N__50953\
        );

    \I__11898\ : Span4Mux_v
    port map (
            O => \N__51051\,
            I => \N__50944\
        );

    \I__11897\ : Span4Mux_h
    port map (
            O => \N__51048\,
            I => \N__50944\
        );

    \I__11896\ : LocalMux
    port map (
            O => \N__51045\,
            I => \N__50944\
        );

    \I__11895\ : LocalMux
    port map (
            O => \N__51042\,
            I => \N__50944\
        );

    \I__11894\ : InMux
    port map (
            O => \N__51041\,
            I => \N__50941\
        );

    \I__11893\ : InMux
    port map (
            O => \N__51040\,
            I => \N__50938\
        );

    \I__11892\ : Span4Mux_v
    port map (
            O => \N__51037\,
            I => \N__50929\
        );

    \I__11891\ : LocalMux
    port map (
            O => \N__51034\,
            I => \N__50929\
        );

    \I__11890\ : LocalMux
    port map (
            O => \N__51031\,
            I => \N__50929\
        );

    \I__11889\ : LocalMux
    port map (
            O => \N__51028\,
            I => \N__50929\
        );

    \I__11888\ : InMux
    port map (
            O => \N__51027\,
            I => \N__50926\
        );

    \I__11887\ : InMux
    port map (
            O => \N__51026\,
            I => \N__50923\
        );

    \I__11886\ : InMux
    port map (
            O => \N__51025\,
            I => \N__50920\
        );

    \I__11885\ : InMux
    port map (
            O => \N__51024\,
            I => \N__50917\
        );

    \I__11884\ : Span4Mux_v
    port map (
            O => \N__51017\,
            I => \N__50914\
        );

    \I__11883\ : Span4Mux_v
    port map (
            O => \N__51010\,
            I => \N__50905\
        );

    \I__11882\ : LocalMux
    port map (
            O => \N__51007\,
            I => \N__50905\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__51004\,
            I => \N__50905\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__51001\,
            I => \N__50905\
        );

    \I__11879\ : Span4Mux_v
    port map (
            O => \N__50994\,
            I => \N__50898\
        );

    \I__11878\ : LocalMux
    port map (
            O => \N__50991\,
            I => \N__50898\
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__50988\,
            I => \N__50898\
        );

    \I__11876\ : InMux
    port map (
            O => \N__50987\,
            I => \N__50895\
        );

    \I__11875\ : InMux
    port map (
            O => \N__50986\,
            I => \N__50892\
        );

    \I__11874\ : LocalMux
    port map (
            O => \N__50983\,
            I => \N__50889\
        );

    \I__11873\ : InMux
    port map (
            O => \N__50982\,
            I => \N__50886\
        );

    \I__11872\ : InMux
    port map (
            O => \N__50981\,
            I => \N__50883\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__50978\,
            I => \N__50874\
        );

    \I__11870\ : LocalMux
    port map (
            O => \N__50975\,
            I => \N__50874\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__50972\,
            I => \N__50874\
        );

    \I__11868\ : Span4Mux_v
    port map (
            O => \N__50967\,
            I => \N__50867\
        );

    \I__11867\ : Span4Mux_v
    port map (
            O => \N__50956\,
            I => \N__50867\
        );

    \I__11866\ : Span4Mux_h
    port map (
            O => \N__50953\,
            I => \N__50860\
        );

    \I__11865\ : Span4Mux_v
    port map (
            O => \N__50944\,
            I => \N__50860\
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__50941\,
            I => \N__50860\
        );

    \I__11863\ : LocalMux
    port map (
            O => \N__50938\,
            I => \N__50857\
        );

    \I__11862\ : Span4Mux_v
    port map (
            O => \N__50929\,
            I => \N__50846\
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__50926\,
            I => \N__50846\
        );

    \I__11860\ : LocalMux
    port map (
            O => \N__50923\,
            I => \N__50846\
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__50920\,
            I => \N__50846\
        );

    \I__11858\ : LocalMux
    port map (
            O => \N__50917\,
            I => \N__50846\
        );

    \I__11857\ : Span4Mux_h
    port map (
            O => \N__50914\,
            I => \N__50835\
        );

    \I__11856\ : Span4Mux_v
    port map (
            O => \N__50905\,
            I => \N__50835\
        );

    \I__11855\ : Span4Mux_h
    port map (
            O => \N__50898\,
            I => \N__50835\
        );

    \I__11854\ : LocalMux
    port map (
            O => \N__50895\,
            I => \N__50835\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__50892\,
            I => \N__50835\
        );

    \I__11852\ : Sp12to4
    port map (
            O => \N__50889\,
            I => \N__50828\
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__50886\,
            I => \N__50828\
        );

    \I__11850\ : LocalMux
    port map (
            O => \N__50883\,
            I => \N__50828\
        );

    \I__11849\ : InMux
    port map (
            O => \N__50882\,
            I => \N__50825\
        );

    \I__11848\ : InMux
    port map (
            O => \N__50881\,
            I => \N__50822\
        );

    \I__11847\ : Span4Mux_v
    port map (
            O => \N__50874\,
            I => \N__50819\
        );

    \I__11846\ : InMux
    port map (
            O => \N__50873\,
            I => \N__50814\
        );

    \I__11845\ : InMux
    port map (
            O => \N__50872\,
            I => \N__50814\
        );

    \I__11844\ : Span4Mux_h
    port map (
            O => \N__50867\,
            I => \N__50807\
        );

    \I__11843\ : Span4Mux_v
    port map (
            O => \N__50860\,
            I => \N__50807\
        );

    \I__11842\ : Span4Mux_v
    port map (
            O => \N__50857\,
            I => \N__50807\
        );

    \I__11841\ : Span4Mux_v
    port map (
            O => \N__50846\,
            I => \N__50804\
        );

    \I__11840\ : Span4Mux_h
    port map (
            O => \N__50835\,
            I => \N__50801\
        );

    \I__11839\ : Span12Mux_v
    port map (
            O => \N__50828\,
            I => \N__50796\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__50825\,
            I => \N__50796\
        );

    \I__11837\ : LocalMux
    port map (
            O => \N__50822\,
            I => \N__50789\
        );

    \I__11836\ : Sp12to4
    port map (
            O => \N__50819\,
            I => \N__50789\
        );

    \I__11835\ : LocalMux
    port map (
            O => \N__50814\,
            I => \N__50789\
        );

    \I__11834\ : Odrv4
    port map (
            O => \N__50807\,
            I => spi_data_mosi_0
        );

    \I__11833\ : Odrv4
    port map (
            O => \N__50804\,
            I => spi_data_mosi_0
        );

    \I__11832\ : Odrv4
    port map (
            O => \N__50801\,
            I => spi_data_mosi_0
        );

    \I__11831\ : Odrv12
    port map (
            O => \N__50796\,
            I => spi_data_mosi_0
        );

    \I__11830\ : Odrv12
    port map (
            O => \N__50789\,
            I => spi_data_mosi_0
        );

    \I__11829\ : InMux
    port map (
            O => \N__50778\,
            I => \N__50775\
        );

    \I__11828\ : LocalMux
    port map (
            O => \N__50775\,
            I => \sDAC_mem_13Z0Z_0\
        );

    \I__11827\ : InMux
    port map (
            O => \N__50772\,
            I => \N__50766\
        );

    \I__11826\ : InMux
    port map (
            O => \N__50771\,
            I => \N__50763\
        );

    \I__11825\ : InMux
    port map (
            O => \N__50770\,
            I => \N__50758\
        );

    \I__11824\ : InMux
    port map (
            O => \N__50769\,
            I => \N__50755\
        );

    \I__11823\ : LocalMux
    port map (
            O => \N__50766\,
            I => \N__50750\
        );

    \I__11822\ : LocalMux
    port map (
            O => \N__50763\,
            I => \N__50747\
        );

    \I__11821\ : InMux
    port map (
            O => \N__50762\,
            I => \N__50744\
        );

    \I__11820\ : InMux
    port map (
            O => \N__50761\,
            I => \N__50741\
        );

    \I__11819\ : LocalMux
    port map (
            O => \N__50758\,
            I => \N__50735\
        );

    \I__11818\ : LocalMux
    port map (
            O => \N__50755\,
            I => \N__50735\
        );

    \I__11817\ : InMux
    port map (
            O => \N__50754\,
            I => \N__50729\
        );

    \I__11816\ : InMux
    port map (
            O => \N__50753\,
            I => \N__50726\
        );

    \I__11815\ : Span4Mux_v
    port map (
            O => \N__50750\,
            I => \N__50714\
        );

    \I__11814\ : Span4Mux_v
    port map (
            O => \N__50747\,
            I => \N__50714\
        );

    \I__11813\ : LocalMux
    port map (
            O => \N__50744\,
            I => \N__50714\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__50741\,
            I => \N__50714\
        );

    \I__11811\ : InMux
    port map (
            O => \N__50740\,
            I => \N__50711\
        );

    \I__11810\ : Span4Mux_v
    port map (
            O => \N__50735\,
            I => \N__50704\
        );

    \I__11809\ : InMux
    port map (
            O => \N__50734\,
            I => \N__50701\
        );

    \I__11808\ : InMux
    port map (
            O => \N__50733\,
            I => \N__50698\
        );

    \I__11807\ : InMux
    port map (
            O => \N__50732\,
            I => \N__50695\
        );

    \I__11806\ : LocalMux
    port map (
            O => \N__50729\,
            I => \N__50688\
        );

    \I__11805\ : LocalMux
    port map (
            O => \N__50726\,
            I => \N__50682\
        );

    \I__11804\ : InMux
    port map (
            O => \N__50725\,
            I => \N__50679\
        );

    \I__11803\ : InMux
    port map (
            O => \N__50724\,
            I => \N__50669\
        );

    \I__11802\ : InMux
    port map (
            O => \N__50723\,
            I => \N__50666\
        );

    \I__11801\ : Span4Mux_v
    port map (
            O => \N__50714\,
            I => \N__50659\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__50711\,
            I => \N__50659\
        );

    \I__11799\ : InMux
    port map (
            O => \N__50710\,
            I => \N__50656\
        );

    \I__11798\ : InMux
    port map (
            O => \N__50709\,
            I => \N__50653\
        );

    \I__11797\ : InMux
    port map (
            O => \N__50708\,
            I => \N__50650\
        );

    \I__11796\ : InMux
    port map (
            O => \N__50707\,
            I => \N__50647\
        );

    \I__11795\ : Span4Mux_h
    port map (
            O => \N__50704\,
            I => \N__50638\
        );

    \I__11794\ : LocalMux
    port map (
            O => \N__50701\,
            I => \N__50638\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__50698\,
            I => \N__50638\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__50695\,
            I => \N__50638\
        );

    \I__11791\ : InMux
    port map (
            O => \N__50694\,
            I => \N__50635\
        );

    \I__11790\ : InMux
    port map (
            O => \N__50693\,
            I => \N__50632\
        );

    \I__11789\ : InMux
    port map (
            O => \N__50692\,
            I => \N__50629\
        );

    \I__11788\ : InMux
    port map (
            O => \N__50691\,
            I => \N__50626\
        );

    \I__11787\ : Span4Mux_v
    port map (
            O => \N__50688\,
            I => \N__50622\
        );

    \I__11786\ : InMux
    port map (
            O => \N__50687\,
            I => \N__50619\
        );

    \I__11785\ : InMux
    port map (
            O => \N__50686\,
            I => \N__50616\
        );

    \I__11784\ : InMux
    port map (
            O => \N__50685\,
            I => \N__50613\
        );

    \I__11783\ : Span4Mux_v
    port map (
            O => \N__50682\,
            I => \N__50608\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__50679\,
            I => \N__50608\
        );

    \I__11781\ : InMux
    port map (
            O => \N__50678\,
            I => \N__50605\
        );

    \I__11780\ : InMux
    port map (
            O => \N__50677\,
            I => \N__50602\
        );

    \I__11779\ : InMux
    port map (
            O => \N__50676\,
            I => \N__50596\
        );

    \I__11778\ : InMux
    port map (
            O => \N__50675\,
            I => \N__50593\
        );

    \I__11777\ : InMux
    port map (
            O => \N__50674\,
            I => \N__50589\
        );

    \I__11776\ : InMux
    port map (
            O => \N__50673\,
            I => \N__50586\
        );

    \I__11775\ : InMux
    port map (
            O => \N__50672\,
            I => \N__50577\
        );

    \I__11774\ : LocalMux
    port map (
            O => \N__50669\,
            I => \N__50567\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__50666\,
            I => \N__50567\
        );

    \I__11772\ : InMux
    port map (
            O => \N__50665\,
            I => \N__50564\
        );

    \I__11771\ : InMux
    port map (
            O => \N__50664\,
            I => \N__50561\
        );

    \I__11770\ : Span4Mux_v
    port map (
            O => \N__50659\,
            I => \N__50549\
        );

    \I__11769\ : LocalMux
    port map (
            O => \N__50656\,
            I => \N__50549\
        );

    \I__11768\ : LocalMux
    port map (
            O => \N__50653\,
            I => \N__50549\
        );

    \I__11767\ : LocalMux
    port map (
            O => \N__50650\,
            I => \N__50549\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__50647\,
            I => \N__50549\
        );

    \I__11765\ : Span4Mux_v
    port map (
            O => \N__50638\,
            I => \N__50542\
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__50635\,
            I => \N__50542\
        );

    \I__11763\ : LocalMux
    port map (
            O => \N__50632\,
            I => \N__50542\
        );

    \I__11762\ : LocalMux
    port map (
            O => \N__50629\,
            I => \N__50537\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__50626\,
            I => \N__50537\
        );

    \I__11760\ : InMux
    port map (
            O => \N__50625\,
            I => \N__50534\
        );

    \I__11759\ : Span4Mux_v
    port map (
            O => \N__50622\,
            I => \N__50525\
        );

    \I__11758\ : LocalMux
    port map (
            O => \N__50619\,
            I => \N__50525\
        );

    \I__11757\ : LocalMux
    port map (
            O => \N__50616\,
            I => \N__50525\
        );

    \I__11756\ : LocalMux
    port map (
            O => \N__50613\,
            I => \N__50525\
        );

    \I__11755\ : Span4Mux_v
    port map (
            O => \N__50608\,
            I => \N__50518\
        );

    \I__11754\ : LocalMux
    port map (
            O => \N__50605\,
            I => \N__50518\
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__50602\,
            I => \N__50518\
        );

    \I__11752\ : InMux
    port map (
            O => \N__50601\,
            I => \N__50515\
        );

    \I__11751\ : InMux
    port map (
            O => \N__50600\,
            I => \N__50512\
        );

    \I__11750\ : InMux
    port map (
            O => \N__50599\,
            I => \N__50509\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__50596\,
            I => \N__50504\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__50593\,
            I => \N__50504\
        );

    \I__11747\ : InMux
    port map (
            O => \N__50592\,
            I => \N__50501\
        );

    \I__11746\ : LocalMux
    port map (
            O => \N__50589\,
            I => \N__50497\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__50586\,
            I => \N__50494\
        );

    \I__11744\ : InMux
    port map (
            O => \N__50585\,
            I => \N__50491\
        );

    \I__11743\ : InMux
    port map (
            O => \N__50584\,
            I => \N__50488\
        );

    \I__11742\ : InMux
    port map (
            O => \N__50583\,
            I => \N__50485\
        );

    \I__11741\ : InMux
    port map (
            O => \N__50582\,
            I => \N__50482\
        );

    \I__11740\ : InMux
    port map (
            O => \N__50581\,
            I => \N__50479\
        );

    \I__11739\ : InMux
    port map (
            O => \N__50580\,
            I => \N__50476\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__50577\,
            I => \N__50473\
        );

    \I__11737\ : InMux
    port map (
            O => \N__50576\,
            I => \N__50470\
        );

    \I__11736\ : InMux
    port map (
            O => \N__50575\,
            I => \N__50467\
        );

    \I__11735\ : InMux
    port map (
            O => \N__50574\,
            I => \N__50464\
        );

    \I__11734\ : InMux
    port map (
            O => \N__50573\,
            I => \N__50461\
        );

    \I__11733\ : InMux
    port map (
            O => \N__50572\,
            I => \N__50458\
        );

    \I__11732\ : Span4Mux_v
    port map (
            O => \N__50567\,
            I => \N__50451\
        );

    \I__11731\ : LocalMux
    port map (
            O => \N__50564\,
            I => \N__50448\
        );

    \I__11730\ : LocalMux
    port map (
            O => \N__50561\,
            I => \N__50445\
        );

    \I__11729\ : InMux
    port map (
            O => \N__50560\,
            I => \N__50442\
        );

    \I__11728\ : Span4Mux_v
    port map (
            O => \N__50549\,
            I => \N__50439\
        );

    \I__11727\ : Span4Mux_v
    port map (
            O => \N__50542\,
            I => \N__50432\
        );

    \I__11726\ : Span4Mux_h
    port map (
            O => \N__50537\,
            I => \N__50432\
        );

    \I__11725\ : LocalMux
    port map (
            O => \N__50534\,
            I => \N__50432\
        );

    \I__11724\ : Span4Mux_v
    port map (
            O => \N__50525\,
            I => \N__50423\
        );

    \I__11723\ : Span4Mux_h
    port map (
            O => \N__50518\,
            I => \N__50423\
        );

    \I__11722\ : LocalMux
    port map (
            O => \N__50515\,
            I => \N__50423\
        );

    \I__11721\ : LocalMux
    port map (
            O => \N__50512\,
            I => \N__50423\
        );

    \I__11720\ : LocalMux
    port map (
            O => \N__50509\,
            I => \N__50415\
        );

    \I__11719\ : Sp12to4
    port map (
            O => \N__50504\,
            I => \N__50415\
        );

    \I__11718\ : LocalMux
    port map (
            O => \N__50501\,
            I => \N__50415\
        );

    \I__11717\ : InMux
    port map (
            O => \N__50500\,
            I => \N__50412\
        );

    \I__11716\ : Span12Mux_s11_v
    port map (
            O => \N__50497\,
            I => \N__50393\
        );

    \I__11715\ : Sp12to4
    port map (
            O => \N__50494\,
            I => \N__50393\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__50491\,
            I => \N__50393\
        );

    \I__11713\ : LocalMux
    port map (
            O => \N__50488\,
            I => \N__50393\
        );

    \I__11712\ : LocalMux
    port map (
            O => \N__50485\,
            I => \N__50393\
        );

    \I__11711\ : LocalMux
    port map (
            O => \N__50482\,
            I => \N__50393\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__50479\,
            I => \N__50393\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__50476\,
            I => \N__50393\
        );

    \I__11708\ : Sp12to4
    port map (
            O => \N__50473\,
            I => \N__50393\
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__50470\,
            I => \N__50386\
        );

    \I__11706\ : LocalMux
    port map (
            O => \N__50467\,
            I => \N__50386\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__50464\,
            I => \N__50386\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__50461\,
            I => \N__50381\
        );

    \I__11703\ : LocalMux
    port map (
            O => \N__50458\,
            I => \N__50381\
        );

    \I__11702\ : InMux
    port map (
            O => \N__50457\,
            I => \N__50378\
        );

    \I__11701\ : InMux
    port map (
            O => \N__50456\,
            I => \N__50375\
        );

    \I__11700\ : InMux
    port map (
            O => \N__50455\,
            I => \N__50372\
        );

    \I__11699\ : InMux
    port map (
            O => \N__50454\,
            I => \N__50369\
        );

    \I__11698\ : Span4Mux_h
    port map (
            O => \N__50451\,
            I => \N__50360\
        );

    \I__11697\ : Span4Mux_h
    port map (
            O => \N__50448\,
            I => \N__50360\
        );

    \I__11696\ : Span4Mux_v
    port map (
            O => \N__50445\,
            I => \N__50360\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__50442\,
            I => \N__50360\
        );

    \I__11694\ : Span4Mux_h
    port map (
            O => \N__50439\,
            I => \N__50355\
        );

    \I__11693\ : Span4Mux_v
    port map (
            O => \N__50432\,
            I => \N__50355\
        );

    \I__11692\ : Span4Mux_h
    port map (
            O => \N__50423\,
            I => \N__50352\
        );

    \I__11691\ : InMux
    port map (
            O => \N__50422\,
            I => \N__50349\
        );

    \I__11690\ : Span12Mux_v
    port map (
            O => \N__50415\,
            I => \N__50342\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__50412\,
            I => \N__50342\
        );

    \I__11688\ : Span12Mux_v
    port map (
            O => \N__50393\,
            I => \N__50342\
        );

    \I__11687\ : Span12Mux_h
    port map (
            O => \N__50386\,
            I => \N__50327\
        );

    \I__11686\ : Span12Mux_v
    port map (
            O => \N__50381\,
            I => \N__50327\
        );

    \I__11685\ : LocalMux
    port map (
            O => \N__50378\,
            I => \N__50327\
        );

    \I__11684\ : LocalMux
    port map (
            O => \N__50375\,
            I => \N__50327\
        );

    \I__11683\ : LocalMux
    port map (
            O => \N__50372\,
            I => \N__50327\
        );

    \I__11682\ : LocalMux
    port map (
            O => \N__50369\,
            I => \N__50327\
        );

    \I__11681\ : Sp12to4
    port map (
            O => \N__50360\,
            I => \N__50327\
        );

    \I__11680\ : Odrv4
    port map (
            O => \N__50355\,
            I => spi_data_mosi_1
        );

    \I__11679\ : Odrv4
    port map (
            O => \N__50352\,
            I => spi_data_mosi_1
        );

    \I__11678\ : LocalMux
    port map (
            O => \N__50349\,
            I => spi_data_mosi_1
        );

    \I__11677\ : Odrv12
    port map (
            O => \N__50342\,
            I => spi_data_mosi_1
        );

    \I__11676\ : Odrv12
    port map (
            O => \N__50327\,
            I => spi_data_mosi_1
        );

    \I__11675\ : InMux
    port map (
            O => \N__50316\,
            I => \N__50313\
        );

    \I__11674\ : LocalMux
    port map (
            O => \N__50313\,
            I => \sDAC_mem_13Z0Z_1\
        );

    \I__11673\ : InMux
    port map (
            O => \N__50310\,
            I => \N__50302\
        );

    \I__11672\ : InMux
    port map (
            O => \N__50309\,
            I => \N__50296\
        );

    \I__11671\ : InMux
    port map (
            O => \N__50308\,
            I => \N__50293\
        );

    \I__11670\ : InMux
    port map (
            O => \N__50307\,
            I => \N__50288\
        );

    \I__11669\ : InMux
    port map (
            O => \N__50306\,
            I => \N__50278\
        );

    \I__11668\ : InMux
    port map (
            O => \N__50305\,
            I => \N__50275\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__50302\,
            I => \N__50271\
        );

    \I__11666\ : InMux
    port map (
            O => \N__50301\,
            I => \N__50268\
        );

    \I__11665\ : InMux
    port map (
            O => \N__50300\,
            I => \N__50265\
        );

    \I__11664\ : InMux
    port map (
            O => \N__50299\,
            I => \N__50258\
        );

    \I__11663\ : LocalMux
    port map (
            O => \N__50296\,
            I => \N__50250\
        );

    \I__11662\ : LocalMux
    port map (
            O => \N__50293\,
            I => \N__50250\
        );

    \I__11661\ : InMux
    port map (
            O => \N__50292\,
            I => \N__50247\
        );

    \I__11660\ : InMux
    port map (
            O => \N__50291\,
            I => \N__50244\
        );

    \I__11659\ : LocalMux
    port map (
            O => \N__50288\,
            I => \N__50237\
        );

    \I__11658\ : InMux
    port map (
            O => \N__50287\,
            I => \N__50234\
        );

    \I__11657\ : InMux
    port map (
            O => \N__50286\,
            I => \N__50231\
        );

    \I__11656\ : InMux
    port map (
            O => \N__50285\,
            I => \N__50227\
        );

    \I__11655\ : InMux
    port map (
            O => \N__50284\,
            I => \N__50224\
        );

    \I__11654\ : InMux
    port map (
            O => \N__50283\,
            I => \N__50221\
        );

    \I__11653\ : InMux
    port map (
            O => \N__50282\,
            I => \N__50218\
        );

    \I__11652\ : InMux
    port map (
            O => \N__50281\,
            I => \N__50215\
        );

    \I__11651\ : LocalMux
    port map (
            O => \N__50278\,
            I => \N__50210\
        );

    \I__11650\ : LocalMux
    port map (
            O => \N__50275\,
            I => \N__50210\
        );

    \I__11649\ : InMux
    port map (
            O => \N__50274\,
            I => \N__50207\
        );

    \I__11648\ : Span4Mux_v
    port map (
            O => \N__50271\,
            I => \N__50200\
        );

    \I__11647\ : LocalMux
    port map (
            O => \N__50268\,
            I => \N__50200\
        );

    \I__11646\ : LocalMux
    port map (
            O => \N__50265\,
            I => \N__50200\
        );

    \I__11645\ : InMux
    port map (
            O => \N__50264\,
            I => \N__50197\
        );

    \I__11644\ : InMux
    port map (
            O => \N__50263\,
            I => \N__50194\
        );

    \I__11643\ : InMux
    port map (
            O => \N__50262\,
            I => \N__50191\
        );

    \I__11642\ : InMux
    port map (
            O => \N__50261\,
            I => \N__50188\
        );

    \I__11641\ : LocalMux
    port map (
            O => \N__50258\,
            I => \N__50184\
        );

    \I__11640\ : InMux
    port map (
            O => \N__50257\,
            I => \N__50181\
        );

    \I__11639\ : InMux
    port map (
            O => \N__50256\,
            I => \N__50175\
        );

    \I__11638\ : InMux
    port map (
            O => \N__50255\,
            I => \N__50171\
        );

    \I__11637\ : Span4Mux_v
    port map (
            O => \N__50250\,
            I => \N__50164\
        );

    \I__11636\ : LocalMux
    port map (
            O => \N__50247\,
            I => \N__50164\
        );

    \I__11635\ : LocalMux
    port map (
            O => \N__50244\,
            I => \N__50164\
        );

    \I__11634\ : InMux
    port map (
            O => \N__50243\,
            I => \N__50161\
        );

    \I__11633\ : InMux
    port map (
            O => \N__50242\,
            I => \N__50158\
        );

    \I__11632\ : InMux
    port map (
            O => \N__50241\,
            I => \N__50155\
        );

    \I__11631\ : InMux
    port map (
            O => \N__50240\,
            I => \N__50152\
        );

    \I__11630\ : Span4Mux_v
    port map (
            O => \N__50237\,
            I => \N__50144\
        );

    \I__11629\ : LocalMux
    port map (
            O => \N__50234\,
            I => \N__50144\
        );

    \I__11628\ : LocalMux
    port map (
            O => \N__50231\,
            I => \N__50144\
        );

    \I__11627\ : InMux
    port map (
            O => \N__50230\,
            I => \N__50141\
        );

    \I__11626\ : LocalMux
    port map (
            O => \N__50227\,
            I => \N__50132\
        );

    \I__11625\ : LocalMux
    port map (
            O => \N__50224\,
            I => \N__50132\
        );

    \I__11624\ : LocalMux
    port map (
            O => \N__50221\,
            I => \N__50132\
        );

    \I__11623\ : LocalMux
    port map (
            O => \N__50218\,
            I => \N__50132\
        );

    \I__11622\ : LocalMux
    port map (
            O => \N__50215\,
            I => \N__50129\
        );

    \I__11621\ : Span4Mux_v
    port map (
            O => \N__50210\,
            I => \N__50124\
        );

    \I__11620\ : LocalMux
    port map (
            O => \N__50207\,
            I => \N__50124\
        );

    \I__11619\ : Span4Mux_v
    port map (
            O => \N__50200\,
            I => \N__50112\
        );

    \I__11618\ : LocalMux
    port map (
            O => \N__50197\,
            I => \N__50112\
        );

    \I__11617\ : LocalMux
    port map (
            O => \N__50194\,
            I => \N__50112\
        );

    \I__11616\ : LocalMux
    port map (
            O => \N__50191\,
            I => \N__50112\
        );

    \I__11615\ : LocalMux
    port map (
            O => \N__50188\,
            I => \N__50112\
        );

    \I__11614\ : InMux
    port map (
            O => \N__50187\,
            I => \N__50109\
        );

    \I__11613\ : Span4Mux_h
    port map (
            O => \N__50184\,
            I => \N__50100\
        );

    \I__11612\ : LocalMux
    port map (
            O => \N__50181\,
            I => \N__50100\
        );

    \I__11611\ : InMux
    port map (
            O => \N__50180\,
            I => \N__50097\
        );

    \I__11610\ : InMux
    port map (
            O => \N__50179\,
            I => \N__50094\
        );

    \I__11609\ : InMux
    port map (
            O => \N__50178\,
            I => \N__50087\
        );

    \I__11608\ : LocalMux
    port map (
            O => \N__50175\,
            I => \N__50084\
        );

    \I__11607\ : InMux
    port map (
            O => \N__50174\,
            I => \N__50081\
        );

    \I__11606\ : LocalMux
    port map (
            O => \N__50171\,
            I => \N__50074\
        );

    \I__11605\ : Span4Mux_h
    port map (
            O => \N__50164\,
            I => \N__50063\
        );

    \I__11604\ : LocalMux
    port map (
            O => \N__50161\,
            I => \N__50063\
        );

    \I__11603\ : LocalMux
    port map (
            O => \N__50158\,
            I => \N__50063\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__50155\,
            I => \N__50063\
        );

    \I__11601\ : LocalMux
    port map (
            O => \N__50152\,
            I => \N__50063\
        );

    \I__11600\ : InMux
    port map (
            O => \N__50151\,
            I => \N__50060\
        );

    \I__11599\ : Span4Mux_v
    port map (
            O => \N__50144\,
            I => \N__50055\
        );

    \I__11598\ : LocalMux
    port map (
            O => \N__50141\,
            I => \N__50055\
        );

    \I__11597\ : Span4Mux_v
    port map (
            O => \N__50132\,
            I => \N__50052\
        );

    \I__11596\ : Span4Mux_h
    port map (
            O => \N__50129\,
            I => \N__50047\
        );

    \I__11595\ : Span4Mux_v
    port map (
            O => \N__50124\,
            I => \N__50047\
        );

    \I__11594\ : InMux
    port map (
            O => \N__50123\,
            I => \N__50044\
        );

    \I__11593\ : Span4Mux_v
    port map (
            O => \N__50112\,
            I => \N__50039\
        );

    \I__11592\ : LocalMux
    port map (
            O => \N__50109\,
            I => \N__50039\
        );

    \I__11591\ : InMux
    port map (
            O => \N__50108\,
            I => \N__50036\
        );

    \I__11590\ : InMux
    port map (
            O => \N__50107\,
            I => \N__50033\
        );

    \I__11589\ : InMux
    port map (
            O => \N__50106\,
            I => \N__50030\
        );

    \I__11588\ : InMux
    port map (
            O => \N__50105\,
            I => \N__50027\
        );

    \I__11587\ : Span4Mux_v
    port map (
            O => \N__50100\,
            I => \N__50016\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__50097\,
            I => \N__50016\
        );

    \I__11585\ : LocalMux
    port map (
            O => \N__50094\,
            I => \N__50016\
        );

    \I__11584\ : InMux
    port map (
            O => \N__50093\,
            I => \N__50013\
        );

    \I__11583\ : InMux
    port map (
            O => \N__50092\,
            I => \N__50010\
        );

    \I__11582\ : InMux
    port map (
            O => \N__50091\,
            I => \N__50007\
        );

    \I__11581\ : InMux
    port map (
            O => \N__50090\,
            I => \N__50001\
        );

    \I__11580\ : LocalMux
    port map (
            O => \N__50087\,
            I => \N__49998\
        );

    \I__11579\ : Span4Mux_v
    port map (
            O => \N__50084\,
            I => \N__49993\
        );

    \I__11578\ : LocalMux
    port map (
            O => \N__50081\,
            I => \N__49993\
        );

    \I__11577\ : InMux
    port map (
            O => \N__50080\,
            I => \N__49990\
        );

    \I__11576\ : InMux
    port map (
            O => \N__50079\,
            I => \N__49987\
        );

    \I__11575\ : InMux
    port map (
            O => \N__50078\,
            I => \N__49984\
        );

    \I__11574\ : InMux
    port map (
            O => \N__50077\,
            I => \N__49981\
        );

    \I__11573\ : Span4Mux_h
    port map (
            O => \N__50074\,
            I => \N__49974\
        );

    \I__11572\ : Span4Mux_v
    port map (
            O => \N__50063\,
            I => \N__49974\
        );

    \I__11571\ : LocalMux
    port map (
            O => \N__50060\,
            I => \N__49974\
        );

    \I__11570\ : Span4Mux_v
    port map (
            O => \N__50055\,
            I => \N__49971\
        );

    \I__11569\ : Span4Mux_h
    port map (
            O => \N__50052\,
            I => \N__49964\
        );

    \I__11568\ : Span4Mux_v
    port map (
            O => \N__50047\,
            I => \N__49964\
        );

    \I__11567\ : LocalMux
    port map (
            O => \N__50044\,
            I => \N__49964\
        );

    \I__11566\ : Span4Mux_v
    port map (
            O => \N__50039\,
            I => \N__49955\
        );

    \I__11565\ : LocalMux
    port map (
            O => \N__50036\,
            I => \N__49955\
        );

    \I__11564\ : LocalMux
    port map (
            O => \N__50033\,
            I => \N__49955\
        );

    \I__11563\ : LocalMux
    port map (
            O => \N__50030\,
            I => \N__49955\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__50027\,
            I => \N__49952\
        );

    \I__11561\ : InMux
    port map (
            O => \N__50026\,
            I => \N__49949\
        );

    \I__11560\ : InMux
    port map (
            O => \N__50025\,
            I => \N__49946\
        );

    \I__11559\ : InMux
    port map (
            O => \N__50024\,
            I => \N__49943\
        );

    \I__11558\ : InMux
    port map (
            O => \N__50023\,
            I => \N__49940\
        );

    \I__11557\ : Span4Mux_v
    port map (
            O => \N__50016\,
            I => \N__49931\
        );

    \I__11556\ : LocalMux
    port map (
            O => \N__50013\,
            I => \N__49931\
        );

    \I__11555\ : LocalMux
    port map (
            O => \N__50010\,
            I => \N__49931\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__50007\,
            I => \N__49931\
        );

    \I__11553\ : InMux
    port map (
            O => \N__50006\,
            I => \N__49928\
        );

    \I__11552\ : InMux
    port map (
            O => \N__50005\,
            I => \N__49925\
        );

    \I__11551\ : InMux
    port map (
            O => \N__50004\,
            I => \N__49922\
        );

    \I__11550\ : LocalMux
    port map (
            O => \N__50001\,
            I => \N__49907\
        );

    \I__11549\ : Span12Mux_h
    port map (
            O => \N__49998\,
            I => \N__49907\
        );

    \I__11548\ : Sp12to4
    port map (
            O => \N__49993\,
            I => \N__49907\
        );

    \I__11547\ : LocalMux
    port map (
            O => \N__49990\,
            I => \N__49907\
        );

    \I__11546\ : LocalMux
    port map (
            O => \N__49987\,
            I => \N__49907\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__49984\,
            I => \N__49907\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__49981\,
            I => \N__49907\
        );

    \I__11543\ : Span4Mux_h
    port map (
            O => \N__49974\,
            I => \N__49903\
        );

    \I__11542\ : Span4Mux_h
    port map (
            O => \N__49971\,
            I => \N__49896\
        );

    \I__11541\ : Span4Mux_v
    port map (
            O => \N__49964\,
            I => \N__49896\
        );

    \I__11540\ : Span4Mux_v
    port map (
            O => \N__49955\,
            I => \N__49896\
        );

    \I__11539\ : Span12Mux_h
    port map (
            O => \N__49952\,
            I => \N__49885\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__49949\,
            I => \N__49885\
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__49946\,
            I => \N__49885\
        );

    \I__11536\ : LocalMux
    port map (
            O => \N__49943\,
            I => \N__49885\
        );

    \I__11535\ : LocalMux
    port map (
            O => \N__49940\,
            I => \N__49885\
        );

    \I__11534\ : Span4Mux_v
    port map (
            O => \N__49931\,
            I => \N__49878\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__49928\,
            I => \N__49878\
        );

    \I__11532\ : LocalMux
    port map (
            O => \N__49925\,
            I => \N__49878\
        );

    \I__11531\ : LocalMux
    port map (
            O => \N__49922\,
            I => \N__49873\
        );

    \I__11530\ : Span12Mux_v
    port map (
            O => \N__49907\,
            I => \N__49873\
        );

    \I__11529\ : InMux
    port map (
            O => \N__49906\,
            I => \N__49870\
        );

    \I__11528\ : Odrv4
    port map (
            O => \N__49903\,
            I => spi_data_mosi_2
        );

    \I__11527\ : Odrv4
    port map (
            O => \N__49896\,
            I => spi_data_mosi_2
        );

    \I__11526\ : Odrv12
    port map (
            O => \N__49885\,
            I => spi_data_mosi_2
        );

    \I__11525\ : Odrv4
    port map (
            O => \N__49878\,
            I => spi_data_mosi_2
        );

    \I__11524\ : Odrv12
    port map (
            O => \N__49873\,
            I => spi_data_mosi_2
        );

    \I__11523\ : LocalMux
    port map (
            O => \N__49870\,
            I => spi_data_mosi_2
        );

    \I__11522\ : InMux
    port map (
            O => \N__49857\,
            I => \N__49854\
        );

    \I__11521\ : LocalMux
    port map (
            O => \N__49854\,
            I => \N__49851\
        );

    \I__11520\ : Span12Mux_v
    port map (
            O => \N__49851\,
            I => \N__49848\
        );

    \I__11519\ : Odrv12
    port map (
            O => \N__49848\,
            I => \sDAC_mem_13Z0Z_2\
        );

    \I__11518\ : InMux
    port map (
            O => \N__49845\,
            I => \N__49838\
        );

    \I__11517\ : InMux
    port map (
            O => \N__49844\,
            I => \N__49830\
        );

    \I__11516\ : InMux
    port map (
            O => \N__49843\,
            I => \N__49827\
        );

    \I__11515\ : InMux
    port map (
            O => \N__49842\,
            I => \N__49815\
        );

    \I__11514\ : InMux
    port map (
            O => \N__49841\,
            I => \N__49812\
        );

    \I__11513\ : LocalMux
    port map (
            O => \N__49838\,
            I => \N__49808\
        );

    \I__11512\ : InMux
    port map (
            O => \N__49837\,
            I => \N__49805\
        );

    \I__11511\ : InMux
    port map (
            O => \N__49836\,
            I => \N__49802\
        );

    \I__11510\ : InMux
    port map (
            O => \N__49835\,
            I => \N__49799\
        );

    \I__11509\ : InMux
    port map (
            O => \N__49834\,
            I => \N__49791\
        );

    \I__11508\ : InMux
    port map (
            O => \N__49833\,
            I => \N__49787\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__49830\,
            I => \N__49779\
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__49827\,
            I => \N__49779\
        );

    \I__11505\ : InMux
    port map (
            O => \N__49826\,
            I => \N__49776\
        );

    \I__11504\ : InMux
    port map (
            O => \N__49825\,
            I => \N__49773\
        );

    \I__11503\ : InMux
    port map (
            O => \N__49824\,
            I => \N__49770\
        );

    \I__11502\ : InMux
    port map (
            O => \N__49823\,
            I => \N__49762\
        );

    \I__11501\ : InMux
    port map (
            O => \N__49822\,
            I => \N__49759\
        );

    \I__11500\ : InMux
    port map (
            O => \N__49821\,
            I => \N__49756\
        );

    \I__11499\ : InMux
    port map (
            O => \N__49820\,
            I => \N__49753\
        );

    \I__11498\ : InMux
    port map (
            O => \N__49819\,
            I => \N__49750\
        );

    \I__11497\ : InMux
    port map (
            O => \N__49818\,
            I => \N__49747\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__49815\,
            I => \N__49744\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__49812\,
            I => \N__49741\
        );

    \I__11494\ : InMux
    port map (
            O => \N__49811\,
            I => \N__49738\
        );

    \I__11493\ : Span4Mux_h
    port map (
            O => \N__49808\,
            I => \N__49729\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__49805\,
            I => \N__49729\
        );

    \I__11491\ : LocalMux
    port map (
            O => \N__49802\,
            I => \N__49726\
        );

    \I__11490\ : LocalMux
    port map (
            O => \N__49799\,
            I => \N__49723\
        );

    \I__11489\ : InMux
    port map (
            O => \N__49798\,
            I => \N__49720\
        );

    \I__11488\ : InMux
    port map (
            O => \N__49797\,
            I => \N__49717\
        );

    \I__11487\ : InMux
    port map (
            O => \N__49796\,
            I => \N__49714\
        );

    \I__11486\ : InMux
    port map (
            O => \N__49795\,
            I => \N__49711\
        );

    \I__11485\ : InMux
    port map (
            O => \N__49794\,
            I => \N__49708\
        );

    \I__11484\ : LocalMux
    port map (
            O => \N__49791\,
            I => \N__49705\
        );

    \I__11483\ : InMux
    port map (
            O => \N__49790\,
            I => \N__49699\
        );

    \I__11482\ : LocalMux
    port map (
            O => \N__49787\,
            I => \N__49696\
        );

    \I__11481\ : InMux
    port map (
            O => \N__49786\,
            I => \N__49693\
        );

    \I__11480\ : InMux
    port map (
            O => \N__49785\,
            I => \N__49690\
        );

    \I__11479\ : InMux
    port map (
            O => \N__49784\,
            I => \N__49686\
        );

    \I__11478\ : Span4Mux_v
    port map (
            O => \N__49779\,
            I => \N__49677\
        );

    \I__11477\ : LocalMux
    port map (
            O => \N__49776\,
            I => \N__49677\
        );

    \I__11476\ : LocalMux
    port map (
            O => \N__49773\,
            I => \N__49677\
        );

    \I__11475\ : LocalMux
    port map (
            O => \N__49770\,
            I => \N__49677\
        );

    \I__11474\ : InMux
    port map (
            O => \N__49769\,
            I => \N__49674\
        );

    \I__11473\ : InMux
    port map (
            O => \N__49768\,
            I => \N__49671\
        );

    \I__11472\ : InMux
    port map (
            O => \N__49767\,
            I => \N__49668\
        );

    \I__11471\ : InMux
    port map (
            O => \N__49766\,
            I => \N__49665\
        );

    \I__11470\ : InMux
    port map (
            O => \N__49765\,
            I => \N__49662\
        );

    \I__11469\ : LocalMux
    port map (
            O => \N__49762\,
            I => \N__49652\
        );

    \I__11468\ : LocalMux
    port map (
            O => \N__49759\,
            I => \N__49652\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__49756\,
            I => \N__49652\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__49753\,
            I => \N__49652\
        );

    \I__11465\ : LocalMux
    port map (
            O => \N__49750\,
            I => \N__49646\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__49747\,
            I => \N__49646\
        );

    \I__11463\ : Span4Mux_v
    port map (
            O => \N__49744\,
            I => \N__49639\
        );

    \I__11462\ : Span4Mux_v
    port map (
            O => \N__49741\,
            I => \N__49639\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__49738\,
            I => \N__49639\
        );

    \I__11460\ : InMux
    port map (
            O => \N__49737\,
            I => \N__49636\
        );

    \I__11459\ : InMux
    port map (
            O => \N__49736\,
            I => \N__49633\
        );

    \I__11458\ : InMux
    port map (
            O => \N__49735\,
            I => \N__49630\
        );

    \I__11457\ : InMux
    port map (
            O => \N__49734\,
            I => \N__49627\
        );

    \I__11456\ : Span4Mux_v
    port map (
            O => \N__49729\,
            I => \N__49611\
        );

    \I__11455\ : Span4Mux_h
    port map (
            O => \N__49726\,
            I => \N__49611\
        );

    \I__11454\ : Span4Mux_v
    port map (
            O => \N__49723\,
            I => \N__49611\
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__49720\,
            I => \N__49611\
        );

    \I__11452\ : LocalMux
    port map (
            O => \N__49717\,
            I => \N__49611\
        );

    \I__11451\ : LocalMux
    port map (
            O => \N__49714\,
            I => \N__49611\
        );

    \I__11450\ : LocalMux
    port map (
            O => \N__49711\,
            I => \N__49611\
        );

    \I__11449\ : LocalMux
    port map (
            O => \N__49708\,
            I => \N__49605\
        );

    \I__11448\ : Span4Mux_h
    port map (
            O => \N__49705\,
            I => \N__49602\
        );

    \I__11447\ : InMux
    port map (
            O => \N__49704\,
            I => \N__49599\
        );

    \I__11446\ : InMux
    port map (
            O => \N__49703\,
            I => \N__49596\
        );

    \I__11445\ : InMux
    port map (
            O => \N__49702\,
            I => \N__49593\
        );

    \I__11444\ : LocalMux
    port map (
            O => \N__49699\,
            I => \N__49587\
        );

    \I__11443\ : Span4Mux_v
    port map (
            O => \N__49696\,
            I => \N__49582\
        );

    \I__11442\ : LocalMux
    port map (
            O => \N__49693\,
            I => \N__49582\
        );

    \I__11441\ : LocalMux
    port map (
            O => \N__49690\,
            I => \N__49579\
        );

    \I__11440\ : InMux
    port map (
            O => \N__49689\,
            I => \N__49576\
        );

    \I__11439\ : LocalMux
    port map (
            O => \N__49686\,
            I => \N__49568\
        );

    \I__11438\ : Span4Mux_h
    port map (
            O => \N__49677\,
            I => \N__49555\
        );

    \I__11437\ : LocalMux
    port map (
            O => \N__49674\,
            I => \N__49555\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__49671\,
            I => \N__49555\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__49668\,
            I => \N__49555\
        );

    \I__11434\ : LocalMux
    port map (
            O => \N__49665\,
            I => \N__49555\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__49662\,
            I => \N__49555\
        );

    \I__11432\ : InMux
    port map (
            O => \N__49661\,
            I => \N__49552\
        );

    \I__11431\ : Span4Mux_v
    port map (
            O => \N__49652\,
            I => \N__49549\
        );

    \I__11430\ : InMux
    port map (
            O => \N__49651\,
            I => \N__49546\
        );

    \I__11429\ : Span4Mux_v
    port map (
            O => \N__49646\,
            I => \N__49533\
        );

    \I__11428\ : Span4Mux_v
    port map (
            O => \N__49639\,
            I => \N__49533\
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__49636\,
            I => \N__49533\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__49633\,
            I => \N__49533\
        );

    \I__11425\ : LocalMux
    port map (
            O => \N__49630\,
            I => \N__49533\
        );

    \I__11424\ : LocalMux
    port map (
            O => \N__49627\,
            I => \N__49533\
        );

    \I__11423\ : InMux
    port map (
            O => \N__49626\,
            I => \N__49530\
        );

    \I__11422\ : Span4Mux_v
    port map (
            O => \N__49611\,
            I => \N__49527\
        );

    \I__11421\ : InMux
    port map (
            O => \N__49610\,
            I => \N__49524\
        );

    \I__11420\ : InMux
    port map (
            O => \N__49609\,
            I => \N__49521\
        );

    \I__11419\ : InMux
    port map (
            O => \N__49608\,
            I => \N__49518\
        );

    \I__11418\ : Span4Mux_v
    port map (
            O => \N__49605\,
            I => \N__49515\
        );

    \I__11417\ : Span4Mux_v
    port map (
            O => \N__49602\,
            I => \N__49506\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__49599\,
            I => \N__49506\
        );

    \I__11415\ : LocalMux
    port map (
            O => \N__49596\,
            I => \N__49506\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__49593\,
            I => \N__49506\
        );

    \I__11413\ : InMux
    port map (
            O => \N__49592\,
            I => \N__49503\
        );

    \I__11412\ : InMux
    port map (
            O => \N__49591\,
            I => \N__49500\
        );

    \I__11411\ : InMux
    port map (
            O => \N__49590\,
            I => \N__49497\
        );

    \I__11410\ : Span4Mux_h
    port map (
            O => \N__49587\,
            I => \N__49493\
        );

    \I__11409\ : Span4Mux_h
    port map (
            O => \N__49582\,
            I => \N__49486\
        );

    \I__11408\ : Span4Mux_h
    port map (
            O => \N__49579\,
            I => \N__49486\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__49576\,
            I => \N__49486\
        );

    \I__11406\ : InMux
    port map (
            O => \N__49575\,
            I => \N__49483\
        );

    \I__11405\ : InMux
    port map (
            O => \N__49574\,
            I => \N__49480\
        );

    \I__11404\ : InMux
    port map (
            O => \N__49573\,
            I => \N__49477\
        );

    \I__11403\ : InMux
    port map (
            O => \N__49572\,
            I => \N__49474\
        );

    \I__11402\ : InMux
    port map (
            O => \N__49571\,
            I => \N__49471\
        );

    \I__11401\ : Span4Mux_h
    port map (
            O => \N__49568\,
            I => \N__49464\
        );

    \I__11400\ : Span4Mux_v
    port map (
            O => \N__49555\,
            I => \N__49464\
        );

    \I__11399\ : LocalMux
    port map (
            O => \N__49552\,
            I => \N__49464\
        );

    \I__11398\ : Span4Mux_h
    port map (
            O => \N__49549\,
            I => \N__49459\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__49546\,
            I => \N__49459\
        );

    \I__11396\ : Span4Mux_v
    port map (
            O => \N__49533\,
            I => \N__49454\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__49530\,
            I => \N__49454\
        );

    \I__11394\ : Span4Mux_v
    port map (
            O => \N__49527\,
            I => \N__49445\
        );

    \I__11393\ : LocalMux
    port map (
            O => \N__49524\,
            I => \N__49445\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__49521\,
            I => \N__49445\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__49518\,
            I => \N__49445\
        );

    \I__11390\ : Span4Mux_h
    port map (
            O => \N__49515\,
            I => \N__49434\
        );

    \I__11389\ : Span4Mux_v
    port map (
            O => \N__49506\,
            I => \N__49434\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__49503\,
            I => \N__49434\
        );

    \I__11387\ : LocalMux
    port map (
            O => \N__49500\,
            I => \N__49434\
        );

    \I__11386\ : LocalMux
    port map (
            O => \N__49497\,
            I => \N__49434\
        );

    \I__11385\ : InMux
    port map (
            O => \N__49496\,
            I => \N__49431\
        );

    \I__11384\ : Sp12to4
    port map (
            O => \N__49493\,
            I => \N__49416\
        );

    \I__11383\ : Sp12to4
    port map (
            O => \N__49486\,
            I => \N__49416\
        );

    \I__11382\ : LocalMux
    port map (
            O => \N__49483\,
            I => \N__49416\
        );

    \I__11381\ : LocalMux
    port map (
            O => \N__49480\,
            I => \N__49416\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__49477\,
            I => \N__49416\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__49474\,
            I => \N__49416\
        );

    \I__11378\ : LocalMux
    port map (
            O => \N__49471\,
            I => \N__49416\
        );

    \I__11377\ : Span4Mux_h
    port map (
            O => \N__49464\,
            I => \N__49412\
        );

    \I__11376\ : Span4Mux_v
    port map (
            O => \N__49459\,
            I => \N__49405\
        );

    \I__11375\ : Span4Mux_h
    port map (
            O => \N__49454\,
            I => \N__49405\
        );

    \I__11374\ : Span4Mux_v
    port map (
            O => \N__49445\,
            I => \N__49405\
        );

    \I__11373\ : Span4Mux_v
    port map (
            O => \N__49434\,
            I => \N__49400\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__49431\,
            I => \N__49400\
        );

    \I__11371\ : Span12Mux_v
    port map (
            O => \N__49416\,
            I => \N__49397\
        );

    \I__11370\ : InMux
    port map (
            O => \N__49415\,
            I => \N__49394\
        );

    \I__11369\ : Odrv4
    port map (
            O => \N__49412\,
            I => spi_data_mosi_3
        );

    \I__11368\ : Odrv4
    port map (
            O => \N__49405\,
            I => spi_data_mosi_3
        );

    \I__11367\ : Odrv4
    port map (
            O => \N__49400\,
            I => spi_data_mosi_3
        );

    \I__11366\ : Odrv12
    port map (
            O => \N__49397\,
            I => spi_data_mosi_3
        );

    \I__11365\ : LocalMux
    port map (
            O => \N__49394\,
            I => spi_data_mosi_3
        );

    \I__11364\ : InMux
    port map (
            O => \N__49383\,
            I => \N__49380\
        );

    \I__11363\ : LocalMux
    port map (
            O => \N__49380\,
            I => \N__49377\
        );

    \I__11362\ : Span4Mux_h
    port map (
            O => \N__49377\,
            I => \N__49374\
        );

    \I__11361\ : Span4Mux_h
    port map (
            O => \N__49374\,
            I => \N__49371\
        );

    \I__11360\ : Odrv4
    port map (
            O => \N__49371\,
            I => \sDAC_mem_13Z0Z_3\
        );

    \I__11359\ : InMux
    port map (
            O => \N__49368\,
            I => \N__49364\
        );

    \I__11358\ : InMux
    port map (
            O => \N__49367\,
            I => \N__49351\
        );

    \I__11357\ : LocalMux
    port map (
            O => \N__49364\,
            I => \N__49348\
        );

    \I__11356\ : InMux
    port map (
            O => \N__49363\,
            I => \N__49340\
        );

    \I__11355\ : InMux
    port map (
            O => \N__49362\,
            I => \N__49337\
        );

    \I__11354\ : InMux
    port map (
            O => \N__49361\,
            I => \N__49331\
        );

    \I__11353\ : InMux
    port map (
            O => \N__49360\,
            I => \N__49328\
        );

    \I__11352\ : InMux
    port map (
            O => \N__49359\,
            I => \N__49323\
        );

    \I__11351\ : InMux
    port map (
            O => \N__49358\,
            I => \N__49319\
        );

    \I__11350\ : InMux
    port map (
            O => \N__49357\,
            I => \N__49316\
        );

    \I__11349\ : InMux
    port map (
            O => \N__49356\,
            I => \N__49313\
        );

    \I__11348\ : InMux
    port map (
            O => \N__49355\,
            I => \N__49309\
        );

    \I__11347\ : InMux
    port map (
            O => \N__49354\,
            I => \N__49302\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__49351\,
            I => \N__49297\
        );

    \I__11345\ : Span4Mux_v
    port map (
            O => \N__49348\,
            I => \N__49297\
        );

    \I__11344\ : InMux
    port map (
            O => \N__49347\,
            I => \N__49294\
        );

    \I__11343\ : InMux
    port map (
            O => \N__49346\,
            I => \N__49291\
        );

    \I__11342\ : InMux
    port map (
            O => \N__49345\,
            I => \N__49288\
        );

    \I__11341\ : InMux
    port map (
            O => \N__49344\,
            I => \N__49285\
        );

    \I__11340\ : InMux
    port map (
            O => \N__49343\,
            I => \N__49282\
        );

    \I__11339\ : LocalMux
    port map (
            O => \N__49340\,
            I => \N__49276\
        );

    \I__11338\ : LocalMux
    port map (
            O => \N__49337\,
            I => \N__49276\
        );

    \I__11337\ : InMux
    port map (
            O => \N__49336\,
            I => \N__49273\
        );

    \I__11336\ : InMux
    port map (
            O => \N__49335\,
            I => \N__49270\
        );

    \I__11335\ : InMux
    port map (
            O => \N__49334\,
            I => \N__49267\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__49331\,
            I => \N__49264\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__49328\,
            I => \N__49261\
        );

    \I__11332\ : InMux
    port map (
            O => \N__49327\,
            I => \N__49257\
        );

    \I__11331\ : InMux
    port map (
            O => \N__49326\,
            I => \N__49254\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__49323\,
            I => \N__49251\
        );

    \I__11329\ : InMux
    port map (
            O => \N__49322\,
            I => \N__49248\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__49319\,
            I => \N__49241\
        );

    \I__11327\ : LocalMux
    port map (
            O => \N__49316\,
            I => \N__49241\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__49313\,
            I => \N__49241\
        );

    \I__11325\ : InMux
    port map (
            O => \N__49312\,
            I => \N__49238\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__49309\,
            I => \N__49235\
        );

    \I__11323\ : InMux
    port map (
            O => \N__49308\,
            I => \N__49232\
        );

    \I__11322\ : InMux
    port map (
            O => \N__49307\,
            I => \N__49227\
        );

    \I__11321\ : InMux
    port map (
            O => \N__49306\,
            I => \N__49223\
        );

    \I__11320\ : InMux
    port map (
            O => \N__49305\,
            I => \N__49219\
        );

    \I__11319\ : LocalMux
    port map (
            O => \N__49302\,
            I => \N__49208\
        );

    \I__11318\ : Span4Mux_h
    port map (
            O => \N__49297\,
            I => \N__49208\
        );

    \I__11317\ : LocalMux
    port map (
            O => \N__49294\,
            I => \N__49208\
        );

    \I__11316\ : LocalMux
    port map (
            O => \N__49291\,
            I => \N__49208\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__49288\,
            I => \N__49208\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__49285\,
            I => \N__49202\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__49282\,
            I => \N__49202\
        );

    \I__11312\ : InMux
    port map (
            O => \N__49281\,
            I => \N__49199\
        );

    \I__11311\ : Span4Mux_v
    port map (
            O => \N__49276\,
            I => \N__49190\
        );

    \I__11310\ : LocalMux
    port map (
            O => \N__49273\,
            I => \N__49190\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__49270\,
            I => \N__49190\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__49267\,
            I => \N__49190\
        );

    \I__11307\ : Span4Mux_h
    port map (
            O => \N__49264\,
            I => \N__49181\
        );

    \I__11306\ : Span4Mux_v
    port map (
            O => \N__49261\,
            I => \N__49181\
        );

    \I__11305\ : InMux
    port map (
            O => \N__49260\,
            I => \N__49178\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__49257\,
            I => \N__49172\
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__49254\,
            I => \N__49172\
        );

    \I__11302\ : Span4Mux_h
    port map (
            O => \N__49251\,
            I => \N__49167\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__49248\,
            I => \N__49167\
        );

    \I__11300\ : Span4Mux_v
    port map (
            O => \N__49241\,
            I => \N__49160\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__49238\,
            I => \N__49160\
        );

    \I__11298\ : Span4Mux_v
    port map (
            O => \N__49235\,
            I => \N__49155\
        );

    \I__11297\ : LocalMux
    port map (
            O => \N__49232\,
            I => \N__49155\
        );

    \I__11296\ : InMux
    port map (
            O => \N__49231\,
            I => \N__49152\
        );

    \I__11295\ : InMux
    port map (
            O => \N__49230\,
            I => \N__49149\
        );

    \I__11294\ : LocalMux
    port map (
            O => \N__49227\,
            I => \N__49146\
        );

    \I__11293\ : InMux
    port map (
            O => \N__49226\,
            I => \N__49141\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__49223\,
            I => \N__49138\
        );

    \I__11291\ : InMux
    port map (
            O => \N__49222\,
            I => \N__49135\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__49219\,
            I => \N__49132\
        );

    \I__11289\ : Span4Mux_v
    port map (
            O => \N__49208\,
            I => \N__49126\
        );

    \I__11288\ : InMux
    port map (
            O => \N__49207\,
            I => \N__49123\
        );

    \I__11287\ : Span4Mux_v
    port map (
            O => \N__49202\,
            I => \N__49120\
        );

    \I__11286\ : LocalMux
    port map (
            O => \N__49199\,
            I => \N__49115\
        );

    \I__11285\ : Span4Mux_v
    port map (
            O => \N__49190\,
            I => \N__49115\
        );

    \I__11284\ : InMux
    port map (
            O => \N__49189\,
            I => \N__49112\
        );

    \I__11283\ : InMux
    port map (
            O => \N__49188\,
            I => \N__49106\
        );

    \I__11282\ : InMux
    port map (
            O => \N__49187\,
            I => \N__49103\
        );

    \I__11281\ : InMux
    port map (
            O => \N__49186\,
            I => \N__49100\
        );

    \I__11280\ : Span4Mux_h
    port map (
            O => \N__49181\,
            I => \N__49095\
        );

    \I__11279\ : LocalMux
    port map (
            O => \N__49178\,
            I => \N__49095\
        );

    \I__11278\ : InMux
    port map (
            O => \N__49177\,
            I => \N__49092\
        );

    \I__11277\ : Span4Mux_v
    port map (
            O => \N__49172\,
            I => \N__49088\
        );

    \I__11276\ : Span4Mux_v
    port map (
            O => \N__49167\,
            I => \N__49085\
        );

    \I__11275\ : InMux
    port map (
            O => \N__49166\,
            I => \N__49082\
        );

    \I__11274\ : InMux
    port map (
            O => \N__49165\,
            I => \N__49079\
        );

    \I__11273\ : Span4Mux_v
    port map (
            O => \N__49160\,
            I => \N__49068\
        );

    \I__11272\ : Span4Mux_h
    port map (
            O => \N__49155\,
            I => \N__49068\
        );

    \I__11271\ : LocalMux
    port map (
            O => \N__49152\,
            I => \N__49068\
        );

    \I__11270\ : LocalMux
    port map (
            O => \N__49149\,
            I => \N__49063\
        );

    \I__11269\ : Span4Mux_v
    port map (
            O => \N__49146\,
            I => \N__49063\
        );

    \I__11268\ : InMux
    port map (
            O => \N__49145\,
            I => \N__49060\
        );

    \I__11267\ : InMux
    port map (
            O => \N__49144\,
            I => \N__49057\
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__49141\,
            I => \N__49052\
        );

    \I__11265\ : Span4Mux_h
    port map (
            O => \N__49138\,
            I => \N__49052\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__49135\,
            I => \N__49047\
        );

    \I__11263\ : Span4Mux_v
    port map (
            O => \N__49132\,
            I => \N__49047\
        );

    \I__11262\ : InMux
    port map (
            O => \N__49131\,
            I => \N__49044\
        );

    \I__11261\ : InMux
    port map (
            O => \N__49130\,
            I => \N__49041\
        );

    \I__11260\ : InMux
    port map (
            O => \N__49129\,
            I => \N__49038\
        );

    \I__11259\ : Sp12to4
    port map (
            O => \N__49126\,
            I => \N__49035\
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__49123\,
            I => \N__49028\
        );

    \I__11257\ : Sp12to4
    port map (
            O => \N__49120\,
            I => \N__49028\
        );

    \I__11256\ : Sp12to4
    port map (
            O => \N__49115\,
            I => \N__49028\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__49112\,
            I => \N__49025\
        );

    \I__11254\ : InMux
    port map (
            O => \N__49111\,
            I => \N__49022\
        );

    \I__11253\ : InMux
    port map (
            O => \N__49110\,
            I => \N__49019\
        );

    \I__11252\ : InMux
    port map (
            O => \N__49109\,
            I => \N__49016\
        );

    \I__11251\ : LocalMux
    port map (
            O => \N__49106\,
            I => \N__49009\
        );

    \I__11250\ : LocalMux
    port map (
            O => \N__49103\,
            I => \N__49009\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__49100\,
            I => \N__49009\
        );

    \I__11248\ : Span4Mux_v
    port map (
            O => \N__49095\,
            I => \N__49004\
        );

    \I__11247\ : LocalMux
    port map (
            O => \N__49092\,
            I => \N__49004\
        );

    \I__11246\ : InMux
    port map (
            O => \N__49091\,
            I => \N__49001\
        );

    \I__11245\ : Sp12to4
    port map (
            O => \N__49088\,
            I => \N__48998\
        );

    \I__11244\ : Sp12to4
    port map (
            O => \N__49085\,
            I => \N__48993\
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__49082\,
            I => \N__48993\
        );

    \I__11242\ : LocalMux
    port map (
            O => \N__49079\,
            I => \N__48990\
        );

    \I__11241\ : InMux
    port map (
            O => \N__49078\,
            I => \N__48985\
        );

    \I__11240\ : InMux
    port map (
            O => \N__49077\,
            I => \N__48982\
        );

    \I__11239\ : InMux
    port map (
            O => \N__49076\,
            I => \N__48979\
        );

    \I__11238\ : InMux
    port map (
            O => \N__49075\,
            I => \N__48976\
        );

    \I__11237\ : Span4Mux_v
    port map (
            O => \N__49068\,
            I => \N__48973\
        );

    \I__11236\ : Span4Mux_h
    port map (
            O => \N__49063\,
            I => \N__48962\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__49060\,
            I => \N__48962\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__49057\,
            I => \N__48962\
        );

    \I__11233\ : Span4Mux_v
    port map (
            O => \N__49052\,
            I => \N__48962\
        );

    \I__11232\ : Span4Mux_h
    port map (
            O => \N__49047\,
            I => \N__48962\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__49044\,
            I => \N__48949\
        );

    \I__11230\ : LocalMux
    port map (
            O => \N__49041\,
            I => \N__48949\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__49038\,
            I => \N__48949\
        );

    \I__11228\ : Span12Mux_h
    port map (
            O => \N__49035\,
            I => \N__48949\
        );

    \I__11227\ : Span12Mux_h
    port map (
            O => \N__49028\,
            I => \N__48949\
        );

    \I__11226\ : Span12Mux_h
    port map (
            O => \N__49025\,
            I => \N__48949\
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__49022\,
            I => \N__48930\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__49019\,
            I => \N__48930\
        );

    \I__11223\ : LocalMux
    port map (
            O => \N__49016\,
            I => \N__48930\
        );

    \I__11222\ : Sp12to4
    port map (
            O => \N__49009\,
            I => \N__48930\
        );

    \I__11221\ : Sp12to4
    port map (
            O => \N__49004\,
            I => \N__48930\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__49001\,
            I => \N__48930\
        );

    \I__11219\ : Span12Mux_s11_v
    port map (
            O => \N__48998\,
            I => \N__48930\
        );

    \I__11218\ : Span12Mux_h
    port map (
            O => \N__48993\,
            I => \N__48930\
        );

    \I__11217\ : Span12Mux_h
    port map (
            O => \N__48990\,
            I => \N__48930\
        );

    \I__11216\ : InMux
    port map (
            O => \N__48989\,
            I => \N__48927\
        );

    \I__11215\ : InMux
    port map (
            O => \N__48988\,
            I => \N__48924\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__48985\,
            I => \N__48911\
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__48982\,
            I => \N__48911\
        );

    \I__11212\ : LocalMux
    port map (
            O => \N__48979\,
            I => \N__48911\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__48976\,
            I => \N__48911\
        );

    \I__11210\ : Span4Mux_h
    port map (
            O => \N__48973\,
            I => \N__48911\
        );

    \I__11209\ : Span4Mux_v
    port map (
            O => \N__48962\,
            I => \N__48911\
        );

    \I__11208\ : Span12Mux_v
    port map (
            O => \N__48949\,
            I => \N__48907\
        );

    \I__11207\ : Span12Mux_v
    port map (
            O => \N__48930\,
            I => \N__48904\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__48927\,
            I => \N__48897\
        );

    \I__11205\ : LocalMux
    port map (
            O => \N__48924\,
            I => \N__48897\
        );

    \I__11204\ : Span4Mux_v
    port map (
            O => \N__48911\,
            I => \N__48897\
        );

    \I__11203\ : InMux
    port map (
            O => \N__48910\,
            I => \N__48894\
        );

    \I__11202\ : Odrv12
    port map (
            O => \N__48907\,
            I => spi_data_mosi_4
        );

    \I__11201\ : Odrv12
    port map (
            O => \N__48904\,
            I => spi_data_mosi_4
        );

    \I__11200\ : Odrv4
    port map (
            O => \N__48897\,
            I => spi_data_mosi_4
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__48894\,
            I => spi_data_mosi_4
        );

    \I__11198\ : InMux
    port map (
            O => \N__48885\,
            I => \N__48882\
        );

    \I__11197\ : LocalMux
    port map (
            O => \N__48882\,
            I => \N__48879\
        );

    \I__11196\ : Span4Mux_h
    port map (
            O => \N__48879\,
            I => \N__48876\
        );

    \I__11195\ : Odrv4
    port map (
            O => \N__48876\,
            I => \sDAC_mem_13Z0Z_4\
        );

    \I__11194\ : InMux
    port map (
            O => \N__48873\,
            I => \N__48870\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__48870\,
            I => \sDAC_mem_13Z0Z_7\
        );

    \I__11192\ : CEMux
    port map (
            O => \N__48867\,
            I => \N__48863\
        );

    \I__11191\ : CEMux
    port map (
            O => \N__48866\,
            I => \N__48860\
        );

    \I__11190\ : LocalMux
    port map (
            O => \N__48863\,
            I => \N__48857\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__48860\,
            I => \N__48854\
        );

    \I__11188\ : Span4Mux_v
    port map (
            O => \N__48857\,
            I => \N__48851\
        );

    \I__11187\ : Span4Mux_v
    port map (
            O => \N__48854\,
            I => \N__48848\
        );

    \I__11186\ : Odrv4
    port map (
            O => \N__48851\,
            I => \sDAC_mem_13_1_sqmuxa\
        );

    \I__11185\ : Odrv4
    port map (
            O => \N__48848\,
            I => \sDAC_mem_13_1_sqmuxa\
        );

    \I__11184\ : InMux
    port map (
            O => \N__48843\,
            I => \N__48838\
        );

    \I__11183\ : InMux
    port map (
            O => \N__48842\,
            I => \N__48835\
        );

    \I__11182\ : InMux
    port map (
            O => \N__48841\,
            I => \N__48827\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__48838\,
            I => \N__48822\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__48835\,
            I => \N__48822\
        );

    \I__11179\ : InMux
    port map (
            O => \N__48834\,
            I => \N__48819\
        );

    \I__11178\ : InMux
    port map (
            O => \N__48833\,
            I => \N__48813\
        );

    \I__11177\ : InMux
    port map (
            O => \N__48832\,
            I => \N__48809\
        );

    \I__11176\ : InMux
    port map (
            O => \N__48831\,
            I => \N__48805\
        );

    \I__11175\ : InMux
    port map (
            O => \N__48830\,
            I => \N__48802\
        );

    \I__11174\ : LocalMux
    port map (
            O => \N__48827\,
            I => \N__48790\
        );

    \I__11173\ : Span4Mux_h
    port map (
            O => \N__48822\,
            I => \N__48790\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__48819\,
            I => \N__48790\
        );

    \I__11171\ : InMux
    port map (
            O => \N__48818\,
            I => \N__48787\
        );

    \I__11170\ : InMux
    port map (
            O => \N__48817\,
            I => \N__48783\
        );

    \I__11169\ : InMux
    port map (
            O => \N__48816\,
            I => \N__48780\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__48813\,
            I => \N__48773\
        );

    \I__11167\ : InMux
    port map (
            O => \N__48812\,
            I => \N__48770\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__48809\,
            I => \N__48765\
        );

    \I__11165\ : InMux
    port map (
            O => \N__48808\,
            I => \N__48762\
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__48805\,
            I => \N__48757\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__48802\,
            I => \N__48757\
        );

    \I__11162\ : InMux
    port map (
            O => \N__48801\,
            I => \N__48754\
        );

    \I__11161\ : InMux
    port map (
            O => \N__48800\,
            I => \N__48751\
        );

    \I__11160\ : InMux
    port map (
            O => \N__48799\,
            I => \N__48748\
        );

    \I__11159\ : InMux
    port map (
            O => \N__48798\,
            I => \N__48733\
        );

    \I__11158\ : InMux
    port map (
            O => \N__48797\,
            I => \N__48730\
        );

    \I__11157\ : Span4Mux_v
    port map (
            O => \N__48790\,
            I => \N__48723\
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__48787\,
            I => \N__48723\
        );

    \I__11155\ : InMux
    port map (
            O => \N__48786\,
            I => \N__48720\
        );

    \I__11154\ : LocalMux
    port map (
            O => \N__48783\,
            I => \N__48713\
        );

    \I__11153\ : LocalMux
    port map (
            O => \N__48780\,
            I => \N__48713\
        );

    \I__11152\ : InMux
    port map (
            O => \N__48779\,
            I => \N__48710\
        );

    \I__11151\ : InMux
    port map (
            O => \N__48778\,
            I => \N__48707\
        );

    \I__11150\ : InMux
    port map (
            O => \N__48777\,
            I => \N__48702\
        );

    \I__11149\ : InMux
    port map (
            O => \N__48776\,
            I => \N__48699\
        );

    \I__11148\ : Span4Mux_v
    port map (
            O => \N__48773\,
            I => \N__48694\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__48770\,
            I => \N__48694\
        );

    \I__11146\ : InMux
    port map (
            O => \N__48769\,
            I => \N__48691\
        );

    \I__11145\ : InMux
    port map (
            O => \N__48768\,
            I => \N__48688\
        );

    \I__11144\ : Span4Mux_h
    port map (
            O => \N__48765\,
            I => \N__48683\
        );

    \I__11143\ : LocalMux
    port map (
            O => \N__48762\,
            I => \N__48683\
        );

    \I__11142\ : Span4Mux_v
    port map (
            O => \N__48757\,
            I => \N__48678\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__48754\,
            I => \N__48678\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__48751\,
            I => \N__48673\
        );

    \I__11139\ : LocalMux
    port map (
            O => \N__48748\,
            I => \N__48673\
        );

    \I__11138\ : InMux
    port map (
            O => \N__48747\,
            I => \N__48664\
        );

    \I__11137\ : InMux
    port map (
            O => \N__48746\,
            I => \N__48661\
        );

    \I__11136\ : InMux
    port map (
            O => \N__48745\,
            I => \N__48658\
        );

    \I__11135\ : InMux
    port map (
            O => \N__48744\,
            I => \N__48655\
        );

    \I__11134\ : InMux
    port map (
            O => \N__48743\,
            I => \N__48652\
        );

    \I__11133\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48649\
        );

    \I__11132\ : InMux
    port map (
            O => \N__48741\,
            I => \N__48646\
        );

    \I__11131\ : InMux
    port map (
            O => \N__48740\,
            I => \N__48643\
        );

    \I__11130\ : InMux
    port map (
            O => \N__48739\,
            I => \N__48640\
        );

    \I__11129\ : InMux
    port map (
            O => \N__48738\,
            I => \N__48637\
        );

    \I__11128\ : InMux
    port map (
            O => \N__48737\,
            I => \N__48634\
        );

    \I__11127\ : InMux
    port map (
            O => \N__48736\,
            I => \N__48630\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__48733\,
            I => \N__48627\
        );

    \I__11125\ : LocalMux
    port map (
            O => \N__48730\,
            I => \N__48624\
        );

    \I__11124\ : InMux
    port map (
            O => \N__48729\,
            I => \N__48621\
        );

    \I__11123\ : InMux
    port map (
            O => \N__48728\,
            I => \N__48618\
        );

    \I__11122\ : Span4Mux_v
    port map (
            O => \N__48723\,
            I => \N__48613\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__48720\,
            I => \N__48613\
        );

    \I__11120\ : InMux
    port map (
            O => \N__48719\,
            I => \N__48610\
        );

    \I__11119\ : InMux
    port map (
            O => \N__48718\,
            I => \N__48607\
        );

    \I__11118\ : Span4Mux_h
    port map (
            O => \N__48713\,
            I => \N__48600\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__48710\,
            I => \N__48600\
        );

    \I__11116\ : LocalMux
    port map (
            O => \N__48707\,
            I => \N__48600\
        );

    \I__11115\ : InMux
    port map (
            O => \N__48706\,
            I => \N__48594\
        );

    \I__11114\ : InMux
    port map (
            O => \N__48705\,
            I => \N__48589\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__48702\,
            I => \N__48586\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__48699\,
            I => \N__48583\
        );

    \I__11111\ : Span4Mux_h
    port map (
            O => \N__48694\,
            I => \N__48580\
        );

    \I__11110\ : LocalMux
    port map (
            O => \N__48691\,
            I => \N__48577\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__48688\,
            I => \N__48572\
        );

    \I__11108\ : Span4Mux_v
    port map (
            O => \N__48683\,
            I => \N__48569\
        );

    \I__11107\ : Span4Mux_v
    port map (
            O => \N__48678\,
            I => \N__48564\
        );

    \I__11106\ : Span4Mux_h
    port map (
            O => \N__48673\,
            I => \N__48564\
        );

    \I__11105\ : CascadeMux
    port map (
            O => \N__48672\,
            I => \N__48561\
        );

    \I__11104\ : InMux
    port map (
            O => \N__48671\,
            I => \N__48558\
        );

    \I__11103\ : InMux
    port map (
            O => \N__48670\,
            I => \N__48555\
        );

    \I__11102\ : InMux
    port map (
            O => \N__48669\,
            I => \N__48552\
        );

    \I__11101\ : InMux
    port map (
            O => \N__48668\,
            I => \N__48549\
        );

    \I__11100\ : InMux
    port map (
            O => \N__48667\,
            I => \N__48546\
        );

    \I__11099\ : LocalMux
    port map (
            O => \N__48664\,
            I => \N__48540\
        );

    \I__11098\ : LocalMux
    port map (
            O => \N__48661\,
            I => \N__48540\
        );

    \I__11097\ : LocalMux
    port map (
            O => \N__48658\,
            I => \N__48531\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__48655\,
            I => \N__48531\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__48652\,
            I => \N__48531\
        );

    \I__11094\ : LocalMux
    port map (
            O => \N__48649\,
            I => \N__48531\
        );

    \I__11093\ : LocalMux
    port map (
            O => \N__48646\,
            I => \N__48520\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__48643\,
            I => \N__48520\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__48640\,
            I => \N__48520\
        );

    \I__11090\ : LocalMux
    port map (
            O => \N__48637\,
            I => \N__48520\
        );

    \I__11089\ : LocalMux
    port map (
            O => \N__48634\,
            I => \N__48520\
        );

    \I__11088\ : InMux
    port map (
            O => \N__48633\,
            I => \N__48517\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__48630\,
            I => \N__48512\
        );

    \I__11086\ : Span4Mux_h
    port map (
            O => \N__48627\,
            I => \N__48512\
        );

    \I__11085\ : Span4Mux_h
    port map (
            O => \N__48624\,
            I => \N__48507\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__48621\,
            I => \N__48507\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__48618\,
            I => \N__48502\
        );

    \I__11082\ : Span4Mux_h
    port map (
            O => \N__48613\,
            I => \N__48502\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__48610\,
            I => \N__48495\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__48607\,
            I => \N__48495\
        );

    \I__11079\ : Span4Mux_h
    port map (
            O => \N__48600\,
            I => \N__48495\
        );

    \I__11078\ : InMux
    port map (
            O => \N__48599\,
            I => \N__48492\
        );

    \I__11077\ : InMux
    port map (
            O => \N__48598\,
            I => \N__48489\
        );

    \I__11076\ : InMux
    port map (
            O => \N__48597\,
            I => \N__48486\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__48594\,
            I => \N__48483\
        );

    \I__11074\ : InMux
    port map (
            O => \N__48593\,
            I => \N__48480\
        );

    \I__11073\ : InMux
    port map (
            O => \N__48592\,
            I => \N__48477\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__48589\,
            I => \N__48474\
        );

    \I__11071\ : Span4Mux_h
    port map (
            O => \N__48586\,
            I => \N__48465\
        );

    \I__11070\ : Span4Mux_v
    port map (
            O => \N__48583\,
            I => \N__48465\
        );

    \I__11069\ : Span4Mux_h
    port map (
            O => \N__48580\,
            I => \N__48465\
        );

    \I__11068\ : Span4Mux_h
    port map (
            O => \N__48577\,
            I => \N__48465\
        );

    \I__11067\ : InMux
    port map (
            O => \N__48576\,
            I => \N__48462\
        );

    \I__11066\ : InMux
    port map (
            O => \N__48575\,
            I => \N__48459\
        );

    \I__11065\ : Span4Mux_h
    port map (
            O => \N__48572\,
            I => \N__48456\
        );

    \I__11064\ : Sp12to4
    port map (
            O => \N__48569\,
            I => \N__48453\
        );

    \I__11063\ : Span4Mux_h
    port map (
            O => \N__48564\,
            I => \N__48450\
        );

    \I__11062\ : InMux
    port map (
            O => \N__48561\,
            I => \N__48447\
        );

    \I__11061\ : LocalMux
    port map (
            O => \N__48558\,
            I => \N__48436\
        );

    \I__11060\ : LocalMux
    port map (
            O => \N__48555\,
            I => \N__48436\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__48552\,
            I => \N__48436\
        );

    \I__11058\ : LocalMux
    port map (
            O => \N__48549\,
            I => \N__48436\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__48546\,
            I => \N__48436\
        );

    \I__11056\ : InMux
    port map (
            O => \N__48545\,
            I => \N__48433\
        );

    \I__11055\ : Span4Mux_v
    port map (
            O => \N__48540\,
            I => \N__48428\
        );

    \I__11054\ : Span4Mux_v
    port map (
            O => \N__48531\,
            I => \N__48428\
        );

    \I__11053\ : Span4Mux_v
    port map (
            O => \N__48520\,
            I => \N__48425\
        );

    \I__11052\ : LocalMux
    port map (
            O => \N__48517\,
            I => \N__48420\
        );

    \I__11051\ : Sp12to4
    port map (
            O => \N__48512\,
            I => \N__48420\
        );

    \I__11050\ : Sp12to4
    port map (
            O => \N__48507\,
            I => \N__48413\
        );

    \I__11049\ : Sp12to4
    port map (
            O => \N__48502\,
            I => \N__48413\
        );

    \I__11048\ : Sp12to4
    port map (
            O => \N__48495\,
            I => \N__48413\
        );

    \I__11047\ : LocalMux
    port map (
            O => \N__48492\,
            I => \N__48404\
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__48489\,
            I => \N__48404\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__48486\,
            I => \N__48404\
        );

    \I__11044\ : Span4Mux_h
    port map (
            O => \N__48483\,
            I => \N__48404\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__48480\,
            I => \N__48401\
        );

    \I__11042\ : LocalMux
    port map (
            O => \N__48477\,
            I => \N__48394\
        );

    \I__11041\ : Span4Mux_v
    port map (
            O => \N__48474\,
            I => \N__48394\
        );

    \I__11040\ : Span4Mux_h
    port map (
            O => \N__48465\,
            I => \N__48394\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__48462\,
            I => \N__48381\
        );

    \I__11038\ : LocalMux
    port map (
            O => \N__48459\,
            I => \N__48381\
        );

    \I__11037\ : Sp12to4
    port map (
            O => \N__48456\,
            I => \N__48381\
        );

    \I__11036\ : Span12Mux_h
    port map (
            O => \N__48453\,
            I => \N__48381\
        );

    \I__11035\ : Sp12to4
    port map (
            O => \N__48450\,
            I => \N__48381\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__48447\,
            I => \N__48381\
        );

    \I__11033\ : Span12Mux_v
    port map (
            O => \N__48436\,
            I => \N__48378\
        );

    \I__11032\ : LocalMux
    port map (
            O => \N__48433\,
            I => \N__48367\
        );

    \I__11031\ : Sp12to4
    port map (
            O => \N__48428\,
            I => \N__48367\
        );

    \I__11030\ : Sp12to4
    port map (
            O => \N__48425\,
            I => \N__48367\
        );

    \I__11029\ : Span12Mux_v
    port map (
            O => \N__48420\,
            I => \N__48367\
        );

    \I__11028\ : Span12Mux_v
    port map (
            O => \N__48413\,
            I => \N__48367\
        );

    \I__11027\ : Sp12to4
    port map (
            O => \N__48404\,
            I => \N__48358\
        );

    \I__11026\ : Span12Mux_h
    port map (
            O => \N__48401\,
            I => \N__48358\
        );

    \I__11025\ : Sp12to4
    port map (
            O => \N__48394\,
            I => \N__48358\
        );

    \I__11024\ : Span12Mux_v
    port map (
            O => \N__48381\,
            I => \N__48358\
        );

    \I__11023\ : Odrv12
    port map (
            O => \N__48378\,
            I => spi_data_mosi_7
        );

    \I__11022\ : Odrv12
    port map (
            O => \N__48367\,
            I => spi_data_mosi_7
        );

    \I__11021\ : Odrv12
    port map (
            O => \N__48358\,
            I => spi_data_mosi_7
        );

    \I__11020\ : InMux
    port map (
            O => \N__48351\,
            I => \N__48348\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__48348\,
            I => \N__48345\
        );

    \I__11018\ : Odrv4
    port map (
            O => \N__48345\,
            I => \sDAC_mem_12Z0Z_7\
        );

    \I__11017\ : InMux
    port map (
            O => \N__48342\,
            I => \N__48333\
        );

    \I__11016\ : InMux
    port map (
            O => \N__48341\,
            I => \N__48326\
        );

    \I__11015\ : InMux
    port map (
            O => \N__48340\,
            I => \N__48321\
        );

    \I__11014\ : InMux
    port map (
            O => \N__48339\,
            I => \N__48318\
        );

    \I__11013\ : InMux
    port map (
            O => \N__48338\,
            I => \N__48315\
        );

    \I__11012\ : InMux
    port map (
            O => \N__48337\,
            I => \N__48312\
        );

    \I__11011\ : InMux
    port map (
            O => \N__48336\,
            I => \N__48307\
        );

    \I__11010\ : LocalMux
    port map (
            O => \N__48333\,
            I => \N__48300\
        );

    \I__11009\ : InMux
    port map (
            O => \N__48332\,
            I => \N__48297\
        );

    \I__11008\ : InMux
    port map (
            O => \N__48331\,
            I => \N__48294\
        );

    \I__11007\ : InMux
    port map (
            O => \N__48330\,
            I => \N__48291\
        );

    \I__11006\ : InMux
    port map (
            O => \N__48329\,
            I => \N__48288\
        );

    \I__11005\ : LocalMux
    port map (
            O => \N__48326\,
            I => \N__48285\
        );

    \I__11004\ : InMux
    port map (
            O => \N__48325\,
            I => \N__48282\
        );

    \I__11003\ : InMux
    port map (
            O => \N__48324\,
            I => \N__48275\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__48321\,
            I => \N__48269\
        );

    \I__11001\ : LocalMux
    port map (
            O => \N__48318\,
            I => \N__48262\
        );

    \I__11000\ : LocalMux
    port map (
            O => \N__48315\,
            I => \N__48262\
        );

    \I__10999\ : LocalMux
    port map (
            O => \N__48312\,
            I => \N__48262\
        );

    \I__10998\ : InMux
    port map (
            O => \N__48311\,
            I => \N__48259\
        );

    \I__10997\ : InMux
    port map (
            O => \N__48310\,
            I => \N__48256\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__48307\,
            I => \N__48251\
        );

    \I__10995\ : InMux
    port map (
            O => \N__48306\,
            I => \N__48248\
        );

    \I__10994\ : InMux
    port map (
            O => \N__48305\,
            I => \N__48245\
        );

    \I__10993\ : InMux
    port map (
            O => \N__48304\,
            I => \N__48241\
        );

    \I__10992\ : InMux
    port map (
            O => \N__48303\,
            I => \N__48238\
        );

    \I__10991\ : Span4Mux_v
    port map (
            O => \N__48300\,
            I => \N__48220\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__48297\,
            I => \N__48220\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__48294\,
            I => \N__48220\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__48291\,
            I => \N__48215\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__48288\,
            I => \N__48215\
        );

    \I__10986\ : Span4Mux_v
    port map (
            O => \N__48285\,
            I => \N__48205\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__48282\,
            I => \N__48205\
        );

    \I__10984\ : InMux
    port map (
            O => \N__48281\,
            I => \N__48202\
        );

    \I__10983\ : InMux
    port map (
            O => \N__48280\,
            I => \N__48199\
        );

    \I__10982\ : InMux
    port map (
            O => \N__48279\,
            I => \N__48196\
        );

    \I__10981\ : InMux
    port map (
            O => \N__48278\,
            I => \N__48193\
        );

    \I__10980\ : LocalMux
    port map (
            O => \N__48275\,
            I => \N__48186\
        );

    \I__10979\ : InMux
    port map (
            O => \N__48274\,
            I => \N__48183\
        );

    \I__10978\ : InMux
    port map (
            O => \N__48273\,
            I => \N__48180\
        );

    \I__10977\ : InMux
    port map (
            O => \N__48272\,
            I => \N__48177\
        );

    \I__10976\ : Span4Mux_h
    port map (
            O => \N__48269\,
            I => \N__48168\
        );

    \I__10975\ : Span4Mux_v
    port map (
            O => \N__48262\,
            I => \N__48168\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__48259\,
            I => \N__48168\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__48256\,
            I => \N__48168\
        );

    \I__10972\ : InMux
    port map (
            O => \N__48255\,
            I => \N__48165\
        );

    \I__10971\ : InMux
    port map (
            O => \N__48254\,
            I => \N__48162\
        );

    \I__10970\ : Span4Mux_v
    port map (
            O => \N__48251\,
            I => \N__48154\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__48248\,
            I => \N__48154\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__48245\,
            I => \N__48150\
        );

    \I__10967\ : InMux
    port map (
            O => \N__48244\,
            I => \N__48147\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__48241\,
            I => \N__48143\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__48238\,
            I => \N__48140\
        );

    \I__10964\ : InMux
    port map (
            O => \N__48237\,
            I => \N__48137\
        );

    \I__10963\ : InMux
    port map (
            O => \N__48236\,
            I => \N__48134\
        );

    \I__10962\ : InMux
    port map (
            O => \N__48235\,
            I => \N__48131\
        );

    \I__10961\ : InMux
    port map (
            O => \N__48234\,
            I => \N__48128\
        );

    \I__10960\ : InMux
    port map (
            O => \N__48233\,
            I => \N__48125\
        );

    \I__10959\ : InMux
    port map (
            O => \N__48232\,
            I => \N__48121\
        );

    \I__10958\ : InMux
    port map (
            O => \N__48231\,
            I => \N__48118\
        );

    \I__10957\ : InMux
    port map (
            O => \N__48230\,
            I => \N__48115\
        );

    \I__10956\ : InMux
    port map (
            O => \N__48229\,
            I => \N__48112\
        );

    \I__10955\ : InMux
    port map (
            O => \N__48228\,
            I => \N__48109\
        );

    \I__10954\ : InMux
    port map (
            O => \N__48227\,
            I => \N__48106\
        );

    \I__10953\ : Span4Mux_v
    port map (
            O => \N__48220\,
            I => \N__48101\
        );

    \I__10952\ : Span4Mux_h
    port map (
            O => \N__48215\,
            I => \N__48101\
        );

    \I__10951\ : InMux
    port map (
            O => \N__48214\,
            I => \N__48098\
        );

    \I__10950\ : InMux
    port map (
            O => \N__48213\,
            I => \N__48095\
        );

    \I__10949\ : InMux
    port map (
            O => \N__48212\,
            I => \N__48092\
        );

    \I__10948\ : InMux
    port map (
            O => \N__48211\,
            I => \N__48089\
        );

    \I__10947\ : InMux
    port map (
            O => \N__48210\,
            I => \N__48086\
        );

    \I__10946\ : Span4Mux_v
    port map (
            O => \N__48205\,
            I => \N__48075\
        );

    \I__10945\ : LocalMux
    port map (
            O => \N__48202\,
            I => \N__48075\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__48199\,
            I => \N__48075\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__48196\,
            I => \N__48075\
        );

    \I__10942\ : LocalMux
    port map (
            O => \N__48193\,
            I => \N__48075\
        );

    \I__10941\ : InMux
    port map (
            O => \N__48192\,
            I => \N__48072\
        );

    \I__10940\ : InMux
    port map (
            O => \N__48191\,
            I => \N__48069\
        );

    \I__10939\ : InMux
    port map (
            O => \N__48190\,
            I => \N__48066\
        );

    \I__10938\ : InMux
    port map (
            O => \N__48189\,
            I => \N__48063\
        );

    \I__10937\ : Span4Mux_h
    port map (
            O => \N__48186\,
            I => \N__48053\
        );

    \I__10936\ : LocalMux
    port map (
            O => \N__48183\,
            I => \N__48053\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__48180\,
            I => \N__48053\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__48177\,
            I => \N__48053\
        );

    \I__10933\ : Span4Mux_v
    port map (
            O => \N__48168\,
            I => \N__48046\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__48165\,
            I => \N__48046\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__48162\,
            I => \N__48046\
        );

    \I__10930\ : InMux
    port map (
            O => \N__48161\,
            I => \N__48043\
        );

    \I__10929\ : InMux
    port map (
            O => \N__48160\,
            I => \N__48040\
        );

    \I__10928\ : InMux
    port map (
            O => \N__48159\,
            I => \N__48037\
        );

    \I__10927\ : Span4Mux_v
    port map (
            O => \N__48154\,
            I => \N__48034\
        );

    \I__10926\ : InMux
    port map (
            O => \N__48153\,
            I => \N__48031\
        );

    \I__10925\ : Span4Mux_h
    port map (
            O => \N__48150\,
            I => \N__48026\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__48147\,
            I => \N__48026\
        );

    \I__10923\ : InMux
    port map (
            O => \N__48146\,
            I => \N__48023\
        );

    \I__10922\ : Span4Mux_v
    port map (
            O => \N__48143\,
            I => \N__48014\
        );

    \I__10921\ : Span4Mux_v
    port map (
            O => \N__48140\,
            I => \N__48014\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__48137\,
            I => \N__48014\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__48134\,
            I => \N__48014\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__48131\,
            I => \N__48007\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__48128\,
            I => \N__48007\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__48125\,
            I => \N__48007\
        );

    \I__10915\ : InMux
    port map (
            O => \N__48124\,
            I => \N__48004\
        );

    \I__10914\ : LocalMux
    port map (
            O => \N__48121\,
            I => \N__48001\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__48118\,
            I => \N__47996\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__48115\,
            I => \N__47996\
        );

    \I__10911\ : LocalMux
    port map (
            O => \N__48112\,
            I => \N__47989\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__48109\,
            I => \N__47989\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__48106\,
            I => \N__47989\
        );

    \I__10908\ : Span4Mux_v
    port map (
            O => \N__48101\,
            I => \N__47976\
        );

    \I__10907\ : LocalMux
    port map (
            O => \N__48098\,
            I => \N__47976\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__48095\,
            I => \N__47976\
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__48092\,
            I => \N__47976\
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__48089\,
            I => \N__47976\
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__48086\,
            I => \N__47976\
        );

    \I__10902\ : Span4Mux_v
    port map (
            O => \N__48075\,
            I => \N__47972\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__48072\,
            I => \N__47963\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__48069\,
            I => \N__47963\
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__48066\,
            I => \N__47963\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__48063\,
            I => \N__47963\
        );

    \I__10897\ : InMux
    port map (
            O => \N__48062\,
            I => \N__47960\
        );

    \I__10896\ : Span4Mux_v
    port map (
            O => \N__48053\,
            I => \N__47949\
        );

    \I__10895\ : Span4Mux_h
    port map (
            O => \N__48046\,
            I => \N__47949\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__48043\,
            I => \N__47949\
        );

    \I__10893\ : LocalMux
    port map (
            O => \N__48040\,
            I => \N__47949\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__48037\,
            I => \N__47949\
        );

    \I__10891\ : Sp12to4
    port map (
            O => \N__48034\,
            I => \N__47943\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__48031\,
            I => \N__47943\
        );

    \I__10889\ : Span4Mux_v
    port map (
            O => \N__48026\,
            I => \N__47938\
        );

    \I__10888\ : LocalMux
    port map (
            O => \N__48023\,
            I => \N__47938\
        );

    \I__10887\ : Span4Mux_v
    port map (
            O => \N__48014\,
            I => \N__47931\
        );

    \I__10886\ : Span4Mux_h
    port map (
            O => \N__48007\,
            I => \N__47931\
        );

    \I__10885\ : LocalMux
    port map (
            O => \N__48004\,
            I => \N__47931\
        );

    \I__10884\ : Span12Mux_h
    port map (
            O => \N__48001\,
            I => \N__47926\
        );

    \I__10883\ : Span12Mux_s11_v
    port map (
            O => \N__47996\,
            I => \N__47926\
        );

    \I__10882\ : Span4Mux_v
    port map (
            O => \N__47989\,
            I => \N__47923\
        );

    \I__10881\ : Span4Mux_v
    port map (
            O => \N__47976\,
            I => \N__47920\
        );

    \I__10880\ : InMux
    port map (
            O => \N__47975\,
            I => \N__47917\
        );

    \I__10879\ : Span4Mux_h
    port map (
            O => \N__47972\,
            I => \N__47908\
        );

    \I__10878\ : Span4Mux_v
    port map (
            O => \N__47963\,
            I => \N__47908\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__47960\,
            I => \N__47908\
        );

    \I__10876\ : Span4Mux_v
    port map (
            O => \N__47949\,
            I => \N__47908\
        );

    \I__10875\ : CascadeMux
    port map (
            O => \N__47948\,
            I => \N__47905\
        );

    \I__10874\ : Span12Mux_h
    port map (
            O => \N__47943\,
            I => \N__47902\
        );

    \I__10873\ : Span4Mux_v
    port map (
            O => \N__47938\,
            I => \N__47899\
        );

    \I__10872\ : Span4Mux_v
    port map (
            O => \N__47931\,
            I => \N__47896\
        );

    \I__10871\ : Span12Mux_v
    port map (
            O => \N__47926\,
            I => \N__47887\
        );

    \I__10870\ : Sp12to4
    port map (
            O => \N__47923\,
            I => \N__47887\
        );

    \I__10869\ : Sp12to4
    port map (
            O => \N__47920\,
            I => \N__47887\
        );

    \I__10868\ : LocalMux
    port map (
            O => \N__47917\,
            I => \N__47887\
        );

    \I__10867\ : Span4Mux_h
    port map (
            O => \N__47908\,
            I => \N__47884\
        );

    \I__10866\ : InMux
    port map (
            O => \N__47905\,
            I => \N__47881\
        );

    \I__10865\ : Odrv12
    port map (
            O => \N__47902\,
            I => spi_data_mosi_6
        );

    \I__10864\ : Odrv4
    port map (
            O => \N__47899\,
            I => spi_data_mosi_6
        );

    \I__10863\ : Odrv4
    port map (
            O => \N__47896\,
            I => spi_data_mosi_6
        );

    \I__10862\ : Odrv12
    port map (
            O => \N__47887\,
            I => spi_data_mosi_6
        );

    \I__10861\ : Odrv4
    port map (
            O => \N__47884\,
            I => spi_data_mosi_6
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__47881\,
            I => spi_data_mosi_6
        );

    \I__10859\ : InMux
    port map (
            O => \N__47868\,
            I => \N__47865\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__47865\,
            I => \N__47862\
        );

    \I__10857\ : Span4Mux_h
    port map (
            O => \N__47862\,
            I => \N__47859\
        );

    \I__10856\ : Span4Mux_h
    port map (
            O => \N__47859\,
            I => \N__47856\
        );

    \I__10855\ : Odrv4
    port map (
            O => \N__47856\,
            I => \sDAC_mem_12Z0Z_6\
        );

    \I__10854\ : ClkMux
    port map (
            O => \N__47853\,
            I => \N__47397\
        );

    \I__10853\ : ClkMux
    port map (
            O => \N__47852\,
            I => \N__47397\
        );

    \I__10852\ : ClkMux
    port map (
            O => \N__47851\,
            I => \N__47397\
        );

    \I__10851\ : ClkMux
    port map (
            O => \N__47850\,
            I => \N__47397\
        );

    \I__10850\ : ClkMux
    port map (
            O => \N__47849\,
            I => \N__47397\
        );

    \I__10849\ : ClkMux
    port map (
            O => \N__47848\,
            I => \N__47397\
        );

    \I__10848\ : ClkMux
    port map (
            O => \N__47847\,
            I => \N__47397\
        );

    \I__10847\ : ClkMux
    port map (
            O => \N__47846\,
            I => \N__47397\
        );

    \I__10846\ : ClkMux
    port map (
            O => \N__47845\,
            I => \N__47397\
        );

    \I__10845\ : ClkMux
    port map (
            O => \N__47844\,
            I => \N__47397\
        );

    \I__10844\ : ClkMux
    port map (
            O => \N__47843\,
            I => \N__47397\
        );

    \I__10843\ : ClkMux
    port map (
            O => \N__47842\,
            I => \N__47397\
        );

    \I__10842\ : ClkMux
    port map (
            O => \N__47841\,
            I => \N__47397\
        );

    \I__10841\ : ClkMux
    port map (
            O => \N__47840\,
            I => \N__47397\
        );

    \I__10840\ : ClkMux
    port map (
            O => \N__47839\,
            I => \N__47397\
        );

    \I__10839\ : ClkMux
    port map (
            O => \N__47838\,
            I => \N__47397\
        );

    \I__10838\ : ClkMux
    port map (
            O => \N__47837\,
            I => \N__47397\
        );

    \I__10837\ : ClkMux
    port map (
            O => \N__47836\,
            I => \N__47397\
        );

    \I__10836\ : ClkMux
    port map (
            O => \N__47835\,
            I => \N__47397\
        );

    \I__10835\ : ClkMux
    port map (
            O => \N__47834\,
            I => \N__47397\
        );

    \I__10834\ : ClkMux
    port map (
            O => \N__47833\,
            I => \N__47397\
        );

    \I__10833\ : ClkMux
    port map (
            O => \N__47832\,
            I => \N__47397\
        );

    \I__10832\ : ClkMux
    port map (
            O => \N__47831\,
            I => \N__47397\
        );

    \I__10831\ : ClkMux
    port map (
            O => \N__47830\,
            I => \N__47397\
        );

    \I__10830\ : ClkMux
    port map (
            O => \N__47829\,
            I => \N__47397\
        );

    \I__10829\ : ClkMux
    port map (
            O => \N__47828\,
            I => \N__47397\
        );

    \I__10828\ : ClkMux
    port map (
            O => \N__47827\,
            I => \N__47397\
        );

    \I__10827\ : ClkMux
    port map (
            O => \N__47826\,
            I => \N__47397\
        );

    \I__10826\ : ClkMux
    port map (
            O => \N__47825\,
            I => \N__47397\
        );

    \I__10825\ : ClkMux
    port map (
            O => \N__47824\,
            I => \N__47397\
        );

    \I__10824\ : ClkMux
    port map (
            O => \N__47823\,
            I => \N__47397\
        );

    \I__10823\ : ClkMux
    port map (
            O => \N__47822\,
            I => \N__47397\
        );

    \I__10822\ : ClkMux
    port map (
            O => \N__47821\,
            I => \N__47397\
        );

    \I__10821\ : ClkMux
    port map (
            O => \N__47820\,
            I => \N__47397\
        );

    \I__10820\ : ClkMux
    port map (
            O => \N__47819\,
            I => \N__47397\
        );

    \I__10819\ : ClkMux
    port map (
            O => \N__47818\,
            I => \N__47397\
        );

    \I__10818\ : ClkMux
    port map (
            O => \N__47817\,
            I => \N__47397\
        );

    \I__10817\ : ClkMux
    port map (
            O => \N__47816\,
            I => \N__47397\
        );

    \I__10816\ : ClkMux
    port map (
            O => \N__47815\,
            I => \N__47397\
        );

    \I__10815\ : ClkMux
    port map (
            O => \N__47814\,
            I => \N__47397\
        );

    \I__10814\ : ClkMux
    port map (
            O => \N__47813\,
            I => \N__47397\
        );

    \I__10813\ : ClkMux
    port map (
            O => \N__47812\,
            I => \N__47397\
        );

    \I__10812\ : ClkMux
    port map (
            O => \N__47811\,
            I => \N__47397\
        );

    \I__10811\ : ClkMux
    port map (
            O => \N__47810\,
            I => \N__47397\
        );

    \I__10810\ : ClkMux
    port map (
            O => \N__47809\,
            I => \N__47397\
        );

    \I__10809\ : ClkMux
    port map (
            O => \N__47808\,
            I => \N__47397\
        );

    \I__10808\ : ClkMux
    port map (
            O => \N__47807\,
            I => \N__47397\
        );

    \I__10807\ : ClkMux
    port map (
            O => \N__47806\,
            I => \N__47397\
        );

    \I__10806\ : ClkMux
    port map (
            O => \N__47805\,
            I => \N__47397\
        );

    \I__10805\ : ClkMux
    port map (
            O => \N__47804\,
            I => \N__47397\
        );

    \I__10804\ : ClkMux
    port map (
            O => \N__47803\,
            I => \N__47397\
        );

    \I__10803\ : ClkMux
    port map (
            O => \N__47802\,
            I => \N__47397\
        );

    \I__10802\ : ClkMux
    port map (
            O => \N__47801\,
            I => \N__47397\
        );

    \I__10801\ : ClkMux
    port map (
            O => \N__47800\,
            I => \N__47397\
        );

    \I__10800\ : ClkMux
    port map (
            O => \N__47799\,
            I => \N__47397\
        );

    \I__10799\ : ClkMux
    port map (
            O => \N__47798\,
            I => \N__47397\
        );

    \I__10798\ : ClkMux
    port map (
            O => \N__47797\,
            I => \N__47397\
        );

    \I__10797\ : ClkMux
    port map (
            O => \N__47796\,
            I => \N__47397\
        );

    \I__10796\ : ClkMux
    port map (
            O => \N__47795\,
            I => \N__47397\
        );

    \I__10795\ : ClkMux
    port map (
            O => \N__47794\,
            I => \N__47397\
        );

    \I__10794\ : ClkMux
    port map (
            O => \N__47793\,
            I => \N__47397\
        );

    \I__10793\ : ClkMux
    port map (
            O => \N__47792\,
            I => \N__47397\
        );

    \I__10792\ : ClkMux
    port map (
            O => \N__47791\,
            I => \N__47397\
        );

    \I__10791\ : ClkMux
    port map (
            O => \N__47790\,
            I => \N__47397\
        );

    \I__10790\ : ClkMux
    port map (
            O => \N__47789\,
            I => \N__47397\
        );

    \I__10789\ : ClkMux
    port map (
            O => \N__47788\,
            I => \N__47397\
        );

    \I__10788\ : ClkMux
    port map (
            O => \N__47787\,
            I => \N__47397\
        );

    \I__10787\ : ClkMux
    port map (
            O => \N__47786\,
            I => \N__47397\
        );

    \I__10786\ : ClkMux
    port map (
            O => \N__47785\,
            I => \N__47397\
        );

    \I__10785\ : ClkMux
    port map (
            O => \N__47784\,
            I => \N__47397\
        );

    \I__10784\ : ClkMux
    port map (
            O => \N__47783\,
            I => \N__47397\
        );

    \I__10783\ : ClkMux
    port map (
            O => \N__47782\,
            I => \N__47397\
        );

    \I__10782\ : ClkMux
    port map (
            O => \N__47781\,
            I => \N__47397\
        );

    \I__10781\ : ClkMux
    port map (
            O => \N__47780\,
            I => \N__47397\
        );

    \I__10780\ : ClkMux
    port map (
            O => \N__47779\,
            I => \N__47397\
        );

    \I__10779\ : ClkMux
    port map (
            O => \N__47778\,
            I => \N__47397\
        );

    \I__10778\ : ClkMux
    port map (
            O => \N__47777\,
            I => \N__47397\
        );

    \I__10777\ : ClkMux
    port map (
            O => \N__47776\,
            I => \N__47397\
        );

    \I__10776\ : ClkMux
    port map (
            O => \N__47775\,
            I => \N__47397\
        );

    \I__10775\ : ClkMux
    port map (
            O => \N__47774\,
            I => \N__47397\
        );

    \I__10774\ : ClkMux
    port map (
            O => \N__47773\,
            I => \N__47397\
        );

    \I__10773\ : ClkMux
    port map (
            O => \N__47772\,
            I => \N__47397\
        );

    \I__10772\ : ClkMux
    port map (
            O => \N__47771\,
            I => \N__47397\
        );

    \I__10771\ : ClkMux
    port map (
            O => \N__47770\,
            I => \N__47397\
        );

    \I__10770\ : ClkMux
    port map (
            O => \N__47769\,
            I => \N__47397\
        );

    \I__10769\ : ClkMux
    port map (
            O => \N__47768\,
            I => \N__47397\
        );

    \I__10768\ : ClkMux
    port map (
            O => \N__47767\,
            I => \N__47397\
        );

    \I__10767\ : ClkMux
    port map (
            O => \N__47766\,
            I => \N__47397\
        );

    \I__10766\ : ClkMux
    port map (
            O => \N__47765\,
            I => \N__47397\
        );

    \I__10765\ : ClkMux
    port map (
            O => \N__47764\,
            I => \N__47397\
        );

    \I__10764\ : ClkMux
    port map (
            O => \N__47763\,
            I => \N__47397\
        );

    \I__10763\ : ClkMux
    port map (
            O => \N__47762\,
            I => \N__47397\
        );

    \I__10762\ : ClkMux
    port map (
            O => \N__47761\,
            I => \N__47397\
        );

    \I__10761\ : ClkMux
    port map (
            O => \N__47760\,
            I => \N__47397\
        );

    \I__10760\ : ClkMux
    port map (
            O => \N__47759\,
            I => \N__47397\
        );

    \I__10759\ : ClkMux
    port map (
            O => \N__47758\,
            I => \N__47397\
        );

    \I__10758\ : ClkMux
    port map (
            O => \N__47757\,
            I => \N__47397\
        );

    \I__10757\ : ClkMux
    port map (
            O => \N__47756\,
            I => \N__47397\
        );

    \I__10756\ : ClkMux
    port map (
            O => \N__47755\,
            I => \N__47397\
        );

    \I__10755\ : ClkMux
    port map (
            O => \N__47754\,
            I => \N__47397\
        );

    \I__10754\ : ClkMux
    port map (
            O => \N__47753\,
            I => \N__47397\
        );

    \I__10753\ : ClkMux
    port map (
            O => \N__47752\,
            I => \N__47397\
        );

    \I__10752\ : ClkMux
    port map (
            O => \N__47751\,
            I => \N__47397\
        );

    \I__10751\ : ClkMux
    port map (
            O => \N__47750\,
            I => \N__47397\
        );

    \I__10750\ : ClkMux
    port map (
            O => \N__47749\,
            I => \N__47397\
        );

    \I__10749\ : ClkMux
    port map (
            O => \N__47748\,
            I => \N__47397\
        );

    \I__10748\ : ClkMux
    port map (
            O => \N__47747\,
            I => \N__47397\
        );

    \I__10747\ : ClkMux
    port map (
            O => \N__47746\,
            I => \N__47397\
        );

    \I__10746\ : ClkMux
    port map (
            O => \N__47745\,
            I => \N__47397\
        );

    \I__10745\ : ClkMux
    port map (
            O => \N__47744\,
            I => \N__47397\
        );

    \I__10744\ : ClkMux
    port map (
            O => \N__47743\,
            I => \N__47397\
        );

    \I__10743\ : ClkMux
    port map (
            O => \N__47742\,
            I => \N__47397\
        );

    \I__10742\ : ClkMux
    port map (
            O => \N__47741\,
            I => \N__47397\
        );

    \I__10741\ : ClkMux
    port map (
            O => \N__47740\,
            I => \N__47397\
        );

    \I__10740\ : ClkMux
    port map (
            O => \N__47739\,
            I => \N__47397\
        );

    \I__10739\ : ClkMux
    port map (
            O => \N__47738\,
            I => \N__47397\
        );

    \I__10738\ : ClkMux
    port map (
            O => \N__47737\,
            I => \N__47397\
        );

    \I__10737\ : ClkMux
    port map (
            O => \N__47736\,
            I => \N__47397\
        );

    \I__10736\ : ClkMux
    port map (
            O => \N__47735\,
            I => \N__47397\
        );

    \I__10735\ : ClkMux
    port map (
            O => \N__47734\,
            I => \N__47397\
        );

    \I__10734\ : ClkMux
    port map (
            O => \N__47733\,
            I => \N__47397\
        );

    \I__10733\ : ClkMux
    port map (
            O => \N__47732\,
            I => \N__47397\
        );

    \I__10732\ : ClkMux
    port map (
            O => \N__47731\,
            I => \N__47397\
        );

    \I__10731\ : ClkMux
    port map (
            O => \N__47730\,
            I => \N__47397\
        );

    \I__10730\ : ClkMux
    port map (
            O => \N__47729\,
            I => \N__47397\
        );

    \I__10729\ : ClkMux
    port map (
            O => \N__47728\,
            I => \N__47397\
        );

    \I__10728\ : ClkMux
    port map (
            O => \N__47727\,
            I => \N__47397\
        );

    \I__10727\ : ClkMux
    port map (
            O => \N__47726\,
            I => \N__47397\
        );

    \I__10726\ : ClkMux
    port map (
            O => \N__47725\,
            I => \N__47397\
        );

    \I__10725\ : ClkMux
    port map (
            O => \N__47724\,
            I => \N__47397\
        );

    \I__10724\ : ClkMux
    port map (
            O => \N__47723\,
            I => \N__47397\
        );

    \I__10723\ : ClkMux
    port map (
            O => \N__47722\,
            I => \N__47397\
        );

    \I__10722\ : ClkMux
    port map (
            O => \N__47721\,
            I => \N__47397\
        );

    \I__10721\ : ClkMux
    port map (
            O => \N__47720\,
            I => \N__47397\
        );

    \I__10720\ : ClkMux
    port map (
            O => \N__47719\,
            I => \N__47397\
        );

    \I__10719\ : ClkMux
    port map (
            O => \N__47718\,
            I => \N__47397\
        );

    \I__10718\ : ClkMux
    port map (
            O => \N__47717\,
            I => \N__47397\
        );

    \I__10717\ : ClkMux
    port map (
            O => \N__47716\,
            I => \N__47397\
        );

    \I__10716\ : ClkMux
    port map (
            O => \N__47715\,
            I => \N__47397\
        );

    \I__10715\ : ClkMux
    port map (
            O => \N__47714\,
            I => \N__47397\
        );

    \I__10714\ : ClkMux
    port map (
            O => \N__47713\,
            I => \N__47397\
        );

    \I__10713\ : ClkMux
    port map (
            O => \N__47712\,
            I => \N__47397\
        );

    \I__10712\ : ClkMux
    port map (
            O => \N__47711\,
            I => \N__47397\
        );

    \I__10711\ : ClkMux
    port map (
            O => \N__47710\,
            I => \N__47397\
        );

    \I__10710\ : ClkMux
    port map (
            O => \N__47709\,
            I => \N__47397\
        );

    \I__10709\ : ClkMux
    port map (
            O => \N__47708\,
            I => \N__47397\
        );

    \I__10708\ : ClkMux
    port map (
            O => \N__47707\,
            I => \N__47397\
        );

    \I__10707\ : ClkMux
    port map (
            O => \N__47706\,
            I => \N__47397\
        );

    \I__10706\ : ClkMux
    port map (
            O => \N__47705\,
            I => \N__47397\
        );

    \I__10705\ : ClkMux
    port map (
            O => \N__47704\,
            I => \N__47397\
        );

    \I__10704\ : ClkMux
    port map (
            O => \N__47703\,
            I => \N__47397\
        );

    \I__10703\ : ClkMux
    port map (
            O => \N__47702\,
            I => \N__47397\
        );

    \I__10702\ : GlobalMux
    port map (
            O => \N__47397\,
            I => \N__47394\
        );

    \I__10701\ : gio2CtrlBuf
    port map (
            O => \N__47394\,
            I => pll_clk128_g
        );

    \I__10700\ : CEMux
    port map (
            O => \N__47391\,
            I => \N__47388\
        );

    \I__10699\ : LocalMux
    port map (
            O => \N__47388\,
            I => \N__47385\
        );

    \I__10698\ : Span4Mux_v
    port map (
            O => \N__47385\,
            I => \N__47381\
        );

    \I__10697\ : CEMux
    port map (
            O => \N__47384\,
            I => \N__47378\
        );

    \I__10696\ : Span4Mux_h
    port map (
            O => \N__47381\,
            I => \N__47372\
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__47378\,
            I => \N__47369\
        );

    \I__10694\ : CEMux
    port map (
            O => \N__47377\,
            I => \N__47366\
        );

    \I__10693\ : CEMux
    port map (
            O => \N__47376\,
            I => \N__47363\
        );

    \I__10692\ : CEMux
    port map (
            O => \N__47375\,
            I => \N__47360\
        );

    \I__10691\ : Span4Mux_h
    port map (
            O => \N__47372\,
            I => \N__47353\
        );

    \I__10690\ : Span4Mux_h
    port map (
            O => \N__47369\,
            I => \N__47353\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__47366\,
            I => \N__47353\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__47363\,
            I => \N__47350\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__47360\,
            I => \N__47347\
        );

    \I__10686\ : Odrv4
    port map (
            O => \N__47353\,
            I => \sDAC_mem_12_1_sqmuxa\
        );

    \I__10685\ : Odrv4
    port map (
            O => \N__47350\,
            I => \sDAC_mem_12_1_sqmuxa\
        );

    \I__10684\ : Odrv4
    port map (
            O => \N__47347\,
            I => \sDAC_mem_12_1_sqmuxa\
        );

    \I__10683\ : InMux
    port map (
            O => \N__47340\,
            I => \N__47337\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__47337\,
            I => \N__47334\
        );

    \I__10681\ : Span4Mux_h
    port map (
            O => \N__47334\,
            I => \N__47331\
        );

    \I__10680\ : Span4Mux_h
    port map (
            O => \N__47331\,
            I => \N__47328\
        );

    \I__10679\ : Odrv4
    port map (
            O => \N__47328\,
            I => \sDAC_mem_9Z0Z_7\
        );

    \I__10678\ : CEMux
    port map (
            O => \N__47325\,
            I => \N__47322\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__47322\,
            I => \N__47319\
        );

    \I__10676\ : Span4Mux_v
    port map (
            O => \N__47319\,
            I => \N__47316\
        );

    \I__10675\ : Odrv4
    port map (
            O => \N__47316\,
            I => \sDAC_mem_9_1_sqmuxa\
        );

    \I__10674\ : CascadeMux
    port map (
            O => \N__47313\,
            I => \N_14_3_cascade_\
        );

    \I__10673\ : CascadeMux
    port map (
            O => \N__47310\,
            I => \N_8_cascade_\
        );

    \I__10672\ : InMux
    port map (
            O => \N__47307\,
            I => \N__47301\
        );

    \I__10671\ : InMux
    port map (
            O => \N__47306\,
            I => \N__47301\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__47301\,
            I => \N__47297\
        );

    \I__10669\ : InMux
    port map (
            O => \N__47300\,
            I => \N__47294\
        );

    \I__10668\ : Span12Mux_h
    port map (
            O => \N__47297\,
            I => \N__47291\
        );

    \I__10667\ : LocalMux
    port map (
            O => \N__47294\,
            I => \sDAC_spi_startZ0\
        );

    \I__10666\ : Odrv12
    port map (
            O => \N__47291\,
            I => \sDAC_spi_startZ0\
        );

    \I__10665\ : InMux
    port map (
            O => \N__47286\,
            I => \N__47283\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__47283\,
            I => un1_scounterdac8_i_a2_1_2
        );

    \I__10663\ : InMux
    port map (
            O => \N__47280\,
            I => \N__47277\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__47277\,
            I => un1_scounterdac8_i_a2_0
        );

    \I__10661\ : InMux
    port map (
            O => \N__47274\,
            I => \N__47271\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__47271\,
            I => \N__47268\
        );

    \I__10659\ : Span4Mux_h
    port map (
            O => \N__47268\,
            I => \N__47265\
        );

    \I__10658\ : Odrv4
    port map (
            O => \N__47265\,
            I => \sDAC_data_RNO_18Z0Z_10\
        );

    \I__10657\ : InMux
    port map (
            O => \N__47262\,
            I => \N__47259\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__47259\,
            I => \N__47256\
        );

    \I__10655\ : Span4Mux_h
    port map (
            O => \N__47256\,
            I => \N__47253\
        );

    \I__10654\ : Odrv4
    port map (
            O => \N__47253\,
            I => \sEEDACZ0Z_5\
        );

    \I__10653\ : InMux
    port map (
            O => \N__47250\,
            I => \N__47247\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__47247\,
            I => \N__47244\
        );

    \I__10651\ : Span4Mux_h
    port map (
            O => \N__47244\,
            I => \N__47241\
        );

    \I__10650\ : Odrv4
    port map (
            O => \N__47241\,
            I => \sEEDACZ0Z_6\
        );

    \I__10649\ : CEMux
    port map (
            O => \N__47238\,
            I => \N__47235\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__47235\,
            I => \N__47231\
        );

    \I__10647\ : CEMux
    port map (
            O => \N__47234\,
            I => \N__47228\
        );

    \I__10646\ : Span4Mux_h
    port map (
            O => \N__47231\,
            I => \N__47225\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__47228\,
            I => \N__47222\
        );

    \I__10644\ : Odrv4
    port map (
            O => \N__47225\,
            I => \sEEDAC_1_sqmuxa\
        );

    \I__10643\ : Odrv4
    port map (
            O => \N__47222\,
            I => \sEEDAC_1_sqmuxa\
        );

    \I__10642\ : InMux
    port map (
            O => \N__47217\,
            I => \N__47214\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__47214\,
            I => \N__47211\
        );

    \I__10640\ : Span4Mux_h
    port map (
            O => \N__47211\,
            I => \N__47208\
        );

    \I__10639\ : Odrv4
    port map (
            O => \N__47208\,
            I => \sDAC_mem_9Z0Z_0\
        );

    \I__10638\ : InMux
    port map (
            O => \N__47205\,
            I => \N__47202\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__47202\,
            I => \N__47199\
        );

    \I__10636\ : Span4Mux_v
    port map (
            O => \N__47199\,
            I => \N__47196\
        );

    \I__10635\ : Odrv4
    port map (
            O => \N__47196\,
            I => \sDAC_mem_9Z0Z_1\
        );

    \I__10634\ : InMux
    port map (
            O => \N__47193\,
            I => \N__47190\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__47190\,
            I => \N__47187\
        );

    \I__10632\ : Span4Mux_h
    port map (
            O => \N__47187\,
            I => \N__47184\
        );

    \I__10631\ : Span4Mux_h
    port map (
            O => \N__47184\,
            I => \N__47181\
        );

    \I__10630\ : Odrv4
    port map (
            O => \N__47181\,
            I => \sDAC_mem_9Z0Z_2\
        );

    \I__10629\ : InMux
    port map (
            O => \N__47178\,
            I => \N__47175\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__47175\,
            I => \N__47172\
        );

    \I__10627\ : Span4Mux_h
    port map (
            O => \N__47172\,
            I => \N__47169\
        );

    \I__10626\ : Odrv4
    port map (
            O => \N__47169\,
            I => \sDAC_mem_9Z0Z_3\
        );

    \I__10625\ : InMux
    port map (
            O => \N__47166\,
            I => \N__47163\
        );

    \I__10624\ : LocalMux
    port map (
            O => \N__47163\,
            I => \N__47160\
        );

    \I__10623\ : Span4Mux_h
    port map (
            O => \N__47160\,
            I => \N__47157\
        );

    \I__10622\ : Span4Mux_h
    port map (
            O => \N__47157\,
            I => \N__47154\
        );

    \I__10621\ : Odrv4
    port map (
            O => \N__47154\,
            I => \sDAC_mem_9Z0Z_4\
        );

    \I__10620\ : InMux
    port map (
            O => \N__47151\,
            I => \N__47144\
        );

    \I__10619\ : InMux
    port map (
            O => \N__47150\,
            I => \N__47141\
        );

    \I__10618\ : InMux
    port map (
            O => \N__47149\,
            I => \N__47127\
        );

    \I__10617\ : InMux
    port map (
            O => \N__47148\,
            I => \N__47123\
        );

    \I__10616\ : InMux
    port map (
            O => \N__47147\,
            I => \N__47120\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__47144\,
            I => \N__47112\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__47141\,
            I => \N__47112\
        );

    \I__10613\ : InMux
    port map (
            O => \N__47140\,
            I => \N__47109\
        );

    \I__10612\ : InMux
    port map (
            O => \N__47139\,
            I => \N__47106\
        );

    \I__10611\ : InMux
    port map (
            O => \N__47138\,
            I => \N__47103\
        );

    \I__10610\ : InMux
    port map (
            O => \N__47137\,
            I => \N__47100\
        );

    \I__10609\ : InMux
    port map (
            O => \N__47136\,
            I => \N__47096\
        );

    \I__10608\ : InMux
    port map (
            O => \N__47135\,
            I => \N__47093\
        );

    \I__10607\ : InMux
    port map (
            O => \N__47134\,
            I => \N__47090\
        );

    \I__10606\ : InMux
    port map (
            O => \N__47133\,
            I => \N__47085\
        );

    \I__10605\ : InMux
    port map (
            O => \N__47132\,
            I => \N__47082\
        );

    \I__10604\ : InMux
    port map (
            O => \N__47131\,
            I => \N__47078\
        );

    \I__10603\ : InMux
    port map (
            O => \N__47130\,
            I => \N__47075\
        );

    \I__10602\ : LocalMux
    port map (
            O => \N__47127\,
            I => \N__47068\
        );

    \I__10601\ : InMux
    port map (
            O => \N__47126\,
            I => \N__47065\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__47123\,
            I => \N__47057\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__47120\,
            I => \N__47057\
        );

    \I__10598\ : InMux
    port map (
            O => \N__47119\,
            I => \N__47054\
        );

    \I__10597\ : InMux
    port map (
            O => \N__47118\,
            I => \N__47050\
        );

    \I__10596\ : InMux
    port map (
            O => \N__47117\,
            I => \N__47047\
        );

    \I__10595\ : Span4Mux_v
    port map (
            O => \N__47112\,
            I => \N__47034\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__47109\,
            I => \N__47034\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__47106\,
            I => \N__47034\
        );

    \I__10592\ : LocalMux
    port map (
            O => \N__47103\,
            I => \N__47034\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__47100\,
            I => \N__47034\
        );

    \I__10590\ : InMux
    port map (
            O => \N__47099\,
            I => \N__47031\
        );

    \I__10589\ : LocalMux
    port map (
            O => \N__47096\,
            I => \N__47024\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__47093\,
            I => \N__47024\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__47090\,
            I => \N__47024\
        );

    \I__10586\ : InMux
    port map (
            O => \N__47089\,
            I => \N__47021\
        );

    \I__10585\ : InMux
    port map (
            O => \N__47088\,
            I => \N__47018\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__47085\,
            I => \N__47013\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__47082\,
            I => \N__47010\
        );

    \I__10582\ : InMux
    port map (
            O => \N__47081\,
            I => \N__47007\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__47078\,
            I => \N__47004\
        );

    \I__10580\ : LocalMux
    port map (
            O => \N__47075\,
            I => \N__47001\
        );

    \I__10579\ : InMux
    port map (
            O => \N__47074\,
            I => \N__46998\
        );

    \I__10578\ : InMux
    port map (
            O => \N__47073\,
            I => \N__46995\
        );

    \I__10577\ : InMux
    port map (
            O => \N__47072\,
            I => \N__46990\
        );

    \I__10576\ : InMux
    port map (
            O => \N__47071\,
            I => \N__46987\
        );

    \I__10575\ : Span4Mux_h
    port map (
            O => \N__47068\,
            I => \N__46980\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__47065\,
            I => \N__46977\
        );

    \I__10573\ : InMux
    port map (
            O => \N__47064\,
            I => \N__46974\
        );

    \I__10572\ : InMux
    port map (
            O => \N__47063\,
            I => \N__46971\
        );

    \I__10571\ : InMux
    port map (
            O => \N__47062\,
            I => \N__46967\
        );

    \I__10570\ : Span4Mux_h
    port map (
            O => \N__47057\,
            I => \N__46962\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__47054\,
            I => \N__46962\
        );

    \I__10568\ : InMux
    port map (
            O => \N__47053\,
            I => \N__46959\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__47050\,
            I => \N__46953\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__47047\,
            I => \N__46950\
        );

    \I__10565\ : InMux
    port map (
            O => \N__47046\,
            I => \N__46947\
        );

    \I__10564\ : InMux
    port map (
            O => \N__47045\,
            I => \N__46944\
        );

    \I__10563\ : Span4Mux_v
    port map (
            O => \N__47034\,
            I => \N__46939\
        );

    \I__10562\ : LocalMux
    port map (
            O => \N__47031\,
            I => \N__46939\
        );

    \I__10561\ : Span4Mux_v
    port map (
            O => \N__47024\,
            I => \N__46934\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__47021\,
            I => \N__46934\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__47018\,
            I => \N__46931\
        );

    \I__10558\ : InMux
    port map (
            O => \N__47017\,
            I => \N__46928\
        );

    \I__10557\ : InMux
    port map (
            O => \N__47016\,
            I => \N__46925\
        );

    \I__10556\ : Span4Mux_v
    port map (
            O => \N__47013\,
            I => \N__46918\
        );

    \I__10555\ : Span4Mux_h
    port map (
            O => \N__47010\,
            I => \N__46918\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__47007\,
            I => \N__46918\
        );

    \I__10553\ : Span4Mux_h
    port map (
            O => \N__47004\,
            I => \N__46913\
        );

    \I__10552\ : Span4Mux_h
    port map (
            O => \N__47001\,
            I => \N__46913\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__46998\,
            I => \N__46908\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__46995\,
            I => \N__46908\
        );

    \I__10549\ : InMux
    port map (
            O => \N__46994\,
            I => \N__46905\
        );

    \I__10548\ : InMux
    port map (
            O => \N__46993\,
            I => \N__46902\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__46990\,
            I => \N__46899\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__46987\,
            I => \N__46894\
        );

    \I__10545\ : InMux
    port map (
            O => \N__46986\,
            I => \N__46891\
        );

    \I__10544\ : InMux
    port map (
            O => \N__46985\,
            I => \N__46888\
        );

    \I__10543\ : InMux
    port map (
            O => \N__46984\,
            I => \N__46885\
        );

    \I__10542\ : InMux
    port map (
            O => \N__46983\,
            I => \N__46882\
        );

    \I__10541\ : Span4Mux_v
    port map (
            O => \N__46980\,
            I => \N__46871\
        );

    \I__10540\ : Span4Mux_h
    port map (
            O => \N__46977\,
            I => \N__46871\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__46974\,
            I => \N__46868\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__46971\,
            I => \N__46865\
        );

    \I__10537\ : InMux
    port map (
            O => \N__46970\,
            I => \N__46862\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__46967\,
            I => \N__46858\
        );

    \I__10535\ : Span4Mux_h
    port map (
            O => \N__46962\,
            I => \N__46853\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__46959\,
            I => \N__46853\
        );

    \I__10533\ : InMux
    port map (
            O => \N__46958\,
            I => \N__46850\
        );

    \I__10532\ : InMux
    port map (
            O => \N__46957\,
            I => \N__46845\
        );

    \I__10531\ : InMux
    port map (
            O => \N__46956\,
            I => \N__46845\
        );

    \I__10530\ : Span4Mux_h
    port map (
            O => \N__46953\,
            I => \N__46842\
        );

    \I__10529\ : Span4Mux_h
    port map (
            O => \N__46950\,
            I => \N__46835\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__46947\,
            I => \N__46835\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__46944\,
            I => \N__46835\
        );

    \I__10526\ : Span4Mux_h
    port map (
            O => \N__46939\,
            I => \N__46832\
        );

    \I__10525\ : Span4Mux_v
    port map (
            O => \N__46934\,
            I => \N__46823\
        );

    \I__10524\ : Span4Mux_h
    port map (
            O => \N__46931\,
            I => \N__46823\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__46928\,
            I => \N__46823\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__46925\,
            I => \N__46823\
        );

    \I__10521\ : Span4Mux_v
    port map (
            O => \N__46918\,
            I => \N__46820\
        );

    \I__10520\ : Span4Mux_v
    port map (
            O => \N__46913\,
            I => \N__46811\
        );

    \I__10519\ : Span4Mux_h
    port map (
            O => \N__46908\,
            I => \N__46811\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__46905\,
            I => \N__46811\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__46902\,
            I => \N__46811\
        );

    \I__10516\ : Span4Mux_h
    port map (
            O => \N__46899\,
            I => \N__46808\
        );

    \I__10515\ : InMux
    port map (
            O => \N__46898\,
            I => \N__46805\
        );

    \I__10514\ : InMux
    port map (
            O => \N__46897\,
            I => \N__46802\
        );

    \I__10513\ : Span4Mux_h
    port map (
            O => \N__46894\,
            I => \N__46795\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__46891\,
            I => \N__46795\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__46888\,
            I => \N__46795\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__46885\,
            I => \N__46788\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__46882\,
            I => \N__46788\
        );

    \I__10508\ : InMux
    port map (
            O => \N__46881\,
            I => \N__46785\
        );

    \I__10507\ : InMux
    port map (
            O => \N__46880\,
            I => \N__46782\
        );

    \I__10506\ : InMux
    port map (
            O => \N__46879\,
            I => \N__46779\
        );

    \I__10505\ : InMux
    port map (
            O => \N__46878\,
            I => \N__46776\
        );

    \I__10504\ : InMux
    port map (
            O => \N__46877\,
            I => \N__46773\
        );

    \I__10503\ : InMux
    port map (
            O => \N__46876\,
            I => \N__46770\
        );

    \I__10502\ : Span4Mux_v
    port map (
            O => \N__46871\,
            I => \N__46766\
        );

    \I__10501\ : Span4Mux_v
    port map (
            O => \N__46868\,
            I => \N__46759\
        );

    \I__10500\ : Span4Mux_v
    port map (
            O => \N__46865\,
            I => \N__46759\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__46862\,
            I => \N__46759\
        );

    \I__10498\ : InMux
    port map (
            O => \N__46861\,
            I => \N__46756\
        );

    \I__10497\ : Span4Mux_h
    port map (
            O => \N__46858\,
            I => \N__46747\
        );

    \I__10496\ : Span4Mux_v
    port map (
            O => \N__46853\,
            I => \N__46747\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__46850\,
            I => \N__46747\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__46845\,
            I => \N__46747\
        );

    \I__10493\ : Span4Mux_h
    port map (
            O => \N__46842\,
            I => \N__46738\
        );

    \I__10492\ : Span4Mux_v
    port map (
            O => \N__46835\,
            I => \N__46738\
        );

    \I__10491\ : Span4Mux_h
    port map (
            O => \N__46832\,
            I => \N__46738\
        );

    \I__10490\ : Span4Mux_h
    port map (
            O => \N__46823\,
            I => \N__46738\
        );

    \I__10489\ : Span4Mux_h
    port map (
            O => \N__46820\,
            I => \N__46733\
        );

    \I__10488\ : Span4Mux_v
    port map (
            O => \N__46811\,
            I => \N__46733\
        );

    \I__10487\ : Span4Mux_h
    port map (
            O => \N__46808\,
            I => \N__46726\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__46805\,
            I => \N__46726\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__46802\,
            I => \N__46726\
        );

    \I__10484\ : Span4Mux_v
    port map (
            O => \N__46795\,
            I => \N__46723\
        );

    \I__10483\ : InMux
    port map (
            O => \N__46794\,
            I => \N__46720\
        );

    \I__10482\ : InMux
    port map (
            O => \N__46793\,
            I => \N__46717\
        );

    \I__10481\ : Span4Mux_h
    port map (
            O => \N__46788\,
            I => \N__46702\
        );

    \I__10480\ : LocalMux
    port map (
            O => \N__46785\,
            I => \N__46702\
        );

    \I__10479\ : LocalMux
    port map (
            O => \N__46782\,
            I => \N__46702\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__46779\,
            I => \N__46702\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__46776\,
            I => \N__46702\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__46773\,
            I => \N__46702\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__46770\,
            I => \N__46702\
        );

    \I__10474\ : InMux
    port map (
            O => \N__46769\,
            I => \N__46699\
        );

    \I__10473\ : Span4Mux_v
    port map (
            O => \N__46766\,
            I => \N__46690\
        );

    \I__10472\ : Span4Mux_h
    port map (
            O => \N__46759\,
            I => \N__46690\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__46756\,
            I => \N__46690\
        );

    \I__10470\ : Span4Mux_v
    port map (
            O => \N__46747\,
            I => \N__46690\
        );

    \I__10469\ : Span4Mux_v
    port map (
            O => \N__46738\,
            I => \N__46687\
        );

    \I__10468\ : Span4Mux_v
    port map (
            O => \N__46733\,
            I => \N__46676\
        );

    \I__10467\ : Span4Mux_v
    port map (
            O => \N__46726\,
            I => \N__46676\
        );

    \I__10466\ : Span4Mux_h
    port map (
            O => \N__46723\,
            I => \N__46676\
        );

    \I__10465\ : LocalMux
    port map (
            O => \N__46720\,
            I => \N__46676\
        );

    \I__10464\ : LocalMux
    port map (
            O => \N__46717\,
            I => \N__46676\
        );

    \I__10463\ : Span4Mux_v
    port map (
            O => \N__46702\,
            I => \N__46669\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__46699\,
            I => \N__46669\
        );

    \I__10461\ : Span4Mux_v
    port map (
            O => \N__46690\,
            I => \N__46669\
        );

    \I__10460\ : Odrv4
    port map (
            O => \N__46687\,
            I => spi_data_mosi_5
        );

    \I__10459\ : Odrv4
    port map (
            O => \N__46676\,
            I => spi_data_mosi_5
        );

    \I__10458\ : Odrv4
    port map (
            O => \N__46669\,
            I => spi_data_mosi_5
        );

    \I__10457\ : InMux
    port map (
            O => \N__46662\,
            I => \N__46659\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__46659\,
            I => \N__46656\
        );

    \I__10455\ : Span4Mux_v
    port map (
            O => \N__46656\,
            I => \N__46653\
        );

    \I__10454\ : Odrv4
    port map (
            O => \N__46653\,
            I => \sDAC_mem_9Z0Z_5\
        );

    \I__10453\ : InMux
    port map (
            O => \N__46650\,
            I => \N__46647\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__46647\,
            I => \N__46644\
        );

    \I__10451\ : Span4Mux_h
    port map (
            O => \N__46644\,
            I => \N__46641\
        );

    \I__10450\ : Span4Mux_h
    port map (
            O => \N__46641\,
            I => \N__46638\
        );

    \I__10449\ : Odrv4
    port map (
            O => \N__46638\,
            I => \sDAC_mem_9Z0Z_6\
        );

    \I__10448\ : CEMux
    port map (
            O => \N__46635\,
            I => \N__46632\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__46632\,
            I => \N__46626\
        );

    \I__10446\ : CEMux
    port map (
            O => \N__46631\,
            I => \N__46623\
        );

    \I__10445\ : CEMux
    port map (
            O => \N__46630\,
            I => \N__46620\
        );

    \I__10444\ : CEMux
    port map (
            O => \N__46629\,
            I => \N__46617\
        );

    \I__10443\ : Span4Mux_v
    port map (
            O => \N__46626\,
            I => \N__46614\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__46623\,
            I => \N__46611\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__46620\,
            I => \N__46608\
        );

    \I__10440\ : LocalMux
    port map (
            O => \N__46617\,
            I => \N__46605\
        );

    \I__10439\ : Span4Mux_h
    port map (
            O => \N__46614\,
            I => \N__46598\
        );

    \I__10438\ : Span4Mux_v
    port map (
            O => \N__46611\,
            I => \N__46598\
        );

    \I__10437\ : Span4Mux_v
    port map (
            O => \N__46608\,
            I => \N__46598\
        );

    \I__10436\ : Span4Mux_h
    port map (
            O => \N__46605\,
            I => \N__46595\
        );

    \I__10435\ : Span4Mux_v
    port map (
            O => \N__46598\,
            I => \N__46590\
        );

    \I__10434\ : Span4Mux_h
    port map (
            O => \N__46595\,
            I => \N__46590\
        );

    \I__10433\ : Odrv4
    port map (
            O => \N__46590\,
            I => \sDAC_mem_16_1_sqmuxa\
        );

    \I__10432\ : InMux
    port map (
            O => \N__46587\,
            I => \N__46584\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__46584\,
            I => \N__46581\
        );

    \I__10430\ : Span12Mux_v
    port map (
            O => \N__46581\,
            I => \N__46578\
        );

    \I__10429\ : Odrv12
    port map (
            O => \N__46578\,
            I => \sEEDACZ0Z_7\
        );

    \I__10428\ : CascadeMux
    port map (
            O => \N__46575\,
            I => \N__46570\
        );

    \I__10427\ : InMux
    port map (
            O => \N__46574\,
            I => \N__46560\
        );

    \I__10426\ : InMux
    port map (
            O => \N__46573\,
            I => \N__46556\
        );

    \I__10425\ : InMux
    port map (
            O => \N__46570\,
            I => \N__46551\
        );

    \I__10424\ : InMux
    port map (
            O => \N__46569\,
            I => \N__46551\
        );

    \I__10423\ : InMux
    port map (
            O => \N__46568\,
            I => \N__46538\
        );

    \I__10422\ : InMux
    port map (
            O => \N__46567\,
            I => \N__46538\
        );

    \I__10421\ : InMux
    port map (
            O => \N__46566\,
            I => \N__46538\
        );

    \I__10420\ : InMux
    port map (
            O => \N__46565\,
            I => \N__46538\
        );

    \I__10419\ : InMux
    port map (
            O => \N__46564\,
            I => \N__46538\
        );

    \I__10418\ : InMux
    port map (
            O => \N__46563\,
            I => \N__46538\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__46560\,
            I => \N__46535\
        );

    \I__10416\ : InMux
    port map (
            O => \N__46559\,
            I => \N__46532\
        );

    \I__10415\ : LocalMux
    port map (
            O => \N__46556\,
            I => \N__46529\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__46551\,
            I => \N__46525\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__46538\,
            I => \N__46522\
        );

    \I__10412\ : Span4Mux_v
    port map (
            O => \N__46535\,
            I => \N__46519\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__46532\,
            I => \N__46514\
        );

    \I__10410\ : Span4Mux_v
    port map (
            O => \N__46529\,
            I => \N__46514\
        );

    \I__10409\ : InMux
    port map (
            O => \N__46528\,
            I => \N__46508\
        );

    \I__10408\ : Span4Mux_h
    port map (
            O => \N__46525\,
            I => \N__46505\
        );

    \I__10407\ : Span4Mux_h
    port map (
            O => \N__46522\,
            I => \N__46502\
        );

    \I__10406\ : Span4Mux_v
    port map (
            O => \N__46519\,
            I => \N__46497\
        );

    \I__10405\ : Span4Mux_h
    port map (
            O => \N__46514\,
            I => \N__46497\
        );

    \I__10404\ : InMux
    port map (
            O => \N__46513\,
            I => \N__46490\
        );

    \I__10403\ : InMux
    port map (
            O => \N__46512\,
            I => \N__46490\
        );

    \I__10402\ : InMux
    port map (
            O => \N__46511\,
            I => \N__46490\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__46508\,
            I => \N__46487\
        );

    \I__10400\ : Span4Mux_h
    port map (
            O => \N__46505\,
            I => \N__46482\
        );

    \I__10399\ : Span4Mux_h
    port map (
            O => \N__46502\,
            I => \N__46479\
        );

    \I__10398\ : Span4Mux_h
    port map (
            O => \N__46497\,
            I => \N__46474\
        );

    \I__10397\ : LocalMux
    port map (
            O => \N__46490\,
            I => \N__46474\
        );

    \I__10396\ : Span12Mux_v
    port map (
            O => \N__46487\,
            I => \N__46471\
        );

    \I__10395\ : InMux
    port map (
            O => \N__46486\,
            I => \N__46468\
        );

    \I__10394\ : InMux
    port map (
            O => \N__46485\,
            I => \N__46465\
        );

    \I__10393\ : Odrv4
    port map (
            O => \N__46482\,
            I => \sAddressZ0Z_5\
        );

    \I__10392\ : Odrv4
    port map (
            O => \N__46479\,
            I => \sAddressZ0Z_5\
        );

    \I__10391\ : Odrv4
    port map (
            O => \N__46474\,
            I => \sAddressZ0Z_5\
        );

    \I__10390\ : Odrv12
    port map (
            O => \N__46471\,
            I => \sAddressZ0Z_5\
        );

    \I__10389\ : LocalMux
    port map (
            O => \N__46468\,
            I => \sAddressZ0Z_5\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__46465\,
            I => \sAddressZ0Z_5\
        );

    \I__10387\ : CascadeMux
    port map (
            O => \N__46452\,
            I => \N__46446\
        );

    \I__10386\ : InMux
    port map (
            O => \N__46451\,
            I => \N__46442\
        );

    \I__10385\ : CascadeMux
    port map (
            O => \N__46450\,
            I => \N__46439\
        );

    \I__10384\ : CascadeMux
    port map (
            O => \N__46449\,
            I => \N__46435\
        );

    \I__10383\ : InMux
    port map (
            O => \N__46446\,
            I => \N__46432\
        );

    \I__10382\ : CascadeMux
    port map (
            O => \N__46445\,
            I => \N__46429\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__46442\,
            I => \N__46425\
        );

    \I__10380\ : InMux
    port map (
            O => \N__46439\,
            I => \N__46422\
        );

    \I__10379\ : InMux
    port map (
            O => \N__46438\,
            I => \N__46419\
        );

    \I__10378\ : InMux
    port map (
            O => \N__46435\,
            I => \N__46415\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__46432\,
            I => \N__46409\
        );

    \I__10376\ : InMux
    port map (
            O => \N__46429\,
            I => \N__46406\
        );

    \I__10375\ : InMux
    port map (
            O => \N__46428\,
            I => \N__46403\
        );

    \I__10374\ : Span4Mux_v
    port map (
            O => \N__46425\,
            I => \N__46398\
        );

    \I__10373\ : LocalMux
    port map (
            O => \N__46422\,
            I => \N__46398\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__46419\,
            I => \N__46395\
        );

    \I__10371\ : InMux
    port map (
            O => \N__46418\,
            I => \N__46392\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__46415\,
            I => \N__46389\
        );

    \I__10369\ : InMux
    port map (
            O => \N__46414\,
            I => \N__46382\
        );

    \I__10368\ : InMux
    port map (
            O => \N__46413\,
            I => \N__46382\
        );

    \I__10367\ : InMux
    port map (
            O => \N__46412\,
            I => \N__46382\
        );

    \I__10366\ : Span4Mux_h
    port map (
            O => \N__46409\,
            I => \N__46379\
        );

    \I__10365\ : LocalMux
    port map (
            O => \N__46406\,
            I => \N__46376\
        );

    \I__10364\ : LocalMux
    port map (
            O => \N__46403\,
            I => \N__46373\
        );

    \I__10363\ : Span4Mux_h
    port map (
            O => \N__46398\,
            I => \N__46368\
        );

    \I__10362\ : Span4Mux_v
    port map (
            O => \N__46395\,
            I => \N__46368\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__46392\,
            I => \N__46365\
        );

    \I__10360\ : Span4Mux_h
    port map (
            O => \N__46389\,
            I => \N__46362\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__46382\,
            I => \N__46359\
        );

    \I__10358\ : Span4Mux_v
    port map (
            O => \N__46379\,
            I => \N__46354\
        );

    \I__10357\ : Span4Mux_h
    port map (
            O => \N__46376\,
            I => \N__46354\
        );

    \I__10356\ : Span4Mux_v
    port map (
            O => \N__46373\,
            I => \N__46351\
        );

    \I__10355\ : Span4Mux_v
    port map (
            O => \N__46368\,
            I => \N__46348\
        );

    \I__10354\ : Span4Mux_h
    port map (
            O => \N__46365\,
            I => \N__46341\
        );

    \I__10353\ : Span4Mux_v
    port map (
            O => \N__46362\,
            I => \N__46341\
        );

    \I__10352\ : Span4Mux_h
    port map (
            O => \N__46359\,
            I => \N__46341\
        );

    \I__10351\ : Span4Mux_v
    port map (
            O => \N__46354\,
            I => \N__46334\
        );

    \I__10350\ : Span4Mux_h
    port map (
            O => \N__46351\,
            I => \N__46334\
        );

    \I__10349\ : Span4Mux_h
    port map (
            O => \N__46348\,
            I => \N__46334\
        );

    \I__10348\ : Odrv4
    port map (
            O => \N__46341\,
            I => \N_139\
        );

    \I__10347\ : Odrv4
    port map (
            O => \N__46334\,
            I => \N_139\
        );

    \I__10346\ : InMux
    port map (
            O => \N__46329\,
            I => \N__46323\
        );

    \I__10345\ : InMux
    port map (
            O => \N__46328\,
            I => \N__46323\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__46323\,
            I => \N__46316\
        );

    \I__10343\ : InMux
    port map (
            O => \N__46322\,
            I => \N__46313\
        );

    \I__10342\ : InMux
    port map (
            O => \N__46321\,
            I => \N__46308\
        );

    \I__10341\ : InMux
    port map (
            O => \N__46320\,
            I => \N__46308\
        );

    \I__10340\ : InMux
    port map (
            O => \N__46319\,
            I => \N__46305\
        );

    \I__10339\ : Span4Mux_h
    port map (
            O => \N__46316\,
            I => \N__46302\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__46313\,
            I => \N__46297\
        );

    \I__10337\ : LocalMux
    port map (
            O => \N__46308\,
            I => \N__46297\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__46305\,
            I => \N__46289\
        );

    \I__10335\ : Span4Mux_h
    port map (
            O => \N__46302\,
            I => \N__46286\
        );

    \I__10334\ : Span4Mux_h
    port map (
            O => \N__46297\,
            I => \N__46283\
        );

    \I__10333\ : InMux
    port map (
            O => \N__46296\,
            I => \N__46272\
        );

    \I__10332\ : InMux
    port map (
            O => \N__46295\,
            I => \N__46272\
        );

    \I__10331\ : InMux
    port map (
            O => \N__46294\,
            I => \N__46272\
        );

    \I__10330\ : InMux
    port map (
            O => \N__46293\,
            I => \N__46272\
        );

    \I__10329\ : InMux
    port map (
            O => \N__46292\,
            I => \N__46272\
        );

    \I__10328\ : Odrv4
    port map (
            O => \N__46289\,
            I => \N_278\
        );

    \I__10327\ : Odrv4
    port map (
            O => \N__46286\,
            I => \N_278\
        );

    \I__10326\ : Odrv4
    port map (
            O => \N__46283\,
            I => \N_278\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__46272\,
            I => \N_278\
        );

    \I__10324\ : CEMux
    port map (
            O => \N__46263\,
            I => \N__46260\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__46260\,
            I => \N__46257\
        );

    \I__10322\ : Span4Mux_v
    port map (
            O => \N__46257\,
            I => \N__46254\
        );

    \I__10321\ : Odrv4
    port map (
            O => \N__46254\,
            I => \sDAC_mem_41_1_sqmuxa\
        );

    \I__10320\ : CascadeMux
    port map (
            O => \N__46251\,
            I => \N__46240\
        );

    \I__10319\ : InMux
    port map (
            O => \N__46250\,
            I => \N__46237\
        );

    \I__10318\ : InMux
    port map (
            O => \N__46249\,
            I => \N__46234\
        );

    \I__10317\ : InMux
    port map (
            O => \N__46248\,
            I => \N__46231\
        );

    \I__10316\ : CascadeMux
    port map (
            O => \N__46247\,
            I => \N__46228\
        );

    \I__10315\ : CascadeMux
    port map (
            O => \N__46246\,
            I => \N__46225\
        );

    \I__10314\ : CascadeMux
    port map (
            O => \N__46245\,
            I => \N__46222\
        );

    \I__10313\ : InMux
    port map (
            O => \N__46244\,
            I => \N__46217\
        );

    \I__10312\ : InMux
    port map (
            O => \N__46243\,
            I => \N__46217\
        );

    \I__10311\ : InMux
    port map (
            O => \N__46240\,
            I => \N__46214\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__46237\,
            I => \N__46211\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__46234\,
            I => \N__46208\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__46231\,
            I => \N__46204\
        );

    \I__10307\ : InMux
    port map (
            O => \N__46228\,
            I => \N__46201\
        );

    \I__10306\ : InMux
    port map (
            O => \N__46225\,
            I => \N__46196\
        );

    \I__10305\ : InMux
    port map (
            O => \N__46222\,
            I => \N__46196\
        );

    \I__10304\ : LocalMux
    port map (
            O => \N__46217\,
            I => \N__46193\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__46214\,
            I => \N__46190\
        );

    \I__10302\ : Span4Mux_h
    port map (
            O => \N__46211\,
            I => \N__46185\
        );

    \I__10301\ : Span4Mux_h
    port map (
            O => \N__46208\,
            I => \N__46185\
        );

    \I__10300\ : CascadeMux
    port map (
            O => \N__46207\,
            I => \N__46181\
        );

    \I__10299\ : Span4Mux_h
    port map (
            O => \N__46204\,
            I => \N__46176\
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__46201\,
            I => \N__46176\
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__46196\,
            I => \N__46173\
        );

    \I__10296\ : Span4Mux_h
    port map (
            O => \N__46193\,
            I => \N__46170\
        );

    \I__10295\ : Span4Mux_v
    port map (
            O => \N__46190\,
            I => \N__46165\
        );

    \I__10294\ : Span4Mux_v
    port map (
            O => \N__46185\,
            I => \N__46165\
        );

    \I__10293\ : InMux
    port map (
            O => \N__46184\,
            I => \N__46160\
        );

    \I__10292\ : InMux
    port map (
            O => \N__46181\,
            I => \N__46160\
        );

    \I__10291\ : Span4Mux_v
    port map (
            O => \N__46176\,
            I => \N__46157\
        );

    \I__10290\ : Span4Mux_v
    port map (
            O => \N__46173\,
            I => \N__46154\
        );

    \I__10289\ : Span4Mux_h
    port map (
            O => \N__46170\,
            I => \N__46151\
        );

    \I__10288\ : Span4Mux_h
    port map (
            O => \N__46165\,
            I => \N__46148\
        );

    \I__10287\ : LocalMux
    port map (
            O => \N__46160\,
            I => \N__46141\
        );

    \I__10286\ : Span4Mux_h
    port map (
            O => \N__46157\,
            I => \N__46141\
        );

    \I__10285\ : Span4Mux_v
    port map (
            O => \N__46154\,
            I => \N__46141\
        );

    \I__10284\ : Odrv4
    port map (
            O => \N__46151\,
            I => \N_285\
        );

    \I__10283\ : Odrv4
    port map (
            O => \N__46148\,
            I => \N_285\
        );

    \I__10282\ : Odrv4
    port map (
            O => \N__46141\,
            I => \N_285\
        );

    \I__10281\ : InMux
    port map (
            O => \N__46134\,
            I => \N__46129\
        );

    \I__10280\ : CascadeMux
    port map (
            O => \N__46133\,
            I => \N__46125\
        );

    \I__10279\ : InMux
    port map (
            O => \N__46132\,
            I => \N__46120\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__46129\,
            I => \N__46115\
        );

    \I__10277\ : InMux
    port map (
            O => \N__46128\,
            I => \N__46112\
        );

    \I__10276\ : InMux
    port map (
            O => \N__46125\,
            I => \N__46105\
        );

    \I__10275\ : InMux
    port map (
            O => \N__46124\,
            I => \N__46105\
        );

    \I__10274\ : InMux
    port map (
            O => \N__46123\,
            I => \N__46105\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__46120\,
            I => \N__46102\
        );

    \I__10272\ : InMux
    port map (
            O => \N__46119\,
            I => \N__46097\
        );

    \I__10271\ : InMux
    port map (
            O => \N__46118\,
            I => \N__46097\
        );

    \I__10270\ : Span4Mux_h
    port map (
            O => \N__46115\,
            I => \N__46093\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__46112\,
            I => \N__46088\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__46105\,
            I => \N__46088\
        );

    \I__10267\ : Span4Mux_v
    port map (
            O => \N__46102\,
            I => \N__46085\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__46097\,
            I => \N__46082\
        );

    \I__10265\ : InMux
    port map (
            O => \N__46096\,
            I => \N__46079\
        );

    \I__10264\ : Span4Mux_v
    port map (
            O => \N__46093\,
            I => \N__46074\
        );

    \I__10263\ : Span4Mux_v
    port map (
            O => \N__46088\,
            I => \N__46074\
        );

    \I__10262\ : Span4Mux_v
    port map (
            O => \N__46085\,
            I => \N__46069\
        );

    \I__10261\ : Span4Mux_h
    port map (
            O => \N__46082\,
            I => \N__46069\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__46079\,
            I => \N__46062\
        );

    \I__10259\ : Span4Mux_h
    port map (
            O => \N__46074\,
            I => \N__46062\
        );

    \I__10258\ : Span4Mux_h
    port map (
            O => \N__46069\,
            I => \N__46059\
        );

    \I__10257\ : InMux
    port map (
            O => \N__46068\,
            I => \N__46056\
        );

    \I__10256\ : InMux
    port map (
            O => \N__46067\,
            I => \N__46053\
        );

    \I__10255\ : Odrv4
    port map (
            O => \N__46062\,
            I => \N_1480\
        );

    \I__10254\ : Odrv4
    port map (
            O => \N__46059\,
            I => \N_1480\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__46056\,
            I => \N_1480\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__46053\,
            I => \N_1480\
        );

    \I__10251\ : InMux
    port map (
            O => \N__46044\,
            I => \N__46040\
        );

    \I__10250\ : InMux
    port map (
            O => \N__46043\,
            I => \N__46037\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__46040\,
            I => \N__46034\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__46037\,
            I => \N__46031\
        );

    \I__10247\ : Span4Mux_v
    port map (
            O => \N__46034\,
            I => \N__46028\
        );

    \I__10246\ : Span4Mux_h
    port map (
            O => \N__46031\,
            I => \N__46025\
        );

    \I__10245\ : Span4Mux_h
    port map (
            O => \N__46028\,
            I => \N__46020\
        );

    \I__10244\ : Span4Mux_h
    port map (
            O => \N__46025\,
            I => \N__46020\
        );

    \I__10243\ : Odrv4
    port map (
            O => \N__46020\,
            I => \N_360\
        );

    \I__10242\ : InMux
    port map (
            O => \N__46017\,
            I => \N__46014\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__46014\,
            I => \N__46011\
        );

    \I__10240\ : Span4Mux_v
    port map (
            O => \N__46011\,
            I => \N__46008\
        );

    \I__10239\ : Span4Mux_h
    port map (
            O => \N__46008\,
            I => \N__46005\
        );

    \I__10238\ : Odrv4
    port map (
            O => \N__46005\,
            I => \sEEDACZ0Z_0\
        );

    \I__10237\ : InMux
    port map (
            O => \N__46002\,
            I => \N__45999\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__45999\,
            I => \N__45996\
        );

    \I__10235\ : Span4Mux_v
    port map (
            O => \N__45996\,
            I => \N__45993\
        );

    \I__10234\ : Odrv4
    port map (
            O => \N__45993\,
            I => \sEEDACZ0Z_1\
        );

    \I__10233\ : InMux
    port map (
            O => \N__45990\,
            I => \N__45987\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__45987\,
            I => \N__45984\
        );

    \I__10231\ : Span4Mux_h
    port map (
            O => \N__45984\,
            I => \N__45981\
        );

    \I__10230\ : Span4Mux_h
    port map (
            O => \N__45981\,
            I => \N__45978\
        );

    \I__10229\ : Odrv4
    port map (
            O => \N__45978\,
            I => \sEEDACZ0Z_2\
        );

    \I__10228\ : InMux
    port map (
            O => \N__45975\,
            I => \N__45972\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__45972\,
            I => \N__45969\
        );

    \I__10226\ : Span4Mux_v
    port map (
            O => \N__45969\,
            I => \N__45966\
        );

    \I__10225\ : Sp12to4
    port map (
            O => \N__45966\,
            I => \N__45963\
        );

    \I__10224\ : Odrv12
    port map (
            O => \N__45963\,
            I => \sEEDACZ0Z_3\
        );

    \I__10223\ : InMux
    port map (
            O => \N__45960\,
            I => \N__45957\
        );

    \I__10222\ : LocalMux
    port map (
            O => \N__45957\,
            I => \N__45954\
        );

    \I__10221\ : Span4Mux_h
    port map (
            O => \N__45954\,
            I => \N__45951\
        );

    \I__10220\ : Span4Mux_h
    port map (
            O => \N__45951\,
            I => \N__45948\
        );

    \I__10219\ : Odrv4
    port map (
            O => \N__45948\,
            I => \sEEDACZ0Z_4\
        );

    \I__10218\ : CascadeMux
    port map (
            O => \N__45945\,
            I => \N__45939\
        );

    \I__10217\ : CascadeMux
    port map (
            O => \N__45944\,
            I => \N__45935\
        );

    \I__10216\ : InMux
    port map (
            O => \N__45943\,
            I => \N__45922\
        );

    \I__10215\ : InMux
    port map (
            O => \N__45942\,
            I => \N__45922\
        );

    \I__10214\ : InMux
    port map (
            O => \N__45939\,
            I => \N__45922\
        );

    \I__10213\ : InMux
    port map (
            O => \N__45938\,
            I => \N__45922\
        );

    \I__10212\ : InMux
    port map (
            O => \N__45935\,
            I => \N__45919\
        );

    \I__10211\ : InMux
    port map (
            O => \N__45934\,
            I => \N__45912\
        );

    \I__10210\ : InMux
    port map (
            O => \N__45933\,
            I => \N__45912\
        );

    \I__10209\ : InMux
    port map (
            O => \N__45932\,
            I => \N__45912\
        );

    \I__10208\ : InMux
    port map (
            O => \N__45931\,
            I => \N__45905\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__45922\,
            I => \N__45902\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__45919\,
            I => \N__45897\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__45912\,
            I => \N__45897\
        );

    \I__10204\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45892\
        );

    \I__10203\ : InMux
    port map (
            O => \N__45910\,
            I => \N__45892\
        );

    \I__10202\ : CascadeMux
    port map (
            O => \N__45909\,
            I => \N__45884\
        );

    \I__10201\ : CascadeMux
    port map (
            O => \N__45908\,
            I => \N__45862\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__45905\,
            I => \N__45856\
        );

    \I__10199\ : Span4Mux_h
    port map (
            O => \N__45902\,
            I => \N__45849\
        );

    \I__10198\ : Span4Mux_v
    port map (
            O => \N__45897\,
            I => \N__45849\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__45892\,
            I => \N__45849\
        );

    \I__10196\ : InMux
    port map (
            O => \N__45891\,
            I => \N__45842\
        );

    \I__10195\ : InMux
    port map (
            O => \N__45890\,
            I => \N__45842\
        );

    \I__10194\ : InMux
    port map (
            O => \N__45889\,
            I => \N__45838\
        );

    \I__10193\ : InMux
    port map (
            O => \N__45888\,
            I => \N__45829\
        );

    \I__10192\ : InMux
    port map (
            O => \N__45887\,
            I => \N__45829\
        );

    \I__10191\ : InMux
    port map (
            O => \N__45884\,
            I => \N__45829\
        );

    \I__10190\ : InMux
    port map (
            O => \N__45883\,
            I => \N__45829\
        );

    \I__10189\ : CascadeMux
    port map (
            O => \N__45882\,
            I => \N__45825\
        );

    \I__10188\ : InMux
    port map (
            O => \N__45881\,
            I => \N__45822\
        );

    \I__10187\ : InMux
    port map (
            O => \N__45880\,
            I => \N__45817\
        );

    \I__10186\ : InMux
    port map (
            O => \N__45879\,
            I => \N__45817\
        );

    \I__10185\ : InMux
    port map (
            O => \N__45878\,
            I => \N__45814\
        );

    \I__10184\ : InMux
    port map (
            O => \N__45877\,
            I => \N__45809\
        );

    \I__10183\ : InMux
    port map (
            O => \N__45876\,
            I => \N__45809\
        );

    \I__10182\ : CascadeMux
    port map (
            O => \N__45875\,
            I => \N__45804\
        );

    \I__10181\ : InMux
    port map (
            O => \N__45874\,
            I => \N__45800\
        );

    \I__10180\ : InMux
    port map (
            O => \N__45873\,
            I => \N__45796\
        );

    \I__10179\ : InMux
    port map (
            O => \N__45872\,
            I => \N__45793\
        );

    \I__10178\ : InMux
    port map (
            O => \N__45871\,
            I => \N__45784\
        );

    \I__10177\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45784\
        );

    \I__10176\ : InMux
    port map (
            O => \N__45869\,
            I => \N__45784\
        );

    \I__10175\ : InMux
    port map (
            O => \N__45868\,
            I => \N__45784\
        );

    \I__10174\ : InMux
    port map (
            O => \N__45867\,
            I => \N__45780\
        );

    \I__10173\ : InMux
    port map (
            O => \N__45866\,
            I => \N__45777\
        );

    \I__10172\ : InMux
    port map (
            O => \N__45865\,
            I => \N__45770\
        );

    \I__10171\ : InMux
    port map (
            O => \N__45862\,
            I => \N__45770\
        );

    \I__10170\ : InMux
    port map (
            O => \N__45861\,
            I => \N__45770\
        );

    \I__10169\ : InMux
    port map (
            O => \N__45860\,
            I => \N__45765\
        );

    \I__10168\ : InMux
    port map (
            O => \N__45859\,
            I => \N__45765\
        );

    \I__10167\ : Span4Mux_v
    port map (
            O => \N__45856\,
            I => \N__45760\
        );

    \I__10166\ : Span4Mux_v
    port map (
            O => \N__45849\,
            I => \N__45760\
        );

    \I__10165\ : InMux
    port map (
            O => \N__45848\,
            I => \N__45755\
        );

    \I__10164\ : InMux
    port map (
            O => \N__45847\,
            I => \N__45755\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__45842\,
            I => \N__45752\
        );

    \I__10162\ : CascadeMux
    port map (
            O => \N__45841\,
            I => \N__45747\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__45838\,
            I => \N__45741\
        );

    \I__10160\ : LocalMux
    port map (
            O => \N__45829\,
            I => \N__45741\
        );

    \I__10159\ : InMux
    port map (
            O => \N__45828\,
            I => \N__45738\
        );

    \I__10158\ : InMux
    port map (
            O => \N__45825\,
            I => \N__45731\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__45822\,
            I => \N__45723\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__45817\,
            I => \N__45723\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__45814\,
            I => \N__45718\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__45809\,
            I => \N__45718\
        );

    \I__10153\ : CascadeMux
    port map (
            O => \N__45808\,
            I => \N__45713\
        );

    \I__10152\ : CascadeMux
    port map (
            O => \N__45807\,
            I => \N__45706\
        );

    \I__10151\ : InMux
    port map (
            O => \N__45804\,
            I => \N__45701\
        );

    \I__10150\ : InMux
    port map (
            O => \N__45803\,
            I => \N__45701\
        );

    \I__10149\ : LocalMux
    port map (
            O => \N__45800\,
            I => \N__45698\
        );

    \I__10148\ : InMux
    port map (
            O => \N__45799\,
            I => \N__45695\
        );

    \I__10147\ : LocalMux
    port map (
            O => \N__45796\,
            I => \N__45690\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__45793\,
            I => \N__45690\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__45784\,
            I => \N__45687\
        );

    \I__10144\ : InMux
    port map (
            O => \N__45783\,
            I => \N__45684\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__45780\,
            I => \N__45681\
        );

    \I__10142\ : LocalMux
    port map (
            O => \N__45777\,
            I => \N__45676\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__45770\,
            I => \N__45676\
        );

    \I__10140\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45667\
        );

    \I__10139\ : Span4Mux_h
    port map (
            O => \N__45760\,
            I => \N__45667\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__45755\,
            I => \N__45667\
        );

    \I__10137\ : Span4Mux_h
    port map (
            O => \N__45752\,
            I => \N__45667\
        );

    \I__10136\ : InMux
    port map (
            O => \N__45751\,
            I => \N__45664\
        );

    \I__10135\ : InMux
    port map (
            O => \N__45750\,
            I => \N__45661\
        );

    \I__10134\ : InMux
    port map (
            O => \N__45747\,
            I => \N__45656\
        );

    \I__10133\ : InMux
    port map (
            O => \N__45746\,
            I => \N__45656\
        );

    \I__10132\ : Span4Mux_h
    port map (
            O => \N__45741\,
            I => \N__45651\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__45738\,
            I => \N__45651\
        );

    \I__10130\ : InMux
    port map (
            O => \N__45737\,
            I => \N__45648\
        );

    \I__10129\ : InMux
    port map (
            O => \N__45736\,
            I => \N__45645\
        );

    \I__10128\ : InMux
    port map (
            O => \N__45735\,
            I => \N__45640\
        );

    \I__10127\ : InMux
    port map (
            O => \N__45734\,
            I => \N__45640\
        );

    \I__10126\ : LocalMux
    port map (
            O => \N__45731\,
            I => \N__45636\
        );

    \I__10125\ : InMux
    port map (
            O => \N__45730\,
            I => \N__45629\
        );

    \I__10124\ : InMux
    port map (
            O => \N__45729\,
            I => \N__45629\
        );

    \I__10123\ : InMux
    port map (
            O => \N__45728\,
            I => \N__45629\
        );

    \I__10122\ : Span4Mux_h
    port map (
            O => \N__45723\,
            I => \N__45624\
        );

    \I__10121\ : Span4Mux_v
    port map (
            O => \N__45718\,
            I => \N__45624\
        );

    \I__10120\ : InMux
    port map (
            O => \N__45717\,
            I => \N__45621\
        );

    \I__10119\ : InMux
    port map (
            O => \N__45716\,
            I => \N__45618\
        );

    \I__10118\ : InMux
    port map (
            O => \N__45713\,
            I => \N__45611\
        );

    \I__10117\ : InMux
    port map (
            O => \N__45712\,
            I => \N__45611\
        );

    \I__10116\ : InMux
    port map (
            O => \N__45711\,
            I => \N__45611\
        );

    \I__10115\ : InMux
    port map (
            O => \N__45710\,
            I => \N__45606\
        );

    \I__10114\ : InMux
    port map (
            O => \N__45709\,
            I => \N__45606\
        );

    \I__10113\ : InMux
    port map (
            O => \N__45706\,
            I => \N__45603\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__45701\,
            I => \N__45596\
        );

    \I__10111\ : Span4Mux_h
    port map (
            O => \N__45698\,
            I => \N__45596\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__45695\,
            I => \N__45596\
        );

    \I__10109\ : Span4Mux_h
    port map (
            O => \N__45690\,
            I => \N__45591\
        );

    \I__10108\ : Span4Mux_v
    port map (
            O => \N__45687\,
            I => \N__45591\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__45684\,
            I => \N__45582\
        );

    \I__10106\ : Span4Mux_h
    port map (
            O => \N__45681\,
            I => \N__45582\
        );

    \I__10105\ : Span4Mux_h
    port map (
            O => \N__45676\,
            I => \N__45582\
        );

    \I__10104\ : Span4Mux_v
    port map (
            O => \N__45667\,
            I => \N__45582\
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__45664\,
            I => \N__45567\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__45661\,
            I => \N__45567\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__45656\,
            I => \N__45567\
        );

    \I__10100\ : Sp12to4
    port map (
            O => \N__45651\,
            I => \N__45567\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__45648\,
            I => \N__45567\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__45645\,
            I => \N__45567\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__45640\,
            I => \N__45567\
        );

    \I__10096\ : InMux
    port map (
            O => \N__45639\,
            I => \N__45564\
        );

    \I__10095\ : Span4Mux_h
    port map (
            O => \N__45636\,
            I => \N__45557\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__45629\,
            I => \N__45557\
        );

    \I__10093\ : Span4Mux_v
    port map (
            O => \N__45624\,
            I => \N__45557\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__45621\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__45618\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__45611\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__45606\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__45603\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__10087\ : Odrv4
    port map (
            O => \N__45596\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__10086\ : Odrv4
    port map (
            O => \N__45591\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__10085\ : Odrv4
    port map (
            O => \N__45582\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__10084\ : Odrv12
    port map (
            O => \N__45567\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__45564\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__10082\ : Odrv4
    port map (
            O => \N__45557\,
            I => \sDAC_mem_pointerZ0Z_2\
        );

    \I__10081\ : CascadeMux
    port map (
            O => \N__45534\,
            I => \N__45530\
        );

    \I__10080\ : InMux
    port map (
            O => \N__45533\,
            I => \N__45515\
        );

    \I__10079\ : InMux
    port map (
            O => \N__45530\,
            I => \N__45512\
        );

    \I__10078\ : InMux
    port map (
            O => \N__45529\,
            I => \N__45507\
        );

    \I__10077\ : InMux
    port map (
            O => \N__45528\,
            I => \N__45507\
        );

    \I__10076\ : InMux
    port map (
            O => \N__45527\,
            I => \N__45502\
        );

    \I__10075\ : InMux
    port map (
            O => \N__45526\,
            I => \N__45502\
        );

    \I__10074\ : InMux
    port map (
            O => \N__45525\,
            I => \N__45496\
        );

    \I__10073\ : InMux
    port map (
            O => \N__45524\,
            I => \N__45496\
        );

    \I__10072\ : InMux
    port map (
            O => \N__45523\,
            I => \N__45487\
        );

    \I__10071\ : InMux
    port map (
            O => \N__45522\,
            I => \N__45482\
        );

    \I__10070\ : InMux
    port map (
            O => \N__45521\,
            I => \N__45482\
        );

    \I__10069\ : InMux
    port map (
            O => \N__45520\,
            I => \N__45477\
        );

    \I__10068\ : InMux
    port map (
            O => \N__45519\,
            I => \N__45472\
        );

    \I__10067\ : InMux
    port map (
            O => \N__45518\,
            I => \N__45472\
        );

    \I__10066\ : LocalMux
    port map (
            O => \N__45515\,
            I => \N__45465\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__45512\,
            I => \N__45465\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__45507\,
            I => \N__45465\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__45502\,
            I => \N__45462\
        );

    \I__10062\ : InMux
    port map (
            O => \N__45501\,
            I => \N__45459\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__45496\,
            I => \N__45454\
        );

    \I__10060\ : InMux
    port map (
            O => \N__45495\,
            I => \N__45449\
        );

    \I__10059\ : InMux
    port map (
            O => \N__45494\,
            I => \N__45449\
        );

    \I__10058\ : InMux
    port map (
            O => \N__45493\,
            I => \N__45444\
        );

    \I__10057\ : InMux
    port map (
            O => \N__45492\,
            I => \N__45444\
        );

    \I__10056\ : CascadeMux
    port map (
            O => \N__45491\,
            I => \N__45441\
        );

    \I__10055\ : InMux
    port map (
            O => \N__45490\,
            I => \N__45436\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__45487\,
            I => \N__45433\
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__45482\,
            I => \N__45430\
        );

    \I__10052\ : InMux
    port map (
            O => \N__45481\,
            I => \N__45425\
        );

    \I__10051\ : InMux
    port map (
            O => \N__45480\,
            I => \N__45425\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__45477\,
            I => \N__45416\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__45472\,
            I => \N__45416\
        );

    \I__10048\ : Span4Mux_v
    port map (
            O => \N__45465\,
            I => \N__45411\
        );

    \I__10047\ : Span4Mux_v
    port map (
            O => \N__45462\,
            I => \N__45406\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__45459\,
            I => \N__45406\
        );

    \I__10045\ : InMux
    port map (
            O => \N__45458\,
            I => \N__45401\
        );

    \I__10044\ : InMux
    port map (
            O => \N__45457\,
            I => \N__45401\
        );

    \I__10043\ : Span4Mux_v
    port map (
            O => \N__45454\,
            I => \N__45396\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__45449\,
            I => \N__45396\
        );

    \I__10041\ : LocalMux
    port map (
            O => \N__45444\,
            I => \N__45393\
        );

    \I__10040\ : InMux
    port map (
            O => \N__45441\,
            I => \N__45390\
        );

    \I__10039\ : InMux
    port map (
            O => \N__45440\,
            I => \N__45387\
        );

    \I__10038\ : InMux
    port map (
            O => \N__45439\,
            I => \N__45384\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__45436\,
            I => \N__45381\
        );

    \I__10036\ : Span4Mux_v
    port map (
            O => \N__45433\,
            I => \N__45374\
        );

    \I__10035\ : Span4Mux_h
    port map (
            O => \N__45430\,
            I => \N__45374\
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__45425\,
            I => \N__45374\
        );

    \I__10033\ : InMux
    port map (
            O => \N__45424\,
            I => \N__45369\
        );

    \I__10032\ : InMux
    port map (
            O => \N__45423\,
            I => \N__45366\
        );

    \I__10031\ : InMux
    port map (
            O => \N__45422\,
            I => \N__45361\
        );

    \I__10030\ : InMux
    port map (
            O => \N__45421\,
            I => \N__45361\
        );

    \I__10029\ : Span4Mux_v
    port map (
            O => \N__45416\,
            I => \N__45358\
        );

    \I__10028\ : InMux
    port map (
            O => \N__45415\,
            I => \N__45353\
        );

    \I__10027\ : InMux
    port map (
            O => \N__45414\,
            I => \N__45353\
        );

    \I__10026\ : Span4Mux_h
    port map (
            O => \N__45411\,
            I => \N__45348\
        );

    \I__10025\ : Span4Mux_v
    port map (
            O => \N__45406\,
            I => \N__45348\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__45401\,
            I => \N__45341\
        );

    \I__10023\ : Span4Mux_v
    port map (
            O => \N__45396\,
            I => \N__45341\
        );

    \I__10022\ : Span4Mux_v
    port map (
            O => \N__45393\,
            I => \N__45341\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__45390\,
            I => \N__45334\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__45387\,
            I => \N__45334\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__45384\,
            I => \N__45334\
        );

    \I__10018\ : Span4Mux_v
    port map (
            O => \N__45381\,
            I => \N__45329\
        );

    \I__10017\ : Span4Mux_v
    port map (
            O => \N__45374\,
            I => \N__45329\
        );

    \I__10016\ : InMux
    port map (
            O => \N__45373\,
            I => \N__45324\
        );

    \I__10015\ : InMux
    port map (
            O => \N__45372\,
            I => \N__45324\
        );

    \I__10014\ : LocalMux
    port map (
            O => \N__45369\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__45366\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__45361\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__45358\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__45353\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__10009\ : Odrv4
    port map (
            O => \N__45348\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__10008\ : Odrv4
    port map (
            O => \N__45341\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__10007\ : Odrv12
    port map (
            O => \N__45334\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__10006\ : Odrv4
    port map (
            O => \N__45329\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__45324\,
            I => \sDAC_mem_pointerZ0Z_1\
        );

    \I__10004\ : CascadeMux
    port map (
            O => \N__45303\,
            I => \sDAC_data_RNO_18Z0Z_4_cascade_\
        );

    \I__10003\ : InMux
    port map (
            O => \N__45300\,
            I => \N__45297\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__45297\,
            I => \sDAC_data_2_24_ns_1_4\
        );

    \I__10001\ : InMux
    port map (
            O => \N__45294\,
            I => \N__45291\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__45291\,
            I => \sDAC_mem_12Z0Z_0\
        );

    \I__9999\ : InMux
    port map (
            O => \N__45288\,
            I => \N__45285\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__45285\,
            I => \N__45282\
        );

    \I__9997\ : Odrv4
    port map (
            O => \N__45282\,
            I => \sDAC_mem_15Z0Z_1\
        );

    \I__9996\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45276\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__45276\,
            I => \sDAC_mem_14Z0Z_1\
        );

    \I__9994\ : InMux
    port map (
            O => \N__45273\,
            I => \N__45270\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__45270\,
            I => \sDAC_data_RNO_19Z0Z_4\
        );

    \I__9992\ : InMux
    port map (
            O => \N__45267\,
            I => \N__45264\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__45264\,
            I => \sDAC_mem_12Z0Z_1\
        );

    \I__9990\ : InMux
    port map (
            O => \N__45261\,
            I => \N__45258\
        );

    \I__9989\ : LocalMux
    port map (
            O => \N__45258\,
            I => \N__45255\
        );

    \I__9988\ : Span4Mux_v
    port map (
            O => \N__45255\,
            I => \N__45252\
        );

    \I__9987\ : Span4Mux_h
    port map (
            O => \N__45252\,
            I => \N__45249\
        );

    \I__9986\ : Odrv4
    port map (
            O => \N__45249\,
            I => \sDAC_mem_27Z0Z_0\
        );

    \I__9985\ : CEMux
    port map (
            O => \N__45246\,
            I => \N__45242\
        );

    \I__9984\ : CEMux
    port map (
            O => \N__45245\,
            I => \N__45239\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__45242\,
            I => \sDAC_mem_27_1_sqmuxa\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__45239\,
            I => \sDAC_mem_27_1_sqmuxa\
        );

    \I__9981\ : InMux
    port map (
            O => \N__45234\,
            I => \N__45231\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__45231\,
            I => \N__45228\
        );

    \I__9979\ : Odrv12
    port map (
            O => \N__45228\,
            I => \sDAC_mem_13Z0Z_6\
        );

    \I__9978\ : InMux
    port map (
            O => \N__45225\,
            I => \N__45222\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__45222\,
            I => \sDAC_mem_13Z0Z_5\
        );

    \I__9976\ : InMux
    port map (
            O => \N__45219\,
            I => \N__45216\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__45216\,
            I => \N__45213\
        );

    \I__9974\ : Span4Mux_h
    port map (
            O => \N__45213\,
            I => \N__45210\
        );

    \I__9973\ : Odrv4
    port map (
            O => \N__45210\,
            I => \sDAC_mem_16Z0Z_1\
        );

    \I__9972\ : InMux
    port map (
            O => \N__45207\,
            I => \N__45204\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__45204\,
            I => \N__45201\
        );

    \I__9970\ : Span4Mux_v
    port map (
            O => \N__45201\,
            I => \N__45198\
        );

    \I__9969\ : Span4Mux_h
    port map (
            O => \N__45198\,
            I => \N__45195\
        );

    \I__9968\ : Odrv4
    port map (
            O => \N__45195\,
            I => \sDAC_mem_11Z0Z_2\
        );

    \I__9967\ : InMux
    port map (
            O => \N__45192\,
            I => \N__45189\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__45189\,
            I => \N__45186\
        );

    \I__9965\ : Span4Mux_v
    port map (
            O => \N__45186\,
            I => \N__45183\
        );

    \I__9964\ : Odrv4
    port map (
            O => \N__45183\,
            I => \sDAC_mem_11Z0Z_3\
        );

    \I__9963\ : InMux
    port map (
            O => \N__45180\,
            I => \N__45177\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__45177\,
            I => \N__45174\
        );

    \I__9961\ : Span4Mux_h
    port map (
            O => \N__45174\,
            I => \N__45171\
        );

    \I__9960\ : Span4Mux_v
    port map (
            O => \N__45171\,
            I => \N__45168\
        );

    \I__9959\ : Odrv4
    port map (
            O => \N__45168\,
            I => \sDAC_mem_11Z0Z_4\
        );

    \I__9958\ : InMux
    port map (
            O => \N__45165\,
            I => \N__45162\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__45162\,
            I => \N__45159\
        );

    \I__9956\ : Odrv4
    port map (
            O => \N__45159\,
            I => \sDAC_mem_11Z0Z_5\
        );

    \I__9955\ : InMux
    port map (
            O => \N__45156\,
            I => \N__45153\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__45153\,
            I => \N__45150\
        );

    \I__9953\ : Span4Mux_h
    port map (
            O => \N__45150\,
            I => \N__45147\
        );

    \I__9952\ : Span4Mux_v
    port map (
            O => \N__45147\,
            I => \N__45144\
        );

    \I__9951\ : Odrv4
    port map (
            O => \N__45144\,
            I => \sDAC_mem_11Z0Z_6\
        );

    \I__9950\ : InMux
    port map (
            O => \N__45141\,
            I => \N__45138\
        );

    \I__9949\ : LocalMux
    port map (
            O => \N__45138\,
            I => \N__45135\
        );

    \I__9948\ : Span4Mux_v
    port map (
            O => \N__45135\,
            I => \N__45132\
        );

    \I__9947\ : Odrv4
    port map (
            O => \N__45132\,
            I => \sDAC_mem_11Z0Z_7\
        );

    \I__9946\ : CEMux
    port map (
            O => \N__45129\,
            I => \N__45126\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__45126\,
            I => \sDAC_mem_11_1_sqmuxa\
        );

    \I__9944\ : InMux
    port map (
            O => \N__45123\,
            I => \N__45120\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__45120\,
            I => \N__45117\
        );

    \I__9942\ : Odrv12
    port map (
            O => \N__45117\,
            I => \sDAC_mem_15Z0Z_0\
        );

    \I__9941\ : InMux
    port map (
            O => \N__45114\,
            I => \N__45111\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__45111\,
            I => \sDAC_mem_14Z0Z_0\
        );

    \I__9939\ : CascadeMux
    port map (
            O => \N__45108\,
            I => \sDAC_data_RNO_18Z0Z_3_cascade_\
        );

    \I__9938\ : InMux
    port map (
            O => \N__45105\,
            I => \N__45102\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__45102\,
            I => \sDAC_data_RNO_19Z0Z_3\
        );

    \I__9936\ : InMux
    port map (
            O => \N__45099\,
            I => \N__45096\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__45096\,
            I => \N__45093\
        );

    \I__9934\ : Odrv4
    port map (
            O => \N__45093\,
            I => \sDAC_data_2_24_ns_1_3\
        );

    \I__9933\ : InMux
    port map (
            O => \N__45090\,
            I => \N__45087\
        );

    \I__9932\ : LocalMux
    port map (
            O => \N__45087\,
            I => \N__45084\
        );

    \I__9931\ : Span4Mux_v
    port map (
            O => \N__45084\,
            I => \N__45081\
        );

    \I__9930\ : Span4Mux_h
    port map (
            O => \N__45081\,
            I => \N__45078\
        );

    \I__9929\ : Odrv4
    port map (
            O => \N__45078\,
            I => \sDAC_mem_15Z0Z_2\
        );

    \I__9928\ : InMux
    port map (
            O => \N__45075\,
            I => \N__45072\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__45072\,
            I => \N__45069\
        );

    \I__9926\ : Span4Mux_v
    port map (
            O => \N__45069\,
            I => \N__45066\
        );

    \I__9925\ : Span4Mux_h
    port map (
            O => \N__45066\,
            I => \N__45063\
        );

    \I__9924\ : Odrv4
    port map (
            O => \N__45063\,
            I => \sDAC_mem_15Z0Z_3\
        );

    \I__9923\ : InMux
    port map (
            O => \N__45060\,
            I => \N__45057\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__45057\,
            I => \N__45054\
        );

    \I__9921\ : Span4Mux_v
    port map (
            O => \N__45054\,
            I => \N__45051\
        );

    \I__9920\ : Odrv4
    port map (
            O => \N__45051\,
            I => \sDAC_mem_15Z0Z_4\
        );

    \I__9919\ : InMux
    port map (
            O => \N__45048\,
            I => \N__45045\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__45045\,
            I => \N__45042\
        );

    \I__9917\ : Span4Mux_v
    port map (
            O => \N__45042\,
            I => \N__45039\
        );

    \I__9916\ : Odrv4
    port map (
            O => \N__45039\,
            I => \sDAC_mem_15Z0Z_5\
        );

    \I__9915\ : InMux
    port map (
            O => \N__45036\,
            I => \N__45033\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__45033\,
            I => \N__45030\
        );

    \I__9913\ : Span4Mux_v
    port map (
            O => \N__45030\,
            I => \N__45027\
        );

    \I__9912\ : Odrv4
    port map (
            O => \N__45027\,
            I => \sDAC_mem_15Z0Z_6\
        );

    \I__9911\ : CEMux
    port map (
            O => \N__45024\,
            I => \N__45021\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__45021\,
            I => \N__45018\
        );

    \I__9909\ : Span4Mux_h
    port map (
            O => \N__45018\,
            I => \N__45015\
        );

    \I__9908\ : Odrv4
    port map (
            O => \N__45015\,
            I => \sDAC_mem_15_1_sqmuxa\
        );

    \I__9907\ : InMux
    port map (
            O => \N__45012\,
            I => \N__45009\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__45009\,
            I => \sDAC_mem_11Z0Z_0\
        );

    \I__9905\ : InMux
    port map (
            O => \N__45006\,
            I => \N__45003\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__45003\,
            I => \sDAC_mem_11Z0Z_1\
        );

    \I__9903\ : CEMux
    port map (
            O => \N__45000\,
            I => \N__44997\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__44997\,
            I => \N__44994\
        );

    \I__9901\ : Span4Mux_h
    port map (
            O => \N__44994\,
            I => \N__44990\
        );

    \I__9900\ : CEMux
    port map (
            O => \N__44993\,
            I => \N__44987\
        );

    \I__9899\ : Span4Mux_h
    port map (
            O => \N__44990\,
            I => \N__44984\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__44987\,
            I => \N__44981\
        );

    \I__9897\ : Odrv4
    port map (
            O => \N__44984\,
            I => \sDAC_mem_10_1_sqmuxa\
        );

    \I__9896\ : Odrv12
    port map (
            O => \N__44981\,
            I => \sDAC_mem_10_1_sqmuxa\
        );

    \I__9895\ : CEMux
    port map (
            O => \N__44976\,
            I => \N__44973\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__44973\,
            I => \N__44970\
        );

    \I__9893\ : Span4Mux_v
    port map (
            O => \N__44970\,
            I => \N__44967\
        );

    \I__9892\ : Span4Mux_h
    port map (
            O => \N__44967\,
            I => \N__44964\
        );

    \I__9891\ : Odrv4
    port map (
            O => \N__44964\,
            I => \sDAC_mem_42_1_sqmuxa\
        );

    \I__9890\ : CascadeMux
    port map (
            O => \N__44961\,
            I => \N__44954\
        );

    \I__9889\ : InMux
    port map (
            O => \N__44960\,
            I => \N__44949\
        );

    \I__9888\ : InMux
    port map (
            O => \N__44959\,
            I => \N__44946\
        );

    \I__9887\ : InMux
    port map (
            O => \N__44958\,
            I => \N__44943\
        );

    \I__9886\ : InMux
    port map (
            O => \N__44957\,
            I => \N__44940\
        );

    \I__9885\ : InMux
    port map (
            O => \N__44954\,
            I => \N__44935\
        );

    \I__9884\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44935\
        );

    \I__9883\ : InMux
    port map (
            O => \N__44952\,
            I => \N__44932\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__44949\,
            I => \N__44926\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__44946\,
            I => \N__44926\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__44943\,
            I => \N__44923\
        );

    \I__9879\ : LocalMux
    port map (
            O => \N__44940\,
            I => \N__44920\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__44935\,
            I => \N__44915\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__44932\,
            I => \N__44915\
        );

    \I__9876\ : InMux
    port map (
            O => \N__44931\,
            I => \N__44912\
        );

    \I__9875\ : Span4Mux_h
    port map (
            O => \N__44926\,
            I => \N__44909\
        );

    \I__9874\ : Span4Mux_h
    port map (
            O => \N__44923\,
            I => \N__44906\
        );

    \I__9873\ : Span4Mux_v
    port map (
            O => \N__44920\,
            I => \N__44901\
        );

    \I__9872\ : Span4Mux_h
    port map (
            O => \N__44915\,
            I => \N__44901\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__44912\,
            I => \N__44898\
        );

    \I__9870\ : Span4Mux_h
    port map (
            O => \N__44909\,
            I => \N__44893\
        );

    \I__9869\ : Span4Mux_h
    port map (
            O => \N__44906\,
            I => \N__44890\
        );

    \I__9868\ : Span4Mux_h
    port map (
            O => \N__44901\,
            I => \N__44885\
        );

    \I__9867\ : Span4Mux_h
    port map (
            O => \N__44898\,
            I => \N__44885\
        );

    \I__9866\ : InMux
    port map (
            O => \N__44897\,
            I => \N__44880\
        );

    \I__9865\ : InMux
    port map (
            O => \N__44896\,
            I => \N__44880\
        );

    \I__9864\ : Odrv4
    port map (
            O => \N__44893\,
            I => \sAddressZ0Z_2\
        );

    \I__9863\ : Odrv4
    port map (
            O => \N__44890\,
            I => \sAddressZ0Z_2\
        );

    \I__9862\ : Odrv4
    port map (
            O => \N__44885\,
            I => \sAddressZ0Z_2\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__44880\,
            I => \sAddressZ0Z_2\
        );

    \I__9860\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44865\
        );

    \I__9859\ : InMux
    port map (
            O => \N__44870\,
            I => \N__44862\
        );

    \I__9858\ : InMux
    port map (
            O => \N__44869\,
            I => \N__44859\
        );

    \I__9857\ : InMux
    port map (
            O => \N__44868\,
            I => \N__44856\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__44865\,
            I => \N__44848\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__44862\,
            I => \N__44848\
        );

    \I__9854\ : LocalMux
    port map (
            O => \N__44859\,
            I => \N__44848\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__44856\,
            I => \N__44845\
        );

    \I__9852\ : InMux
    port map (
            O => \N__44855\,
            I => \N__44842\
        );

    \I__9851\ : Span4Mux_v
    port map (
            O => \N__44848\,
            I => \N__44839\
        );

    \I__9850\ : Span4Mux_h
    port map (
            O => \N__44845\,
            I => \N__44836\
        );

    \I__9849\ : LocalMux
    port map (
            O => \N__44842\,
            I => \N__44833\
        );

    \I__9848\ : Span4Mux_h
    port map (
            O => \N__44839\,
            I => \N__44828\
        );

    \I__9847\ : Span4Mux_h
    port map (
            O => \N__44836\,
            I => \N__44825\
        );

    \I__9846\ : Span4Mux_v
    port map (
            O => \N__44833\,
            I => \N__44822\
        );

    \I__9845\ : InMux
    port map (
            O => \N__44832\,
            I => \N__44817\
        );

    \I__9844\ : InMux
    port map (
            O => \N__44831\,
            I => \N__44817\
        );

    \I__9843\ : Odrv4
    port map (
            O => \N__44828\,
            I => \sAddressZ0Z_1\
        );

    \I__9842\ : Odrv4
    port map (
            O => \N__44825\,
            I => \sAddressZ0Z_1\
        );

    \I__9841\ : Odrv4
    port map (
            O => \N__44822\,
            I => \sAddressZ0Z_1\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__44817\,
            I => \sAddressZ0Z_1\
        );

    \I__9839\ : CascadeMux
    port map (
            O => \N__44808\,
            I => \N__44804\
        );

    \I__9838\ : CascadeMux
    port map (
            O => \N__44807\,
            I => \N__44801\
        );

    \I__9837\ : InMux
    port map (
            O => \N__44804\,
            I => \N__44798\
        );

    \I__9836\ : InMux
    port map (
            O => \N__44801\,
            I => \N__44794\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__44798\,
            I => \N__44791\
        );

    \I__9834\ : CascadeMux
    port map (
            O => \N__44797\,
            I => \N__44788\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__44794\,
            I => \N__44785\
        );

    \I__9832\ : Span4Mux_h
    port map (
            O => \N__44791\,
            I => \N__44782\
        );

    \I__9831\ : InMux
    port map (
            O => \N__44788\,
            I => \N__44779\
        );

    \I__9830\ : Span4Mux_v
    port map (
            O => \N__44785\,
            I => \N__44775\
        );

    \I__9829\ : Span4Mux_v
    port map (
            O => \N__44782\,
            I => \N__44770\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__44779\,
            I => \N__44770\
        );

    \I__9827\ : InMux
    port map (
            O => \N__44778\,
            I => \N__44767\
        );

    \I__9826\ : Span4Mux_v
    port map (
            O => \N__44775\,
            I => \N__44762\
        );

    \I__9825\ : Span4Mux_v
    port map (
            O => \N__44770\,
            I => \N__44762\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__44767\,
            I => \N__44759\
        );

    \I__9823\ : Sp12to4
    port map (
            O => \N__44762\,
            I => \N__44754\
        );

    \I__9822\ : Sp12to4
    port map (
            O => \N__44759\,
            I => \N__44754\
        );

    \I__9821\ : Odrv12
    port map (
            O => \N__44754\,
            I => \sDAC_mem_30_1_sqmuxa_0_a2_1_0\
        );

    \I__9820\ : InMux
    port map (
            O => \N__44751\,
            I => \N__44746\
        );

    \I__9819\ : InMux
    port map (
            O => \N__44750\,
            I => \N__44742\
        );

    \I__9818\ : InMux
    port map (
            O => \N__44749\,
            I => \N__44738\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__44746\,
            I => \N__44735\
        );

    \I__9816\ : InMux
    port map (
            O => \N__44745\,
            I => \N__44732\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__44742\,
            I => \N__44727\
        );

    \I__9814\ : InMux
    port map (
            O => \N__44741\,
            I => \N__44724\
        );

    \I__9813\ : LocalMux
    port map (
            O => \N__44738\,
            I => \N__44719\
        );

    \I__9812\ : Span4Mux_v
    port map (
            O => \N__44735\,
            I => \N__44711\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__44732\,
            I => \N__44711\
        );

    \I__9810\ : InMux
    port map (
            O => \N__44731\,
            I => \N__44706\
        );

    \I__9809\ : InMux
    port map (
            O => \N__44730\,
            I => \N__44706\
        );

    \I__9808\ : Span4Mux_v
    port map (
            O => \N__44727\,
            I => \N__44701\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__44724\,
            I => \N__44701\
        );

    \I__9806\ : InMux
    port map (
            O => \N__44723\,
            I => \N__44698\
        );

    \I__9805\ : InMux
    port map (
            O => \N__44722\,
            I => \N__44695\
        );

    \I__9804\ : Span4Mux_h
    port map (
            O => \N__44719\,
            I => \N__44690\
        );

    \I__9803\ : InMux
    port map (
            O => \N__44718\,
            I => \N__44687\
        );

    \I__9802\ : InMux
    port map (
            O => \N__44717\,
            I => \N__44682\
        );

    \I__9801\ : InMux
    port map (
            O => \N__44716\,
            I => \N__44682\
        );

    \I__9800\ : Span4Mux_h
    port map (
            O => \N__44711\,
            I => \N__44679\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__44706\,
            I => \N__44674\
        );

    \I__9798\ : Span4Mux_h
    port map (
            O => \N__44701\,
            I => \N__44674\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__44698\,
            I => \N__44669\
        );

    \I__9796\ : LocalMux
    port map (
            O => \N__44695\,
            I => \N__44669\
        );

    \I__9795\ : InMux
    port map (
            O => \N__44694\,
            I => \N__44664\
        );

    \I__9794\ : InMux
    port map (
            O => \N__44693\,
            I => \N__44664\
        );

    \I__9793\ : Odrv4
    port map (
            O => \N__44690\,
            I => \N_275\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__44687\,
            I => \N_275\
        );

    \I__9791\ : LocalMux
    port map (
            O => \N__44682\,
            I => \N_275\
        );

    \I__9790\ : Odrv4
    port map (
            O => \N__44679\,
            I => \N_275\
        );

    \I__9789\ : Odrv4
    port map (
            O => \N__44674\,
            I => \N_275\
        );

    \I__9788\ : Odrv12
    port map (
            O => \N__44669\,
            I => \N_275\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__44664\,
            I => \N_275\
        );

    \I__9786\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44646\
        );

    \I__9785\ : LocalMux
    port map (
            O => \N__44646\,
            I => \N__44641\
        );

    \I__9784\ : InMux
    port map (
            O => \N__44645\,
            I => \N__44638\
        );

    \I__9783\ : InMux
    port map (
            O => \N__44644\,
            I => \N__44633\
        );

    \I__9782\ : Span4Mux_v
    port map (
            O => \N__44641\,
            I => \N__44628\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__44638\,
            I => \N__44628\
        );

    \I__9780\ : InMux
    port map (
            O => \N__44637\,
            I => \N__44625\
        );

    \I__9779\ : InMux
    port map (
            O => \N__44636\,
            I => \N__44622\
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__44633\,
            I => \N__44617\
        );

    \I__9777\ : Span4Mux_h
    port map (
            O => \N__44628\,
            I => \N__44617\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__44625\,
            I => \N__44614\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__44622\,
            I => \N__44610\
        );

    \I__9774\ : Span4Mux_v
    port map (
            O => \N__44617\,
            I => \N__44605\
        );

    \I__9773\ : Span4Mux_v
    port map (
            O => \N__44614\,
            I => \N__44605\
        );

    \I__9772\ : InMux
    port map (
            O => \N__44613\,
            I => \N__44602\
        );

    \I__9771\ : Odrv12
    port map (
            O => \N__44610\,
            I => \sAddressZ0Z_4\
        );

    \I__9770\ : Odrv4
    port map (
            O => \N__44605\,
            I => \sAddressZ0Z_4\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__44602\,
            I => \sAddressZ0Z_4\
        );

    \I__9768\ : CascadeMux
    port map (
            O => \N__44595\,
            I => \N__44589\
        );

    \I__9767\ : CascadeMux
    port map (
            O => \N__44594\,
            I => \N__44583\
        );

    \I__9766\ : CascadeMux
    port map (
            O => \N__44593\,
            I => \N__44580\
        );

    \I__9765\ : InMux
    port map (
            O => \N__44592\,
            I => \N__44577\
        );

    \I__9764\ : InMux
    port map (
            O => \N__44589\,
            I => \N__44572\
        );

    \I__9763\ : InMux
    port map (
            O => \N__44588\,
            I => \N__44572\
        );

    \I__9762\ : CascadeMux
    port map (
            O => \N__44587\,
            I => \N__44568\
        );

    \I__9761\ : CascadeMux
    port map (
            O => \N__44586\,
            I => \N__44565\
        );

    \I__9760\ : InMux
    port map (
            O => \N__44583\,
            I => \N__44560\
        );

    \I__9759\ : InMux
    port map (
            O => \N__44580\,
            I => \N__44560\
        );

    \I__9758\ : LocalMux
    port map (
            O => \N__44577\,
            I => \N__44555\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__44572\,
            I => \N__44555\
        );

    \I__9756\ : CascadeMux
    port map (
            O => \N__44571\,
            I => \N__44550\
        );

    \I__9755\ : InMux
    port map (
            O => \N__44568\,
            I => \N__44546\
        );

    \I__9754\ : InMux
    port map (
            O => \N__44565\,
            I => \N__44543\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__44560\,
            I => \N__44540\
        );

    \I__9752\ : Span4Mux_h
    port map (
            O => \N__44555\,
            I => \N__44536\
        );

    \I__9751\ : CascadeMux
    port map (
            O => \N__44554\,
            I => \N__44533\
        );

    \I__9750\ : InMux
    port map (
            O => \N__44553\,
            I => \N__44528\
        );

    \I__9749\ : InMux
    port map (
            O => \N__44550\,
            I => \N__44528\
        );

    \I__9748\ : InMux
    port map (
            O => \N__44549\,
            I => \N__44525\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__44546\,
            I => \N__44520\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__44543\,
            I => \N__44520\
        );

    \I__9745\ : Span4Mux_h
    port map (
            O => \N__44540\,
            I => \N__44517\
        );

    \I__9744\ : InMux
    port map (
            O => \N__44539\,
            I => \N__44514\
        );

    \I__9743\ : Span4Mux_h
    port map (
            O => \N__44536\,
            I => \N__44511\
        );

    \I__9742\ : InMux
    port map (
            O => \N__44533\,
            I => \N__44508\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__44528\,
            I => \N__44503\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__44525\,
            I => \N__44503\
        );

    \I__9739\ : Span4Mux_h
    port map (
            O => \N__44520\,
            I => \N__44500\
        );

    \I__9738\ : Span4Mux_v
    port map (
            O => \N__44517\,
            I => \N__44497\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__44514\,
            I => \N__44492\
        );

    \I__9736\ : Span4Mux_h
    port map (
            O => \N__44511\,
            I => \N__44492\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__44508\,
            I => \N_286\
        );

    \I__9734\ : Odrv12
    port map (
            O => \N__44503\,
            I => \N_286\
        );

    \I__9733\ : Odrv4
    port map (
            O => \N__44500\,
            I => \N_286\
        );

    \I__9732\ : Odrv4
    port map (
            O => \N__44497\,
            I => \N_286\
        );

    \I__9731\ : Odrv4
    port map (
            O => \N__44492\,
            I => \N_286\
        );

    \I__9730\ : CascadeMux
    port map (
            O => \N__44481\,
            I => \N_278_cascade_\
        );

    \I__9729\ : CascadeMux
    port map (
            O => \N__44478\,
            I => \N__44475\
        );

    \I__9728\ : InMux
    port map (
            O => \N__44475\,
            I => \N__44472\
        );

    \I__9727\ : LocalMux
    port map (
            O => \N__44472\,
            I => \N__44466\
        );

    \I__9726\ : CascadeMux
    port map (
            O => \N__44471\,
            I => \N__44463\
        );

    \I__9725\ : CascadeMux
    port map (
            O => \N__44470\,
            I => \N__44460\
        );

    \I__9724\ : CascadeMux
    port map (
            O => \N__44469\,
            I => \N__44456\
        );

    \I__9723\ : Span4Mux_h
    port map (
            O => \N__44466\,
            I => \N__44453\
        );

    \I__9722\ : InMux
    port map (
            O => \N__44463\,
            I => \N__44446\
        );

    \I__9721\ : InMux
    port map (
            O => \N__44460\,
            I => \N__44446\
        );

    \I__9720\ : InMux
    port map (
            O => \N__44459\,
            I => \N__44446\
        );

    \I__9719\ : InMux
    port map (
            O => \N__44456\,
            I => \N__44440\
        );

    \I__9718\ : Span4Mux_v
    port map (
            O => \N__44453\,
            I => \N__44437\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__44446\,
            I => \N__44434\
        );

    \I__9716\ : InMux
    port map (
            O => \N__44445\,
            I => \N__44431\
        );

    \I__9715\ : InMux
    port map (
            O => \N__44444\,
            I => \N__44425\
        );

    \I__9714\ : InMux
    port map (
            O => \N__44443\,
            I => \N__44425\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__44440\,
            I => \N__44422\
        );

    \I__9712\ : Span4Mux_h
    port map (
            O => \N__44437\,
            I => \N__44415\
        );

    \I__9711\ : Span4Mux_v
    port map (
            O => \N__44434\,
            I => \N__44415\
        );

    \I__9710\ : LocalMux
    port map (
            O => \N__44431\,
            I => \N__44415\
        );

    \I__9709\ : InMux
    port map (
            O => \N__44430\,
            I => \N__44412\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__44425\,
            I => \N__44406\
        );

    \I__9707\ : Span12Mux_v
    port map (
            O => \N__44422\,
            I => \N__44403\
        );

    \I__9706\ : Span4Mux_h
    port map (
            O => \N__44415\,
            I => \N__44400\
        );

    \I__9705\ : LocalMux
    port map (
            O => \N__44412\,
            I => \N__44397\
        );

    \I__9704\ : InMux
    port map (
            O => \N__44411\,
            I => \N__44390\
        );

    \I__9703\ : InMux
    port map (
            O => \N__44410\,
            I => \N__44390\
        );

    \I__9702\ : InMux
    port map (
            O => \N__44409\,
            I => \N__44390\
        );

    \I__9701\ : Span4Mux_h
    port map (
            O => \N__44406\,
            I => \N__44387\
        );

    \I__9700\ : Odrv12
    port map (
            O => \N__44403\,
            I => \N_142\
        );

    \I__9699\ : Odrv4
    port map (
            O => \N__44400\,
            I => \N_142\
        );

    \I__9698\ : Odrv4
    port map (
            O => \N__44397\,
            I => \N_142\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__44390\,
            I => \N_142\
        );

    \I__9696\ : Odrv4
    port map (
            O => \N__44387\,
            I => \N_142\
        );

    \I__9695\ : InMux
    port map (
            O => \N__44376\,
            I => \N__44373\
        );

    \I__9694\ : LocalMux
    port map (
            O => \N__44373\,
            I => \N__44370\
        );

    \I__9693\ : Odrv4
    port map (
            O => \N__44370\,
            I => \sDAC_mem_42Z0Z_5\
        );

    \I__9692\ : InMux
    port map (
            O => \N__44367\,
            I => \N__44364\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__44364\,
            I => \N__44361\
        );

    \I__9690\ : Span4Mux_h
    port map (
            O => \N__44361\,
            I => \N__44358\
        );

    \I__9689\ : Odrv4
    port map (
            O => \N__44358\,
            I => \sDAC_mem_42Z0Z_6\
        );

    \I__9688\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44352\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__44352\,
            I => \N__44349\
        );

    \I__9686\ : Span4Mux_h
    port map (
            O => \N__44349\,
            I => \N__44346\
        );

    \I__9685\ : Span4Mux_h
    port map (
            O => \N__44346\,
            I => \N__44343\
        );

    \I__9684\ : Odrv4
    port map (
            O => \N__44343\,
            I => \sDAC_mem_42Z0Z_7\
        );

    \I__9683\ : InMux
    port map (
            O => \N__44340\,
            I => \N__44337\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__44337\,
            I => \N__44334\
        );

    \I__9681\ : Odrv4
    port map (
            O => \N__44334\,
            I => \sDAC_mem_10Z0Z_0\
        );

    \I__9680\ : InMux
    port map (
            O => \N__44331\,
            I => \N__44328\
        );

    \I__9679\ : LocalMux
    port map (
            O => \N__44328\,
            I => \N__44325\
        );

    \I__9678\ : Span4Mux_v
    port map (
            O => \N__44325\,
            I => \N__44322\
        );

    \I__9677\ : Odrv4
    port map (
            O => \N__44322\,
            I => \sDAC_mem_10Z0Z_1\
        );

    \I__9676\ : InMux
    port map (
            O => \N__44319\,
            I => \N__44316\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__44316\,
            I => \N__44313\
        );

    \I__9674\ : Span4Mux_h
    port map (
            O => \N__44313\,
            I => \N__44310\
        );

    \I__9673\ : Span4Mux_h
    port map (
            O => \N__44310\,
            I => \N__44307\
        );

    \I__9672\ : Odrv4
    port map (
            O => \N__44307\,
            I => \sDAC_mem_10Z0Z_2\
        );

    \I__9671\ : InMux
    port map (
            O => \N__44304\,
            I => \N__44301\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__44301\,
            I => \N__44298\
        );

    \I__9669\ : Span4Mux_h
    port map (
            O => \N__44298\,
            I => \N__44295\
        );

    \I__9668\ : Odrv4
    port map (
            O => \N__44295\,
            I => \sDAC_mem_10Z0Z_3\
        );

    \I__9667\ : InMux
    port map (
            O => \N__44292\,
            I => \N__44289\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__44289\,
            I => \N__44286\
        );

    \I__9665\ : Span4Mux_h
    port map (
            O => \N__44286\,
            I => \N__44283\
        );

    \I__9664\ : Span4Mux_h
    port map (
            O => \N__44283\,
            I => \N__44280\
        );

    \I__9663\ : Odrv4
    port map (
            O => \N__44280\,
            I => \sDAC_mem_10Z0Z_4\
        );

    \I__9662\ : InMux
    port map (
            O => \N__44277\,
            I => \N__44274\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__44274\,
            I => \sDAC_mem_10Z0Z_5\
        );

    \I__9660\ : InMux
    port map (
            O => \N__44271\,
            I => \N__44268\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__44268\,
            I => \N__44265\
        );

    \I__9658\ : Span4Mux_h
    port map (
            O => \N__44265\,
            I => \N__44262\
        );

    \I__9657\ : Odrv4
    port map (
            O => \N__44262\,
            I => \sDAC_mem_10Z0Z_6\
        );

    \I__9656\ : InMux
    port map (
            O => \N__44259\,
            I => \N__44256\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__44256\,
            I => \N__44253\
        );

    \I__9654\ : Span4Mux_v
    port map (
            O => \N__44253\,
            I => \N__44250\
        );

    \I__9653\ : Span4Mux_h
    port map (
            O => \N__44250\,
            I => \N__44247\
        );

    \I__9652\ : Odrv4
    port map (
            O => \N__44247\,
            I => \sDAC_mem_41Z0Z_4\
        );

    \I__9651\ : InMux
    port map (
            O => \N__44244\,
            I => \N__44241\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__44241\,
            I => \N__44238\
        );

    \I__9649\ : Span4Mux_h
    port map (
            O => \N__44238\,
            I => \N__44235\
        );

    \I__9648\ : Odrv4
    port map (
            O => \N__44235\,
            I => \sDAC_mem_41Z0Z_5\
        );

    \I__9647\ : InMux
    port map (
            O => \N__44232\,
            I => \N__44229\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__44229\,
            I => \N__44226\
        );

    \I__9645\ : Span4Mux_h
    port map (
            O => \N__44226\,
            I => \N__44223\
        );

    \I__9644\ : Odrv4
    port map (
            O => \N__44223\,
            I => \sDAC_mem_41Z0Z_6\
        );

    \I__9643\ : InMux
    port map (
            O => \N__44220\,
            I => \N__44217\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__44217\,
            I => \N__44214\
        );

    \I__9641\ : Span4Mux_v
    port map (
            O => \N__44214\,
            I => \N__44211\
        );

    \I__9640\ : Odrv4
    port map (
            O => \N__44211\,
            I => \sDAC_mem_41Z0Z_7\
        );

    \I__9639\ : InMux
    port map (
            O => \N__44208\,
            I => \N__44205\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__44205\,
            I => \N__44202\
        );

    \I__9637\ : Span4Mux_v
    port map (
            O => \N__44202\,
            I => \N__44199\
        );

    \I__9636\ : Odrv4
    port map (
            O => \N__44199\,
            I => \sDAC_mem_42Z0Z_0\
        );

    \I__9635\ : InMux
    port map (
            O => \N__44196\,
            I => \N__44193\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__44193\,
            I => \N__44190\
        );

    \I__9633\ : Span4Mux_v
    port map (
            O => \N__44190\,
            I => \N__44187\
        );

    \I__9632\ : Odrv4
    port map (
            O => \N__44187\,
            I => \sDAC_mem_42Z0Z_1\
        );

    \I__9631\ : InMux
    port map (
            O => \N__44184\,
            I => \N__44181\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__44181\,
            I => \N__44178\
        );

    \I__9629\ : Span12Mux_h
    port map (
            O => \N__44178\,
            I => \N__44175\
        );

    \I__9628\ : Odrv12
    port map (
            O => \N__44175\,
            I => \sDAC_mem_42Z0Z_2\
        );

    \I__9627\ : InMux
    port map (
            O => \N__44172\,
            I => \N__44169\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__44169\,
            I => \N__44166\
        );

    \I__9625\ : Span4Mux_v
    port map (
            O => \N__44166\,
            I => \N__44163\
        );

    \I__9624\ : Span4Mux_h
    port map (
            O => \N__44163\,
            I => \N__44160\
        );

    \I__9623\ : Odrv4
    port map (
            O => \N__44160\,
            I => \sDAC_mem_42Z0Z_3\
        );

    \I__9622\ : InMux
    port map (
            O => \N__44157\,
            I => \N__44154\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__44154\,
            I => \N__44151\
        );

    \I__9620\ : Odrv12
    port map (
            O => \N__44151\,
            I => \sDAC_mem_42Z0Z_4\
        );

    \I__9619\ : InMux
    port map (
            O => \N__44148\,
            I => \N__44145\
        );

    \I__9618\ : LocalMux
    port map (
            O => \N__44145\,
            I => \sDAC_mem_12Z0Z_5\
        );

    \I__9617\ : CascadeMux
    port map (
            O => \N__44142\,
            I => \N__44139\
        );

    \I__9616\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44136\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__44136\,
            I => \N__44133\
        );

    \I__9614\ : Span4Mux_h
    port map (
            O => \N__44133\,
            I => \N__44130\
        );

    \I__9613\ : Odrv4
    port map (
            O => \N__44130\,
            I => \sEEADC_freqZ0Z_1\
        );

    \I__9612\ : CEMux
    port map (
            O => \N__44127\,
            I => \N__44123\
        );

    \I__9611\ : CEMux
    port map (
            O => \N__44126\,
            I => \N__44119\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__44123\,
            I => \N__44116\
        );

    \I__9609\ : CEMux
    port map (
            O => \N__44122\,
            I => \N__44113\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__44119\,
            I => \N__44110\
        );

    \I__9607\ : Span4Mux_h
    port map (
            O => \N__44116\,
            I => \N__44105\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__44113\,
            I => \N__44105\
        );

    \I__9605\ : Span4Mux_h
    port map (
            O => \N__44110\,
            I => \N__44102\
        );

    \I__9604\ : Span4Mux_h
    port map (
            O => \N__44105\,
            I => \N__44099\
        );

    \I__9603\ : Odrv4
    port map (
            O => \N__44102\,
            I => \sEEADC_freq_1_sqmuxa\
        );

    \I__9602\ : Odrv4
    port map (
            O => \N__44099\,
            I => \sEEADC_freq_1_sqmuxa\
        );

    \I__9601\ : InMux
    port map (
            O => \N__44094\,
            I => \N__44091\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__44091\,
            I => \N__44088\
        );

    \I__9599\ : Span12Mux_h
    port map (
            O => \N__44088\,
            I => \N__44085\
        );

    \I__9598\ : Odrv12
    port map (
            O => \N__44085\,
            I => \sDAC_mem_17Z0Z_0\
        );

    \I__9597\ : InMux
    port map (
            O => \N__44082\,
            I => \N__44079\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__44079\,
            I => \N__44076\
        );

    \I__9595\ : Span4Mux_h
    port map (
            O => \N__44076\,
            I => \N__44073\
        );

    \I__9594\ : Odrv4
    port map (
            O => \N__44073\,
            I => \sDAC_mem_16Z0Z_0\
        );

    \I__9593\ : CascadeMux
    port map (
            O => \N__44070\,
            I => \N__44067\
        );

    \I__9592\ : InMux
    port map (
            O => \N__44067\,
            I => \N__44064\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__44064\,
            I => \N__44061\
        );

    \I__9590\ : Span4Mux_v
    port map (
            O => \N__44061\,
            I => \N__44058\
        );

    \I__9589\ : Odrv4
    port map (
            O => \N__44058\,
            I => \sDAC_data_RNO_29Z0Z_3\
        );

    \I__9588\ : InMux
    port map (
            O => \N__44055\,
            I => \N__44052\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__44052\,
            I => \N__44049\
        );

    \I__9586\ : Odrv12
    port map (
            O => \N__44049\,
            I => \sDAC_mem_16Z0Z_3\
        );

    \I__9585\ : InMux
    port map (
            O => \N__44046\,
            I => \N__44043\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__44043\,
            I => \N__44040\
        );

    \I__9583\ : Span4Mux_v
    port map (
            O => \N__44040\,
            I => \N__44037\
        );

    \I__9582\ : Span4Mux_v
    port map (
            O => \N__44037\,
            I => \N__44034\
        );

    \I__9581\ : Odrv4
    port map (
            O => \N__44034\,
            I => \sDAC_mem_20Z0Z_7\
        );

    \I__9580\ : CEMux
    port map (
            O => \N__44031\,
            I => \N__44026\
        );

    \I__9579\ : CEMux
    port map (
            O => \N__44030\,
            I => \N__44023\
        );

    \I__9578\ : CEMux
    port map (
            O => \N__44029\,
            I => \N__44020\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__44026\,
            I => \N__44017\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__44023\,
            I => \N__44014\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__44020\,
            I => \N__44011\
        );

    \I__9574\ : Span4Mux_h
    port map (
            O => \N__44017\,
            I => \N__44008\
        );

    \I__9573\ : Span4Mux_h
    port map (
            O => \N__44014\,
            I => \N__44003\
        );

    \I__9572\ : Span4Mux_h
    port map (
            O => \N__44011\,
            I => \N__44003\
        );

    \I__9571\ : Odrv4
    port map (
            O => \N__44008\,
            I => \sDAC_mem_20_1_sqmuxa\
        );

    \I__9570\ : Odrv4
    port map (
            O => \N__44003\,
            I => \sDAC_mem_20_1_sqmuxa\
        );

    \I__9569\ : InMux
    port map (
            O => \N__43998\,
            I => \N__43995\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__43995\,
            I => \N__43992\
        );

    \I__9567\ : Span4Mux_v
    port map (
            O => \N__43992\,
            I => \N__43989\
        );

    \I__9566\ : Odrv4
    port map (
            O => \N__43989\,
            I => \sDAC_mem_41Z0Z_0\
        );

    \I__9565\ : InMux
    port map (
            O => \N__43986\,
            I => \N__43983\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__43983\,
            I => \N__43980\
        );

    \I__9563\ : Span4Mux_v
    port map (
            O => \N__43980\,
            I => \N__43977\
        );

    \I__9562\ : Odrv4
    port map (
            O => \N__43977\,
            I => \sDAC_mem_41Z0Z_1\
        );

    \I__9561\ : InMux
    port map (
            O => \N__43974\,
            I => \N__43971\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__43971\,
            I => \N__43968\
        );

    \I__9559\ : Span4Mux_h
    port map (
            O => \N__43968\,
            I => \N__43965\
        );

    \I__9558\ : Span4Mux_h
    port map (
            O => \N__43965\,
            I => \N__43962\
        );

    \I__9557\ : Odrv4
    port map (
            O => \N__43962\,
            I => \sDAC_mem_41Z0Z_2\
        );

    \I__9556\ : InMux
    port map (
            O => \N__43959\,
            I => \N__43956\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__43956\,
            I => \N__43953\
        );

    \I__9554\ : Span4Mux_h
    port map (
            O => \N__43953\,
            I => \N__43950\
        );

    \I__9553\ : Odrv4
    port map (
            O => \N__43950\,
            I => \sDAC_mem_41Z0Z_3\
        );

    \I__9552\ : InMux
    port map (
            O => \N__43947\,
            I => \N__43944\
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__43944\,
            I => \N__43941\
        );

    \I__9550\ : Span4Mux_h
    port map (
            O => \N__43941\,
            I => \N__43938\
        );

    \I__9549\ : Odrv4
    port map (
            O => \N__43938\,
            I => \sDAC_mem_14Z0Z_6\
        );

    \I__9548\ : CEMux
    port map (
            O => \N__43935\,
            I => \N__43932\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__43932\,
            I => \sDAC_mem_14_1_sqmuxa\
        );

    \I__9546\ : InMux
    port map (
            O => \N__43929\,
            I => \N__43926\
        );

    \I__9545\ : LocalMux
    port map (
            O => \N__43926\,
            I => \sDAC_mem_14Z0Z_4\
        );

    \I__9544\ : CascadeMux
    port map (
            O => \N__43923\,
            I => \sDAC_data_RNO_18Z0Z_7_cascade_\
        );

    \I__9543\ : InMux
    port map (
            O => \N__43920\,
            I => \N__43917\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__43917\,
            I => \sDAC_data_RNO_19Z0Z_7\
        );

    \I__9541\ : InMux
    port map (
            O => \N__43914\,
            I => \N__43911\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__43911\,
            I => \N__43908\
        );

    \I__9539\ : Span4Mux_h
    port map (
            O => \N__43908\,
            I => \N__43905\
        );

    \I__9538\ : Span4Mux_v
    port map (
            O => \N__43905\,
            I => \N__43902\
        );

    \I__9537\ : Odrv4
    port map (
            O => \N__43902\,
            I => \sDAC_data_2_24_ns_1_7\
        );

    \I__9536\ : CascadeMux
    port map (
            O => \N__43899\,
            I => \sDAC_data_RNO_18Z0Z_8_cascade_\
        );

    \I__9535\ : InMux
    port map (
            O => \N__43896\,
            I => \N__43893\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__43893\,
            I => \N__43890\
        );

    \I__9533\ : Odrv12
    port map (
            O => \N__43890\,
            I => \sDAC_data_2_24_ns_1_8\
        );

    \I__9532\ : InMux
    port map (
            O => \N__43887\,
            I => \N__43884\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__43884\,
            I => \sDAC_mem_12Z0Z_4\
        );

    \I__9530\ : InMux
    port map (
            O => \N__43881\,
            I => \N__43878\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__43878\,
            I => \sDAC_mem_14Z0Z_5\
        );

    \I__9528\ : InMux
    port map (
            O => \N__43875\,
            I => \N__43872\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__43872\,
            I => \sDAC_data_RNO_19Z0Z_8\
        );

    \I__9526\ : InMux
    port map (
            O => \N__43869\,
            I => \N__43863\
        );

    \I__9525\ : InMux
    port map (
            O => \N__43868\,
            I => \N__43863\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__43863\,
            I => \N__43857\
        );

    \I__9523\ : InMux
    port map (
            O => \N__43862\,
            I => \N__43848\
        );

    \I__9522\ : InMux
    port map (
            O => \N__43861\,
            I => \N__43848\
        );

    \I__9521\ : InMux
    port map (
            O => \N__43860\,
            I => \N__43848\
        );

    \I__9520\ : Span4Mux_v
    port map (
            O => \N__43857\,
            I => \N__43840\
        );

    \I__9519\ : InMux
    port map (
            O => \N__43856\,
            I => \N__43837\
        );

    \I__9518\ : InMux
    port map (
            O => \N__43855\,
            I => \N__43834\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__43848\,
            I => \N__43829\
        );

    \I__9516\ : InMux
    port map (
            O => \N__43847\,
            I => \N__43824\
        );

    \I__9515\ : InMux
    port map (
            O => \N__43846\,
            I => \N__43824\
        );

    \I__9514\ : InMux
    port map (
            O => \N__43845\,
            I => \N__43817\
        );

    \I__9513\ : InMux
    port map (
            O => \N__43844\,
            I => \N__43817\
        );

    \I__9512\ : InMux
    port map (
            O => \N__43843\,
            I => \N__43817\
        );

    \I__9511\ : Span4Mux_h
    port map (
            O => \N__43840\,
            I => \N__43812\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__43837\,
            I => \N__43812\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__43834\,
            I => \N__43809\
        );

    \I__9508\ : InMux
    port map (
            O => \N__43833\,
            I => \N__43806\
        );

    \I__9507\ : InMux
    port map (
            O => \N__43832\,
            I => \N__43803\
        );

    \I__9506\ : Span4Mux_v
    port map (
            O => \N__43829\,
            I => \N__43800\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__43824\,
            I => \N__43797\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__43817\,
            I => \N__43792\
        );

    \I__9503\ : Span4Mux_h
    port map (
            O => \N__43812\,
            I => \N__43792\
        );

    \I__9502\ : Odrv12
    port map (
            O => \N__43809\,
            I => \sPointerZ0Z_1\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__43806\,
            I => \sPointerZ0Z_1\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__43803\,
            I => \sPointerZ0Z_1\
        );

    \I__9499\ : Odrv4
    port map (
            O => \N__43800\,
            I => \sPointerZ0Z_1\
        );

    \I__9498\ : Odrv12
    port map (
            O => \N__43797\,
            I => \sPointerZ0Z_1\
        );

    \I__9497\ : Odrv4
    port map (
            O => \N__43792\,
            I => \sPointerZ0Z_1\
        );

    \I__9496\ : CEMux
    port map (
            O => \N__43779\,
            I => \N__43776\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__43776\,
            I => \N__43772\
        );

    \I__9494\ : CEMux
    port map (
            O => \N__43775\,
            I => \N__43768\
        );

    \I__9493\ : Span4Mux_v
    port map (
            O => \N__43772\,
            I => \N__43765\
        );

    \I__9492\ : CEMux
    port map (
            O => \N__43771\,
            I => \N__43762\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__43768\,
            I => \N__43759\
        );

    \I__9490\ : Span4Mux_h
    port map (
            O => \N__43765\,
            I => \N__43754\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__43762\,
            I => \N__43754\
        );

    \I__9488\ : Span4Mux_v
    port map (
            O => \N__43759\,
            I => \N__43751\
        );

    \I__9487\ : Sp12to4
    port map (
            O => \N__43754\,
            I => \N__43748\
        );

    \I__9486\ : Span4Mux_h
    port map (
            O => \N__43751\,
            I => \N__43745\
        );

    \I__9485\ : Odrv12
    port map (
            O => \N__43748\,
            I => un1_spointer11_0
        );

    \I__9484\ : Odrv4
    port map (
            O => \N__43745\,
            I => un1_spointer11_0
        );

    \I__9483\ : InMux
    port map (
            O => \N__43740\,
            I => \N__43737\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__43737\,
            I => \N__43734\
        );

    \I__9481\ : Span4Mux_v
    port map (
            O => \N__43734\,
            I => \N__43731\
        );

    \I__9480\ : Odrv4
    port map (
            O => \N__43731\,
            I => \sDAC_mem_14Z0Z_2\
        );

    \I__9479\ : InMux
    port map (
            O => \N__43728\,
            I => \N__43725\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__43725\,
            I => \N__43722\
        );

    \I__9477\ : Span4Mux_h
    port map (
            O => \N__43722\,
            I => \N__43719\
        );

    \I__9476\ : Odrv4
    port map (
            O => \N__43719\,
            I => \sDAC_mem_14Z0Z_3\
        );

    \I__9475\ : InMux
    port map (
            O => \N__43716\,
            I => \N__43713\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__43713\,
            I => \N__43710\
        );

    \I__9473\ : Odrv12
    port map (
            O => \N__43710\,
            I => \sDAC_mem_40Z0Z_1\
        );

    \I__9472\ : InMux
    port map (
            O => \N__43707\,
            I => \N__43704\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__43704\,
            I => \N__43701\
        );

    \I__9470\ : Span4Mux_h
    port map (
            O => \N__43701\,
            I => \N__43698\
        );

    \I__9469\ : Span4Mux_v
    port map (
            O => \N__43698\,
            I => \N__43695\
        );

    \I__9468\ : Odrv4
    port map (
            O => \N__43695\,
            I => \sDAC_mem_8Z0Z_1\
        );

    \I__9467\ : CascadeMux
    port map (
            O => \N__43692\,
            I => \sDAC_data_2_20_am_1_4_cascade_\
        );

    \I__9466\ : CascadeMux
    port map (
            O => \N__43689\,
            I => \N__43683\
        );

    \I__9465\ : CascadeMux
    port map (
            O => \N__43688\,
            I => \N__43679\
        );

    \I__9464\ : CascadeMux
    port map (
            O => \N__43687\,
            I => \N__43675\
        );

    \I__9463\ : CascadeMux
    port map (
            O => \N__43686\,
            I => \N__43662\
        );

    \I__9462\ : InMux
    port map (
            O => \N__43683\,
            I => \N__43659\
        );

    \I__9461\ : InMux
    port map (
            O => \N__43682\,
            I => \N__43654\
        );

    \I__9460\ : InMux
    port map (
            O => \N__43679\,
            I => \N__43654\
        );

    \I__9459\ : InMux
    port map (
            O => \N__43678\,
            I => \N__43647\
        );

    \I__9458\ : InMux
    port map (
            O => \N__43675\,
            I => \N__43647\
        );

    \I__9457\ : InMux
    port map (
            O => \N__43674\,
            I => \N__43647\
        );

    \I__9456\ : CascadeMux
    port map (
            O => \N__43673\,
            I => \N__43644\
        );

    \I__9455\ : CascadeMux
    port map (
            O => \N__43672\,
            I => \N__43641\
        );

    \I__9454\ : CascadeMux
    port map (
            O => \N__43671\,
            I => \N__43638\
        );

    \I__9453\ : CascadeMux
    port map (
            O => \N__43670\,
            I => \N__43630\
        );

    \I__9452\ : CascadeMux
    port map (
            O => \N__43669\,
            I => \N__43625\
        );

    \I__9451\ : CascadeMux
    port map (
            O => \N__43668\,
            I => \N__43617\
        );

    \I__9450\ : CascadeMux
    port map (
            O => \N__43667\,
            I => \N__43614\
        );

    \I__9449\ : CascadeMux
    port map (
            O => \N__43666\,
            I => \N__43611\
        );

    \I__9448\ : CascadeMux
    port map (
            O => \N__43665\,
            I => \N__43608\
        );

    \I__9447\ : InMux
    port map (
            O => \N__43662\,
            I => \N__43603\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__43659\,
            I => \N__43596\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__43654\,
            I => \N__43596\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__43647\,
            I => \N__43596\
        );

    \I__9443\ : InMux
    port map (
            O => \N__43644\,
            I => \N__43591\
        );

    \I__9442\ : InMux
    port map (
            O => \N__43641\,
            I => \N__43591\
        );

    \I__9441\ : InMux
    port map (
            O => \N__43638\,
            I => \N__43588\
        );

    \I__9440\ : CascadeMux
    port map (
            O => \N__43637\,
            I => \N__43585\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__43636\,
            I => \N__43582\
        );

    \I__9438\ : CascadeMux
    port map (
            O => \N__43635\,
            I => \N__43572\
        );

    \I__9437\ : CascadeMux
    port map (
            O => \N__43634\,
            I => \N__43569\
        );

    \I__9436\ : CascadeMux
    port map (
            O => \N__43633\,
            I => \N__43566\
        );

    \I__9435\ : InMux
    port map (
            O => \N__43630\,
            I => \N__43559\
        );

    \I__9434\ : InMux
    port map (
            O => \N__43629\,
            I => \N__43559\
        );

    \I__9433\ : InMux
    port map (
            O => \N__43628\,
            I => \N__43556\
        );

    \I__9432\ : InMux
    port map (
            O => \N__43625\,
            I => \N__43551\
        );

    \I__9431\ : InMux
    port map (
            O => \N__43624\,
            I => \N__43551\
        );

    \I__9430\ : CascadeMux
    port map (
            O => \N__43623\,
            I => \N__43547\
        );

    \I__9429\ : CascadeMux
    port map (
            O => \N__43622\,
            I => \N__43544\
        );

    \I__9428\ : CascadeMux
    port map (
            O => \N__43621\,
            I => \N__43539\
        );

    \I__9427\ : CascadeMux
    port map (
            O => \N__43620\,
            I => \N__43536\
        );

    \I__9426\ : InMux
    port map (
            O => \N__43617\,
            I => \N__43533\
        );

    \I__9425\ : InMux
    port map (
            O => \N__43614\,
            I => \N__43528\
        );

    \I__9424\ : InMux
    port map (
            O => \N__43611\,
            I => \N__43528\
        );

    \I__9423\ : InMux
    port map (
            O => \N__43608\,
            I => \N__43521\
        );

    \I__9422\ : InMux
    port map (
            O => \N__43607\,
            I => \N__43521\
        );

    \I__9421\ : InMux
    port map (
            O => \N__43606\,
            I => \N__43521\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__43603\,
            I => \N__43508\
        );

    \I__9419\ : Span4Mux_v
    port map (
            O => \N__43596\,
            I => \N__43508\
        );

    \I__9418\ : LocalMux
    port map (
            O => \N__43591\,
            I => \N__43503\
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__43588\,
            I => \N__43503\
        );

    \I__9416\ : InMux
    port map (
            O => \N__43585\,
            I => \N__43495\
        );

    \I__9415\ : InMux
    port map (
            O => \N__43582\,
            I => \N__43495\
        );

    \I__9414\ : InMux
    port map (
            O => \N__43581\,
            I => \N__43492\
        );

    \I__9413\ : InMux
    port map (
            O => \N__43580\,
            I => \N__43489\
        );

    \I__9412\ : InMux
    port map (
            O => \N__43579\,
            I => \N__43480\
        );

    \I__9411\ : InMux
    port map (
            O => \N__43578\,
            I => \N__43480\
        );

    \I__9410\ : InMux
    port map (
            O => \N__43577\,
            I => \N__43480\
        );

    \I__9409\ : InMux
    port map (
            O => \N__43576\,
            I => \N__43480\
        );

    \I__9408\ : CascadeMux
    port map (
            O => \N__43575\,
            I => \N__43476\
        );

    \I__9407\ : InMux
    port map (
            O => \N__43572\,
            I => \N__43473\
        );

    \I__9406\ : InMux
    port map (
            O => \N__43569\,
            I => \N__43468\
        );

    \I__9405\ : InMux
    port map (
            O => \N__43566\,
            I => \N__43468\
        );

    \I__9404\ : CascadeMux
    port map (
            O => \N__43565\,
            I => \N__43465\
        );

    \I__9403\ : CascadeMux
    port map (
            O => \N__43564\,
            I => \N__43462\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__43559\,
            I => \N__43455\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__43556\,
            I => \N__43455\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__43551\,
            I => \N__43455\
        );

    \I__9399\ : CascadeMux
    port map (
            O => \N__43550\,
            I => \N__43452\
        );

    \I__9398\ : InMux
    port map (
            O => \N__43547\,
            I => \N__43441\
        );

    \I__9397\ : InMux
    port map (
            O => \N__43544\,
            I => \N__43441\
        );

    \I__9396\ : InMux
    port map (
            O => \N__43543\,
            I => \N__43441\
        );

    \I__9395\ : InMux
    port map (
            O => \N__43542\,
            I => \N__43434\
        );

    \I__9394\ : InMux
    port map (
            O => \N__43539\,
            I => \N__43434\
        );

    \I__9393\ : InMux
    port map (
            O => \N__43536\,
            I => \N__43434\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__43533\,
            I => \N__43429\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__43528\,
            I => \N__43429\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__43521\,
            I => \N__43426\
        );

    \I__9389\ : InMux
    port map (
            O => \N__43520\,
            I => \N__43417\
        );

    \I__9388\ : InMux
    port map (
            O => \N__43519\,
            I => \N__43417\
        );

    \I__9387\ : InMux
    port map (
            O => \N__43518\,
            I => \N__43417\
        );

    \I__9386\ : InMux
    port map (
            O => \N__43517\,
            I => \N__43417\
        );

    \I__9385\ : InMux
    port map (
            O => \N__43516\,
            I => \N__43408\
        );

    \I__9384\ : InMux
    port map (
            O => \N__43515\,
            I => \N__43408\
        );

    \I__9383\ : InMux
    port map (
            O => \N__43514\,
            I => \N__43408\
        );

    \I__9382\ : InMux
    port map (
            O => \N__43513\,
            I => \N__43408\
        );

    \I__9381\ : Span4Mux_h
    port map (
            O => \N__43508\,
            I => \N__43403\
        );

    \I__9380\ : Span4Mux_h
    port map (
            O => \N__43503\,
            I => \N__43403\
        );

    \I__9379\ : InMux
    port map (
            O => \N__43502\,
            I => \N__43396\
        );

    \I__9378\ : InMux
    port map (
            O => \N__43501\,
            I => \N__43396\
        );

    \I__9377\ : InMux
    port map (
            O => \N__43500\,
            I => \N__43396\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__43495\,
            I => \N__43387\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__43492\,
            I => \N__43387\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__43489\,
            I => \N__43387\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__43480\,
            I => \N__43387\
        );

    \I__9372\ : InMux
    port map (
            O => \N__43479\,
            I => \N__43384\
        );

    \I__9371\ : InMux
    port map (
            O => \N__43476\,
            I => \N__43381\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__43473\,
            I => \N__43376\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__43468\,
            I => \N__43376\
        );

    \I__9368\ : InMux
    port map (
            O => \N__43465\,
            I => \N__43371\
        );

    \I__9367\ : InMux
    port map (
            O => \N__43462\,
            I => \N__43371\
        );

    \I__9366\ : Span4Mux_v
    port map (
            O => \N__43455\,
            I => \N__43368\
        );

    \I__9365\ : InMux
    port map (
            O => \N__43452\,
            I => \N__43365\
        );

    \I__9364\ : InMux
    port map (
            O => \N__43451\,
            I => \N__43356\
        );

    \I__9363\ : InMux
    port map (
            O => \N__43450\,
            I => \N__43356\
        );

    \I__9362\ : InMux
    port map (
            O => \N__43449\,
            I => \N__43356\
        );

    \I__9361\ : InMux
    port map (
            O => \N__43448\,
            I => \N__43356\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__43441\,
            I => \N__43353\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__43434\,
            I => \N__43344\
        );

    \I__9358\ : Span4Mux_v
    port map (
            O => \N__43429\,
            I => \N__43344\
        );

    \I__9357\ : Span4Mux_h
    port map (
            O => \N__43426\,
            I => \N__43344\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__43417\,
            I => \N__43344\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__43408\,
            I => \N__43337\
        );

    \I__9354\ : Span4Mux_v
    port map (
            O => \N__43403\,
            I => \N__43337\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__43396\,
            I => \N__43337\
        );

    \I__9352\ : Span4Mux_h
    port map (
            O => \N__43387\,
            I => \N__43334\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__43384\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__43381\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9349\ : Odrv4
    port map (
            O => \N__43376\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__43371\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9347\ : Odrv4
    port map (
            O => \N__43368\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__43365\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__43356\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9344\ : Odrv12
    port map (
            O => \N__43353\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9343\ : Odrv4
    port map (
            O => \N__43344\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9342\ : Odrv4
    port map (
            O => \N__43337\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9341\ : Odrv4
    port map (
            O => \N__43334\,
            I => \sDAC_mem_pointerZ0Z_5\
        );

    \I__9340\ : CascadeMux
    port map (
            O => \N__43311\,
            I => \sDAC_data_RNO_17Z0Z_4_cascade_\
        );

    \I__9339\ : CascadeMux
    port map (
            O => \N__43308\,
            I => \sDAC_data_RNO_8Z0Z_4_cascade_\
        );

    \I__9338\ : InMux
    port map (
            O => \N__43305\,
            I => \N__43302\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__43302\,
            I => \sDAC_data_RNO_7Z0Z_4\
        );

    \I__9336\ : InMux
    port map (
            O => \N__43299\,
            I => \N__43296\
        );

    \I__9335\ : LocalMux
    port map (
            O => \N__43296\,
            I => \N__43293\
        );

    \I__9334\ : Odrv4
    port map (
            O => \N__43293\,
            I => \sDAC_data_RNO_2Z0Z_4\
        );

    \I__9333\ : CascadeMux
    port map (
            O => \N__43290\,
            I => \N_284_cascade_\
        );

    \I__9332\ : InMux
    port map (
            O => \N__43287\,
            I => \N__43284\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__43284\,
            I => \N__43278\
        );

    \I__9330\ : InMux
    port map (
            O => \N__43283\,
            I => \N__43273\
        );

    \I__9329\ : InMux
    port map (
            O => \N__43282\,
            I => \N__43273\
        );

    \I__9328\ : InMux
    port map (
            O => \N__43281\,
            I => \N__43270\
        );

    \I__9327\ : Span4Mux_v
    port map (
            O => \N__43278\,
            I => \N__43266\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__43273\,
            I => \N__43261\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__43270\,
            I => \N__43261\
        );

    \I__9324\ : InMux
    port map (
            O => \N__43269\,
            I => \N__43257\
        );

    \I__9323\ : Span4Mux_h
    port map (
            O => \N__43266\,
            I => \N__43249\
        );

    \I__9322\ : Span4Mux_v
    port map (
            O => \N__43261\,
            I => \N__43249\
        );

    \I__9321\ : InMux
    port map (
            O => \N__43260\,
            I => \N__43246\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__43257\,
            I => \N__43243\
        );

    \I__9319\ : InMux
    port map (
            O => \N__43256\,
            I => \N__43238\
        );

    \I__9318\ : InMux
    port map (
            O => \N__43255\,
            I => \N__43238\
        );

    \I__9317\ : InMux
    port map (
            O => \N__43254\,
            I => \N__43235\
        );

    \I__9316\ : Span4Mux_h
    port map (
            O => \N__43249\,
            I => \N__43230\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__43246\,
            I => \N__43230\
        );

    \I__9314\ : Span4Mux_h
    port map (
            O => \N__43243\,
            I => \N__43227\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__43238\,
            I => \N__43222\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__43235\,
            I => \N__43219\
        );

    \I__9311\ : Span4Mux_v
    port map (
            O => \N__43230\,
            I => \N__43216\
        );

    \I__9310\ : Span4Mux_h
    port map (
            O => \N__43227\,
            I => \N__43213\
        );

    \I__9309\ : InMux
    port map (
            O => \N__43226\,
            I => \N__43208\
        );

    \I__9308\ : InMux
    port map (
            O => \N__43225\,
            I => \N__43208\
        );

    \I__9307\ : Sp12to4
    port map (
            O => \N__43222\,
            I => \N__43205\
        );

    \I__9306\ : Span4Mux_v
    port map (
            O => \N__43219\,
            I => \N__43200\
        );

    \I__9305\ : Span4Mux_h
    port map (
            O => \N__43216\,
            I => \N__43200\
        );

    \I__9304\ : Odrv4
    port map (
            O => \N__43213\,
            I => \N_284\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__43208\,
            I => \N_284\
        );

    \I__9302\ : Odrv12
    port map (
            O => \N__43205\,
            I => \N_284\
        );

    \I__9301\ : Odrv4
    port map (
            O => \N__43200\,
            I => \N_284\
        );

    \I__9300\ : InMux
    port map (
            O => \N__43191\,
            I => \N__43186\
        );

    \I__9299\ : InMux
    port map (
            O => \N__43190\,
            I => \N__43183\
        );

    \I__9298\ : InMux
    port map (
            O => \N__43189\,
            I => \N__43180\
        );

    \I__9297\ : LocalMux
    port map (
            O => \N__43186\,
            I => \N__43174\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__43183\,
            I => \N__43171\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__43180\,
            I => \N__43168\
        );

    \I__9294\ : InMux
    port map (
            O => \N__43179\,
            I => \N__43161\
        );

    \I__9293\ : InMux
    port map (
            O => \N__43178\,
            I => \N__43161\
        );

    \I__9292\ : InMux
    port map (
            O => \N__43177\,
            I => \N__43161\
        );

    \I__9291\ : Span4Mux_h
    port map (
            O => \N__43174\,
            I => \N__43157\
        );

    \I__9290\ : Span4Mux_v
    port map (
            O => \N__43171\,
            I => \N__43154\
        );

    \I__9289\ : Span4Mux_v
    port map (
            O => \N__43168\,
            I => \N__43149\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__43161\,
            I => \N__43149\
        );

    \I__9287\ : InMux
    port map (
            O => \N__43160\,
            I => \N__43146\
        );

    \I__9286\ : Span4Mux_h
    port map (
            O => \N__43157\,
            I => \N__43135\
        );

    \I__9285\ : Span4Mux_h
    port map (
            O => \N__43154\,
            I => \N__43130\
        );

    \I__9284\ : Span4Mux_h
    port map (
            O => \N__43149\,
            I => \N__43130\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__43146\,
            I => \N__43127\
        );

    \I__9282\ : InMux
    port map (
            O => \N__43145\,
            I => \N__43120\
        );

    \I__9281\ : InMux
    port map (
            O => \N__43144\,
            I => \N__43120\
        );

    \I__9280\ : InMux
    port map (
            O => \N__43143\,
            I => \N__43120\
        );

    \I__9279\ : InMux
    port map (
            O => \N__43142\,
            I => \N__43115\
        );

    \I__9278\ : InMux
    port map (
            O => \N__43141\,
            I => \N__43115\
        );

    \I__9277\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43108\
        );

    \I__9276\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43108\
        );

    \I__9275\ : InMux
    port map (
            O => \N__43138\,
            I => \N__43108\
        );

    \I__9274\ : Odrv4
    port map (
            O => \N__43135\,
            I => \N_280\
        );

    \I__9273\ : Odrv4
    port map (
            O => \N__43130\,
            I => \N_280\
        );

    \I__9272\ : Odrv4
    port map (
            O => \N__43127\,
            I => \N_280\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__43120\,
            I => \N_280\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__43115\,
            I => \N_280\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__43108\,
            I => \N_280\
        );

    \I__9268\ : InMux
    port map (
            O => \N__43095\,
            I => \N__43092\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__43092\,
            I => \sDAC_mem_6Z0Z_6\
        );

    \I__9266\ : CEMux
    port map (
            O => \N__43089\,
            I => \N__43086\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__43086\,
            I => \N__43082\
        );

    \I__9264\ : CEMux
    port map (
            O => \N__43085\,
            I => \N__43079\
        );

    \I__9263\ : Span4Mux_v
    port map (
            O => \N__43082\,
            I => \N__43075\
        );

    \I__9262\ : LocalMux
    port map (
            O => \N__43079\,
            I => \N__43072\
        );

    \I__9261\ : CEMux
    port map (
            O => \N__43078\,
            I => \N__43068\
        );

    \I__9260\ : Span4Mux_v
    port map (
            O => \N__43075\,
            I => \N__43063\
        );

    \I__9259\ : Span4Mux_v
    port map (
            O => \N__43072\,
            I => \N__43063\
        );

    \I__9258\ : CEMux
    port map (
            O => \N__43071\,
            I => \N__43060\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__43068\,
            I => \N__43057\
        );

    \I__9256\ : Sp12to4
    port map (
            O => \N__43063\,
            I => \N__43054\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__43060\,
            I => \N__43051\
        );

    \I__9254\ : Span4Mux_h
    port map (
            O => \N__43057\,
            I => \N__43048\
        );

    \I__9253\ : Odrv12
    port map (
            O => \N__43054\,
            I => \sDAC_mem_6_1_sqmuxa\
        );

    \I__9252\ : Odrv4
    port map (
            O => \N__43051\,
            I => \sDAC_mem_6_1_sqmuxa\
        );

    \I__9251\ : Odrv4
    port map (
            O => \N__43048\,
            I => \sDAC_mem_6_1_sqmuxa\
        );

    \I__9250\ : InMux
    port map (
            O => \N__43041\,
            I => \N__43038\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__43038\,
            I => \N__43035\
        );

    \I__9248\ : Odrv12
    port map (
            O => \N__43035\,
            I => \sDAC_mem_40Z0Z_0\
        );

    \I__9247\ : InMux
    port map (
            O => \N__43032\,
            I => \N__43029\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__43029\,
            I => \N__43026\
        );

    \I__9245\ : Span4Mux_h
    port map (
            O => \N__43026\,
            I => \N__43023\
        );

    \I__9244\ : Span4Mux_v
    port map (
            O => \N__43023\,
            I => \N__43020\
        );

    \I__9243\ : Odrv4
    port map (
            O => \N__43020\,
            I => \sDAC_mem_8Z0Z_0\
        );

    \I__9242\ : CascadeMux
    port map (
            O => \N__43017\,
            I => \sDAC_data_2_20_am_1_3_cascade_\
        );

    \I__9241\ : CascadeMux
    port map (
            O => \N__43014\,
            I => \sDAC_data_RNO_17Z0Z_3_cascade_\
        );

    \I__9240\ : CascadeMux
    port map (
            O => \N__43011\,
            I => \sDAC_data_RNO_8Z0Z_3_cascade_\
        );

    \I__9239\ : InMux
    port map (
            O => \N__43008\,
            I => \N__43005\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__43005\,
            I => \sDAC_data_RNO_7Z0Z_3\
        );

    \I__9237\ : InMux
    port map (
            O => \N__43002\,
            I => \N__42999\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__42999\,
            I => \sDAC_data_RNO_2Z0Z_3\
        );

    \I__9235\ : CEMux
    port map (
            O => \N__42996\,
            I => \N__42993\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__42993\,
            I => \N__42989\
        );

    \I__9233\ : CEMux
    port map (
            O => \N__42992\,
            I => \N__42986\
        );

    \I__9232\ : Span4Mux_h
    port map (
            O => \N__42989\,
            I => \N__42979\
        );

    \I__9231\ : LocalMux
    port map (
            O => \N__42986\,
            I => \N__42979\
        );

    \I__9230\ : CEMux
    port map (
            O => \N__42985\,
            I => \N__42974\
        );

    \I__9229\ : CEMux
    port map (
            O => \N__42984\,
            I => \N__42971\
        );

    \I__9228\ : Span4Mux_v
    port map (
            O => \N__42979\,
            I => \N__42968\
        );

    \I__9227\ : CEMux
    port map (
            O => \N__42978\,
            I => \N__42965\
        );

    \I__9226\ : CEMux
    port map (
            O => \N__42977\,
            I => \N__42962\
        );

    \I__9225\ : LocalMux
    port map (
            O => \N__42974\,
            I => \N__42957\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__42971\,
            I => \N__42954\
        );

    \I__9223\ : Span4Mux_h
    port map (
            O => \N__42968\,
            I => \N__42951\
        );

    \I__9222\ : LocalMux
    port map (
            O => \N__42965\,
            I => \N__42948\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__42962\,
            I => \N__42945\
        );

    \I__9220\ : CEMux
    port map (
            O => \N__42961\,
            I => \N__42942\
        );

    \I__9219\ : CEMux
    port map (
            O => \N__42960\,
            I => \N__42939\
        );

    \I__9218\ : Span4Mux_h
    port map (
            O => \N__42957\,
            I => \N__42936\
        );

    \I__9217\ : Span4Mux_v
    port map (
            O => \N__42954\,
            I => \N__42933\
        );

    \I__9216\ : Span4Mux_h
    port map (
            O => \N__42951\,
            I => \N__42922\
        );

    \I__9215\ : Span4Mux_v
    port map (
            O => \N__42948\,
            I => \N__42922\
        );

    \I__9214\ : Span4Mux_h
    port map (
            O => \N__42945\,
            I => \N__42922\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__42942\,
            I => \N__42922\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__42939\,
            I => \N__42922\
        );

    \I__9211\ : Span4Mux_v
    port map (
            O => \N__42936\,
            I => \N__42919\
        );

    \I__9210\ : Span4Mux_h
    port map (
            O => \N__42933\,
            I => \N__42916\
        );

    \I__9209\ : Sp12to4
    port map (
            O => \N__42922\,
            I => \N__42913\
        );

    \I__9208\ : Odrv4
    port map (
            O => \N__42919\,
            I => \sDAC_mem_3_1_sqmuxa\
        );

    \I__9207\ : Odrv4
    port map (
            O => \N__42916\,
            I => \sDAC_mem_3_1_sqmuxa\
        );

    \I__9206\ : Odrv12
    port map (
            O => \N__42913\,
            I => \sDAC_mem_3_1_sqmuxa\
        );

    \I__9205\ : CascadeMux
    port map (
            O => \N__42906\,
            I => \N__42903\
        );

    \I__9204\ : InMux
    port map (
            O => \N__42903\,
            I => \N__42900\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__42900\,
            I => \N__42897\
        );

    \I__9202\ : Span4Mux_v
    port map (
            O => \N__42897\,
            I => \N__42894\
        );

    \I__9201\ : Span4Mux_h
    port map (
            O => \N__42894\,
            I => \N__42891\
        );

    \I__9200\ : Span4Mux_v
    port map (
            O => \N__42891\,
            I => \N__42888\
        );

    \I__9199\ : Odrv4
    port map (
            O => \N__42888\,
            I => \sDAC_mem_34Z0Z_7\
        );

    \I__9198\ : InMux
    port map (
            O => \N__42885\,
            I => \N__42882\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__42882\,
            I => \N__42879\
        );

    \I__9196\ : Span4Mux_v
    port map (
            O => \N__42879\,
            I => \N__42876\
        );

    \I__9195\ : Span4Mux_h
    port map (
            O => \N__42876\,
            I => \N__42873\
        );

    \I__9194\ : Odrv4
    port map (
            O => \N__42873\,
            I => \sDAC_mem_2Z0Z_7\
        );

    \I__9193\ : InMux
    port map (
            O => \N__42870\,
            I => \N__42867\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__42867\,
            I => \N__42864\
        );

    \I__9191\ : Span4Mux_v
    port map (
            O => \N__42864\,
            I => \N__42861\
        );

    \I__9190\ : Odrv4
    port map (
            O => \N__42861\,
            I => \sDAC_mem_35Z0Z_7\
        );

    \I__9189\ : CascadeMux
    port map (
            O => \N__42858\,
            I => \sDAC_data_2_6_bm_1_10_cascade_\
        );

    \I__9188\ : InMux
    port map (
            O => \N__42855\,
            I => \N__42852\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__42852\,
            I => \sDAC_mem_3Z0Z_7\
        );

    \I__9186\ : CascadeMux
    port map (
            O => \N__42849\,
            I => \N__42846\
        );

    \I__9185\ : InMux
    port map (
            O => \N__42846\,
            I => \N__42843\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__42843\,
            I => \N__42840\
        );

    \I__9183\ : Odrv4
    port map (
            O => \N__42840\,
            I => \sDAC_data_RNO_15Z0Z_10\
        );

    \I__9182\ : InMux
    port map (
            O => \N__42837\,
            I => \N__42834\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__42834\,
            I => \N__42831\
        );

    \I__9180\ : Span4Mux_v
    port map (
            O => \N__42831\,
            I => \N__42828\
        );

    \I__9179\ : Odrv4
    port map (
            O => \N__42828\,
            I => \sDAC_mem_35Z0Z_3\
        );

    \I__9178\ : CascadeMux
    port map (
            O => \N__42825\,
            I => \sDAC_data_2_6_bm_1_6_cascade_\
        );

    \I__9177\ : InMux
    port map (
            O => \N__42822\,
            I => \N__42819\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__42819\,
            I => \sDAC_mem_3Z0Z_3\
        );

    \I__9175\ : CascadeMux
    port map (
            O => \N__42816\,
            I => \N__42813\
        );

    \I__9174\ : InMux
    port map (
            O => \N__42813\,
            I => \N__42810\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__42810\,
            I => \sDAC_data_RNO_15Z0Z_6\
        );

    \I__9172\ : CascadeMux
    port map (
            O => \N__42807\,
            I => \sDAC_data_RNO_17Z0Z_8_cascade_\
        );

    \I__9171\ : InMux
    port map (
            O => \N__42804\,
            I => \N__42801\
        );

    \I__9170\ : LocalMux
    port map (
            O => \N__42801\,
            I => \N__42798\
        );

    \I__9169\ : Odrv12
    port map (
            O => \N__42798\,
            I => \sDAC_mem_40Z0Z_5\
        );

    \I__9168\ : InMux
    port map (
            O => \N__42795\,
            I => \N__42792\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__42792\,
            I => \N__42789\
        );

    \I__9166\ : Span4Mux_v
    port map (
            O => \N__42789\,
            I => \N__42786\
        );

    \I__9165\ : Odrv4
    port map (
            O => \N__42786\,
            I => \sDAC_mem_8Z0Z_5\
        );

    \I__9164\ : CascadeMux
    port map (
            O => \N__42783\,
            I => \sDAC_data_2_20_am_1_8_cascade_\
        );

    \I__9163\ : CascadeMux
    port map (
            O => \N__42780\,
            I => \sDAC_data_RNO_7Z0Z_8_cascade_\
        );

    \I__9162\ : InMux
    port map (
            O => \N__42777\,
            I => \N__42774\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__42774\,
            I => \sDAC_data_RNO_8Z0Z_8\
        );

    \I__9160\ : InMux
    port map (
            O => \N__42771\,
            I => \N__42768\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__42768\,
            I => \sDAC_data_RNO_2Z0Z_8\
        );

    \I__9158\ : InMux
    port map (
            O => \N__42765\,
            I => \N__42762\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__42762\,
            I => \N__42759\
        );

    \I__9156\ : Odrv12
    port map (
            O => \N__42759\,
            I => \sDAC_mem_38Z0Z_6\
        );

    \I__9155\ : InMux
    port map (
            O => \N__42756\,
            I => \N__42753\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__42753\,
            I => \N__42750\
        );

    \I__9153\ : Span4Mux_v
    port map (
            O => \N__42750\,
            I => \N__42747\
        );

    \I__9152\ : Odrv4
    port map (
            O => \N__42747\,
            I => \sDAC_mem_39Z0Z_6\
        );

    \I__9151\ : CascadeMux
    port map (
            O => \N__42744\,
            I => \sDAC_data_2_13_bm_1_9_cascade_\
        );

    \I__9150\ : InMux
    port map (
            O => \N__42741\,
            I => \N__42738\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__42738\,
            I => \N__42735\
        );

    \I__9148\ : Span4Mux_h
    port map (
            O => \N__42735\,
            I => \N__42732\
        );

    \I__9147\ : Span4Mux_v
    port map (
            O => \N__42732\,
            I => \N__42729\
        );

    \I__9146\ : Odrv4
    port map (
            O => \N__42729\,
            I => \sDAC_mem_7Z0Z_6\
        );

    \I__9145\ : InMux
    port map (
            O => \N__42726\,
            I => \N__42723\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__42723\,
            I => \N__42720\
        );

    \I__9143\ : Span4Mux_v
    port map (
            O => \N__42720\,
            I => \N__42717\
        );

    \I__9142\ : Odrv4
    port map (
            O => \N__42717\,
            I => \sDAC_data_RNO_5Z0Z_9\
        );

    \I__9141\ : InMux
    port map (
            O => \N__42714\,
            I => \N__42711\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__42711\,
            I => \sDAC_data_RNO_14Z0Z_6\
        );

    \I__9139\ : InMux
    port map (
            O => \N__42708\,
            I => \N__42705\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__42705\,
            I => \sDAC_data_2_14_ns_1_6\
        );

    \I__9137\ : CascadeMux
    port map (
            O => \N__42702\,
            I => \N__42699\
        );

    \I__9136\ : InMux
    port map (
            O => \N__42699\,
            I => \N__42696\
        );

    \I__9135\ : LocalMux
    port map (
            O => \N__42696\,
            I => \N__42693\
        );

    \I__9134\ : Span4Mux_h
    port map (
            O => \N__42693\,
            I => \N__42690\
        );

    \I__9133\ : Span4Mux_v
    port map (
            O => \N__42690\,
            I => \N__42687\
        );

    \I__9132\ : Span4Mux_v
    port map (
            O => \N__42687\,
            I => \N__42684\
        );

    \I__9131\ : Odrv4
    port map (
            O => \N__42684\,
            I => \sDAC_data_RNO_29Z0Z_6\
        );

    \I__9130\ : InMux
    port map (
            O => \N__42681\,
            I => \N__42678\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__42678\,
            I => \N__42675\
        );

    \I__9128\ : Span4Mux_h
    port map (
            O => \N__42675\,
            I => \N__42672\
        );

    \I__9127\ : Odrv4
    port map (
            O => \N__42672\,
            I => \sDAC_data_RNO_30Z0Z_6\
        );

    \I__9126\ : InMux
    port map (
            O => \N__42669\,
            I => \N__42666\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__42666\,
            I => \N__42663\
        );

    \I__9124\ : Span4Mux_h
    port map (
            O => \N__42663\,
            I => \N__42660\
        );

    \I__9123\ : Span4Mux_h
    port map (
            O => \N__42660\,
            I => \N__42657\
        );

    \I__9122\ : Odrv4
    port map (
            O => \N__42657\,
            I => \sDAC_data_RNO_21Z0Z_6\
        );

    \I__9121\ : CascadeMux
    port map (
            O => \N__42654\,
            I => \sDAC_data_2_32_ns_1_6_cascade_\
        );

    \I__9120\ : InMux
    port map (
            O => \N__42651\,
            I => \N__42648\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__42648\,
            I => \N__42645\
        );

    \I__9118\ : Odrv4
    port map (
            O => \N__42645\,
            I => \sDAC_data_RNO_20Z0Z_6\
        );

    \I__9117\ : InMux
    port map (
            O => \N__42642\,
            I => \N__42635\
        );

    \I__9116\ : InMux
    port map (
            O => \N__42641\,
            I => \N__42632\
        );

    \I__9115\ : InMux
    port map (
            O => \N__42640\,
            I => \N__42627\
        );

    \I__9114\ : InMux
    port map (
            O => \N__42639\,
            I => \N__42624\
        );

    \I__9113\ : InMux
    port map (
            O => \N__42638\,
            I => \N__42620\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__42635\,
            I => \N__42615\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__42632\,
            I => \N__42615\
        );

    \I__9110\ : InMux
    port map (
            O => \N__42631\,
            I => \N__42611\
        );

    \I__9109\ : InMux
    port map (
            O => \N__42630\,
            I => \N__42607\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__42627\,
            I => \N__42604\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__42624\,
            I => \N__42601\
        );

    \I__9106\ : InMux
    port map (
            O => \N__42623\,
            I => \N__42598\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__42620\,
            I => \N__42595\
        );

    \I__9104\ : Span4Mux_v
    port map (
            O => \N__42615\,
            I => \N__42592\
        );

    \I__9103\ : CascadeMux
    port map (
            O => \N__42614\,
            I => \N__42589\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__42611\,
            I => \N__42586\
        );

    \I__9101\ : InMux
    port map (
            O => \N__42610\,
            I => \N__42583\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__42607\,
            I => \N__42576\
        );

    \I__9099\ : Span4Mux_h
    port map (
            O => \N__42604\,
            I => \N__42576\
        );

    \I__9098\ : Span4Mux_h
    port map (
            O => \N__42601\,
            I => \N__42576\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__42598\,
            I => \N__42569\
        );

    \I__9096\ : Span4Mux_v
    port map (
            O => \N__42595\,
            I => \N__42569\
        );

    \I__9095\ : Span4Mux_h
    port map (
            O => \N__42592\,
            I => \N__42569\
        );

    \I__9094\ : InMux
    port map (
            O => \N__42589\,
            I => \N__42566\
        );

    \I__9093\ : Odrv12
    port map (
            O => \N__42586\,
            I => \sDAC_mem_pointerZ0Z_3\
        );

    \I__9092\ : LocalMux
    port map (
            O => \N__42583\,
            I => \sDAC_mem_pointerZ0Z_3\
        );

    \I__9091\ : Odrv4
    port map (
            O => \N__42576\,
            I => \sDAC_mem_pointerZ0Z_3\
        );

    \I__9090\ : Odrv4
    port map (
            O => \N__42569\,
            I => \sDAC_mem_pointerZ0Z_3\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__42566\,
            I => \sDAC_mem_pointerZ0Z_3\
        );

    \I__9088\ : CascadeMux
    port map (
            O => \N__42555\,
            I => \sDAC_data_RNO_10Z0Z_6_cascade_\
        );

    \I__9087\ : InMux
    port map (
            O => \N__42552\,
            I => \N__42549\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__42549\,
            I => \N__42546\
        );

    \I__9085\ : Span4Mux_h
    port map (
            O => \N__42546\,
            I => \N__42543\
        );

    \I__9084\ : Span4Mux_v
    port map (
            O => \N__42543\,
            I => \N__42540\
        );

    \I__9083\ : Span4Mux_h
    port map (
            O => \N__42540\,
            I => \N__42537\
        );

    \I__9082\ : Odrv4
    port map (
            O => \N__42537\,
            I => \sDAC_data_RNO_11Z0Z_6\
        );

    \I__9081\ : CascadeMux
    port map (
            O => \N__42534\,
            I => \N__42519\
        );

    \I__9080\ : InMux
    port map (
            O => \N__42533\,
            I => \N__42514\
        );

    \I__9079\ : InMux
    port map (
            O => \N__42532\,
            I => \N__42511\
        );

    \I__9078\ : InMux
    port map (
            O => \N__42531\,
            I => \N__42508\
        );

    \I__9077\ : InMux
    port map (
            O => \N__42530\,
            I => \N__42505\
        );

    \I__9076\ : InMux
    port map (
            O => \N__42529\,
            I => \N__42500\
        );

    \I__9075\ : InMux
    port map (
            O => \N__42528\,
            I => \N__42500\
        );

    \I__9074\ : InMux
    port map (
            O => \N__42527\,
            I => \N__42497\
        );

    \I__9073\ : InMux
    port map (
            O => \N__42526\,
            I => \N__42492\
        );

    \I__9072\ : InMux
    port map (
            O => \N__42525\,
            I => \N__42492\
        );

    \I__9071\ : InMux
    port map (
            O => \N__42524\,
            I => \N__42489\
        );

    \I__9070\ : InMux
    port map (
            O => \N__42523\,
            I => \N__42484\
        );

    \I__9069\ : InMux
    port map (
            O => \N__42522\,
            I => \N__42484\
        );

    \I__9068\ : InMux
    port map (
            O => \N__42519\,
            I => \N__42480\
        );

    \I__9067\ : InMux
    port map (
            O => \N__42518\,
            I => \N__42476\
        );

    \I__9066\ : InMux
    port map (
            O => \N__42517\,
            I => \N__42473\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__42514\,
            I => \N__42470\
        );

    \I__9064\ : LocalMux
    port map (
            O => \N__42511\,
            I => \N__42467\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__42508\,
            I => \N__42464\
        );

    \I__9062\ : LocalMux
    port map (
            O => \N__42505\,
            I => \N__42461\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__42500\,
            I => \N__42458\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__42497\,
            I => \N__42451\
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__42492\,
            I => \N__42451\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__42489\,
            I => \N__42451\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__42484\,
            I => \N__42448\
        );

    \I__9056\ : InMux
    port map (
            O => \N__42483\,
            I => \N__42444\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__42480\,
            I => \N__42441\
        );

    \I__9054\ : InMux
    port map (
            O => \N__42479\,
            I => \N__42438\
        );

    \I__9053\ : LocalMux
    port map (
            O => \N__42476\,
            I => \N__42429\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__42473\,
            I => \N__42429\
        );

    \I__9051\ : Span4Mux_v
    port map (
            O => \N__42470\,
            I => \N__42429\
        );

    \I__9050\ : Span4Mux_v
    port map (
            O => \N__42467\,
            I => \N__42429\
        );

    \I__9049\ : Span4Mux_h
    port map (
            O => \N__42464\,
            I => \N__42426\
        );

    \I__9048\ : Span4Mux_v
    port map (
            O => \N__42461\,
            I => \N__42417\
        );

    \I__9047\ : Span4Mux_v
    port map (
            O => \N__42458\,
            I => \N__42417\
        );

    \I__9046\ : Span4Mux_v
    port map (
            O => \N__42451\,
            I => \N__42417\
        );

    \I__9045\ : Span4Mux_v
    port map (
            O => \N__42448\,
            I => \N__42417\
        );

    \I__9044\ : InMux
    port map (
            O => \N__42447\,
            I => \N__42414\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__42444\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__9042\ : Odrv12
    port map (
            O => \N__42441\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__42438\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__9040\ : Odrv4
    port map (
            O => \N__42429\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__9039\ : Odrv4
    port map (
            O => \N__42426\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__9038\ : Odrv4
    port map (
            O => \N__42417\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__42414\,
            I => \sDAC_mem_pointerZ0Z_4\
        );

    \I__9036\ : InMux
    port map (
            O => \N__42399\,
            I => \N__42396\
        );

    \I__9035\ : LocalMux
    port map (
            O => \N__42396\,
            I => \sDAC_data_RNO_2Z0Z_6\
        );

    \I__9034\ : CascadeMux
    port map (
            O => \N__42393\,
            I => \sDAC_data_2_41_ns_1_6_cascade_\
        );

    \I__9033\ : InMux
    port map (
            O => \N__42390\,
            I => \N__42387\
        );

    \I__9032\ : LocalMux
    port map (
            O => \N__42387\,
            I => \sDAC_data_RNO_1Z0Z_6\
        );

    \I__9031\ : InMux
    port map (
            O => \N__42384\,
            I => \N__42370\
        );

    \I__9030\ : InMux
    port map (
            O => \N__42383\,
            I => \N__42367\
        );

    \I__9029\ : InMux
    port map (
            O => \N__42382\,
            I => \N__42363\
        );

    \I__9028\ : InMux
    port map (
            O => \N__42381\,
            I => \N__42360\
        );

    \I__9027\ : InMux
    port map (
            O => \N__42380\,
            I => \N__42357\
        );

    \I__9026\ : InMux
    port map (
            O => \N__42379\,
            I => \N__42354\
        );

    \I__9025\ : InMux
    port map (
            O => \N__42378\,
            I => \N__42351\
        );

    \I__9024\ : InMux
    port map (
            O => \N__42377\,
            I => \N__42348\
        );

    \I__9023\ : InMux
    port map (
            O => \N__42376\,
            I => \N__42345\
        );

    \I__9022\ : InMux
    port map (
            O => \N__42375\,
            I => \N__42338\
        );

    \I__9021\ : InMux
    port map (
            O => \N__42374\,
            I => \N__42338\
        );

    \I__9020\ : InMux
    port map (
            O => \N__42373\,
            I => \N__42338\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__42370\,
            I => \N__42333\
        );

    \I__9018\ : LocalMux
    port map (
            O => \N__42367\,
            I => \N__42333\
        );

    \I__9017\ : InMux
    port map (
            O => \N__42366\,
            I => \N__42330\
        );

    \I__9016\ : LocalMux
    port map (
            O => \N__42363\,
            I => \N__42325\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__42360\,
            I => \N__42325\
        );

    \I__9014\ : LocalMux
    port map (
            O => \N__42357\,
            I => \N__42322\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__42354\,
            I => \N__42315\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__42351\,
            I => \N__42315\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__42348\,
            I => \N__42315\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__42345\,
            I => \N__42308\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__42338\,
            I => \N__42308\
        );

    \I__9008\ : Span4Mux_h
    port map (
            O => \N__42333\,
            I => \N__42308\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__42330\,
            I => \N__42305\
        );

    \I__9006\ : Span4Mux_h
    port map (
            O => \N__42325\,
            I => \N__42302\
        );

    \I__9005\ : Span4Mux_v
    port map (
            O => \N__42322\,
            I => \N__42299\
        );

    \I__9004\ : Span4Mux_h
    port map (
            O => \N__42315\,
            I => \N__42295\
        );

    \I__9003\ : Span4Mux_v
    port map (
            O => \N__42308\,
            I => \N__42292\
        );

    \I__9002\ : Span4Mux_h
    port map (
            O => \N__42305\,
            I => \N__42289\
        );

    \I__9001\ : Span4Mux_v
    port map (
            O => \N__42302\,
            I => \N__42286\
        );

    \I__9000\ : Span4Mux_v
    port map (
            O => \N__42299\,
            I => \N__42283\
        );

    \I__8999\ : InMux
    port map (
            O => \N__42298\,
            I => \N__42280\
        );

    \I__8998\ : Span4Mux_v
    port map (
            O => \N__42295\,
            I => \N__42277\
        );

    \I__8997\ : Span4Mux_v
    port map (
            O => \N__42292\,
            I => \N__42274\
        );

    \I__8996\ : Span4Mux_v
    port map (
            O => \N__42289\,
            I => \N__42269\
        );

    \I__8995\ : Span4Mux_v
    port map (
            O => \N__42286\,
            I => \N__42269\
        );

    \I__8994\ : Span4Mux_v
    port map (
            O => \N__42283\,
            I => \N__42266\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__42280\,
            I => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\
        );

    \I__8992\ : Odrv4
    port map (
            O => \N__42277\,
            I => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\
        );

    \I__8991\ : Odrv4
    port map (
            O => \N__42274\,
            I => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\
        );

    \I__8990\ : Odrv4
    port map (
            O => \N__42269\,
            I => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\
        );

    \I__8989\ : Odrv4
    port map (
            O => \N__42266\,
            I => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\
        );

    \I__8988\ : CascadeMux
    port map (
            O => \N__42255\,
            I => \sDAC_data_2_6_cascade_\
        );

    \I__8987\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42249\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__42249\,
            I => \N__42246\
        );

    \I__8985\ : Span4Mux_h
    port map (
            O => \N__42246\,
            I => \N__42243\
        );

    \I__8984\ : Span4Mux_v
    port map (
            O => \N__42243\,
            I => \N__42240\
        );

    \I__8983\ : Span4Mux_h
    port map (
            O => \N__42240\,
            I => \N__42237\
        );

    \I__8982\ : Odrv4
    port map (
            O => \N__42237\,
            I => \sDAC_dataZ0Z_6\
        );

    \I__8981\ : CEMux
    port map (
            O => \N__42234\,
            I => \N__42192\
        );

    \I__8980\ : CEMux
    port map (
            O => \N__42233\,
            I => \N__42192\
        );

    \I__8979\ : CEMux
    port map (
            O => \N__42232\,
            I => \N__42192\
        );

    \I__8978\ : CEMux
    port map (
            O => \N__42231\,
            I => \N__42192\
        );

    \I__8977\ : CEMux
    port map (
            O => \N__42230\,
            I => \N__42192\
        );

    \I__8976\ : CEMux
    port map (
            O => \N__42229\,
            I => \N__42192\
        );

    \I__8975\ : CEMux
    port map (
            O => \N__42228\,
            I => \N__42192\
        );

    \I__8974\ : CEMux
    port map (
            O => \N__42227\,
            I => \N__42192\
        );

    \I__8973\ : CEMux
    port map (
            O => \N__42226\,
            I => \N__42192\
        );

    \I__8972\ : CEMux
    port map (
            O => \N__42225\,
            I => \N__42192\
        );

    \I__8971\ : CEMux
    port map (
            O => \N__42224\,
            I => \N__42192\
        );

    \I__8970\ : CEMux
    port map (
            O => \N__42223\,
            I => \N__42192\
        );

    \I__8969\ : CEMux
    port map (
            O => \N__42222\,
            I => \N__42192\
        );

    \I__8968\ : CEMux
    port map (
            O => \N__42221\,
            I => \N__42192\
        );

    \I__8967\ : GlobalMux
    port map (
            O => \N__42192\,
            I => \N__42189\
        );

    \I__8966\ : gio2CtrlBuf
    port map (
            O => \N__42189\,
            I => op_eq_scounterdac10_g
        );

    \I__8965\ : CascadeMux
    port map (
            O => \N__42186\,
            I => \N__42183\
        );

    \I__8964\ : InMux
    port map (
            O => \N__42183\,
            I => \N__42180\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__42180\,
            I => \N__42177\
        );

    \I__8962\ : Span12Mux_v
    port map (
            O => \N__42177\,
            I => \N__42174\
        );

    \I__8961\ : Odrv12
    port map (
            O => \N__42174\,
            I => \sDAC_mem_2Z0Z_3\
        );

    \I__8960\ : InMux
    port map (
            O => \N__42171\,
            I => \N__42168\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__42168\,
            I => \N__42165\
        );

    \I__8958\ : Span4Mux_v
    port map (
            O => \N__42165\,
            I => \N__42162\
        );

    \I__8957\ : Odrv4
    port map (
            O => \N__42162\,
            I => \sDAC_mem_34Z0Z_3\
        );

    \I__8956\ : InMux
    port map (
            O => \N__42159\,
            I => \N__42156\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__42156\,
            I => \N__42153\
        );

    \I__8954\ : Span4Mux_h
    port map (
            O => \N__42153\,
            I => \N__42150\
        );

    \I__8953\ : Odrv4
    port map (
            O => \N__42150\,
            I => \sDAC_mem_33Z0Z_3\
        );

    \I__8952\ : CascadeMux
    port map (
            O => \N__42147\,
            I => \sDAC_data_RNO_26Z0Z_6_cascade_\
        );

    \I__8951\ : CascadeMux
    port map (
            O => \N__42144\,
            I => \N__42140\
        );

    \I__8950\ : CascadeMux
    port map (
            O => \N__42143\,
            I => \N__42137\
        );

    \I__8949\ : InMux
    port map (
            O => \N__42140\,
            I => \N__42132\
        );

    \I__8948\ : InMux
    port map (
            O => \N__42137\,
            I => \N__42132\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__42132\,
            I => \N__42129\
        );

    \I__8946\ : Span4Mux_v
    port map (
            O => \N__42129\,
            I => \N__42126\
        );

    \I__8945\ : Span4Mux_h
    port map (
            O => \N__42126\,
            I => \N__42123\
        );

    \I__8944\ : Odrv4
    port map (
            O => \N__42123\,
            I => \sDAC_mem_32Z0Z_3\
        );

    \I__8943\ : InMux
    port map (
            O => \N__42120\,
            I => \N__42117\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__42117\,
            I => \sDAC_data_RNO_27Z0Z_6\
        );

    \I__8941\ : InMux
    port map (
            O => \N__42114\,
            I => \N__42108\
        );

    \I__8940\ : InMux
    port map (
            O => \N__42113\,
            I => \N__42108\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__42108\,
            I => \sDAC_mem_1Z0Z_3\
        );

    \I__8938\ : InMux
    port map (
            O => \N__42105\,
            I => \N__42102\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__42102\,
            I => \N__42099\
        );

    \I__8936\ : Odrv12
    port map (
            O => \N__42099\,
            I => \sDAC_mem_33Z0Z_4\
        );

    \I__8935\ : CascadeMux
    port map (
            O => \N__42096\,
            I => \sDAC_data_RNO_26Z0Z_7_cascade_\
        );

    \I__8934\ : CascadeMux
    port map (
            O => \N__42093\,
            I => \N__42090\
        );

    \I__8933\ : InMux
    port map (
            O => \N__42090\,
            I => \N__42087\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__42087\,
            I => \N__42084\
        );

    \I__8931\ : Span4Mux_h
    port map (
            O => \N__42084\,
            I => \N__42081\
        );

    \I__8930\ : Odrv4
    port map (
            O => \N__42081\,
            I => \sDAC_data_RNO_14Z0Z_7\
        );

    \I__8929\ : CascadeMux
    port map (
            O => \N__42078\,
            I => \N__42074\
        );

    \I__8928\ : CascadeMux
    port map (
            O => \N__42077\,
            I => \N__42071\
        );

    \I__8927\ : InMux
    port map (
            O => \N__42074\,
            I => \N__42066\
        );

    \I__8926\ : InMux
    port map (
            O => \N__42071\,
            I => \N__42066\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__42066\,
            I => \N__42063\
        );

    \I__8924\ : Span4Mux_h
    port map (
            O => \N__42063\,
            I => \N__42060\
        );

    \I__8923\ : Span4Mux_h
    port map (
            O => \N__42060\,
            I => \N__42057\
        );

    \I__8922\ : Odrv4
    port map (
            O => \N__42057\,
            I => \sDAC_mem_32Z0Z_4\
        );

    \I__8921\ : InMux
    port map (
            O => \N__42054\,
            I => \N__42051\
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__42051\,
            I => \sDAC_data_RNO_27Z0Z_7\
        );

    \I__8919\ : InMux
    port map (
            O => \N__42048\,
            I => \N__42042\
        );

    \I__8918\ : InMux
    port map (
            O => \N__42047\,
            I => \N__42042\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__42042\,
            I => \sDAC_mem_1Z0Z_4\
        );

    \I__8916\ : CEMux
    port map (
            O => \N__42039\,
            I => \N__42036\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__42036\,
            I => \N__42033\
        );

    \I__8914\ : Span4Mux_h
    port map (
            O => \N__42033\,
            I => \N__42028\
        );

    \I__8913\ : CEMux
    port map (
            O => \N__42032\,
            I => \N__42025\
        );

    \I__8912\ : CEMux
    port map (
            O => \N__42031\,
            I => \N__42022\
        );

    \I__8911\ : Odrv4
    port map (
            O => \N__42028\,
            I => \sDAC_mem_1_1_sqmuxa\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__42025\,
            I => \sDAC_mem_1_1_sqmuxa\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__42022\,
            I => \sDAC_mem_1_1_sqmuxa\
        );

    \I__8908\ : InMux
    port map (
            O => \N__42015\,
            I => \N__42012\
        );

    \I__8907\ : LocalMux
    port map (
            O => \N__42012\,
            I => \sDAC_data_RNO_5Z0Z_6\
        );

    \I__8906\ : InMux
    port map (
            O => \N__42009\,
            I => \N__42006\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__42006\,
            I => \N__42003\
        );

    \I__8904\ : Span4Mux_v
    port map (
            O => \N__42003\,
            I => \N__42000\
        );

    \I__8903\ : Odrv4
    port map (
            O => \N__42000\,
            I => \sDAC_data_RNO_4Z0Z_6\
        );

    \I__8902\ : InMux
    port map (
            O => \N__41997\,
            I => \N__41994\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__41994\,
            I => \N__41991\
        );

    \I__8900\ : Span12Mux_v
    port map (
            O => \N__41991\,
            I => \N__41988\
        );

    \I__8899\ : Odrv12
    port map (
            O => \N__41988\,
            I => \sDAC_mem_40Z0Z_7\
        );

    \I__8898\ : CEMux
    port map (
            O => \N__41985\,
            I => \N__41982\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__41982\,
            I => \N__41979\
        );

    \I__8896\ : Span4Mux_h
    port map (
            O => \N__41979\,
            I => \N__41976\
        );

    \I__8895\ : Odrv4
    port map (
            O => \N__41976\,
            I => \sDAC_mem_40_1_sqmuxa\
        );

    \I__8894\ : InMux
    port map (
            O => \N__41973\,
            I => \N__41970\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__41970\,
            I => \sDAC_mem_21Z0Z_0\
        );

    \I__8892\ : InMux
    port map (
            O => \N__41967\,
            I => \N__41964\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__41964\,
            I => \N__41961\
        );

    \I__8890\ : Span4Mux_v
    port map (
            O => \N__41961\,
            I => \N__41958\
        );

    \I__8889\ : Odrv4
    port map (
            O => \N__41958\,
            I => \sDAC_data_RNO_20Z0Z_3\
        );

    \I__8888\ : InMux
    port map (
            O => \N__41955\,
            I => \N__41952\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__41952\,
            I => \sDAC_mem_20Z0Z_0\
        );

    \I__8886\ : InMux
    port map (
            O => \N__41949\,
            I => \N__41946\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__41946\,
            I => \sDAC_mem_21Z0Z_1\
        );

    \I__8884\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41940\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__41940\,
            I => \N__41937\
        );

    \I__8882\ : Span4Mux_v
    port map (
            O => \N__41937\,
            I => \N__41934\
        );

    \I__8881\ : Odrv4
    port map (
            O => \N__41934\,
            I => \sDAC_data_RNO_20Z0Z_4\
        );

    \I__8880\ : InMux
    port map (
            O => \N__41931\,
            I => \N__41928\
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__41928\,
            I => \sDAC_mem_20Z0Z_1\
        );

    \I__8878\ : InMux
    port map (
            O => \N__41925\,
            I => \N__41922\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__41922\,
            I => \sDAC_mem_21Z0Z_2\
        );

    \I__8876\ : InMux
    port map (
            O => \N__41919\,
            I => \N__41916\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__41916\,
            I => \N__41913\
        );

    \I__8874\ : Odrv12
    port map (
            O => \N__41913\,
            I => \sDAC_data_RNO_20Z0Z_5\
        );

    \I__8873\ : InMux
    port map (
            O => \N__41910\,
            I => \N__41907\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__41907\,
            I => \sDAC_mem_20Z0Z_2\
        );

    \I__8871\ : InMux
    port map (
            O => \N__41904\,
            I => \N__41901\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__41901\,
            I => \N__41898\
        );

    \I__8869\ : Odrv4
    port map (
            O => \N__41898\,
            I => \sDAC_mem_21Z0Z_3\
        );

    \I__8868\ : InMux
    port map (
            O => \N__41895\,
            I => \N__41892\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__41892\,
            I => \sDAC_mem_20Z0Z_3\
        );

    \I__8866\ : InMux
    port map (
            O => \N__41889\,
            I => \N__41886\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__41886\,
            I => \N__41883\
        );

    \I__8864\ : Odrv4
    port map (
            O => \N__41883\,
            I => \sDAC_mem_38Z0Z_5\
        );

    \I__8863\ : InMux
    port map (
            O => \N__41880\,
            I => \N__41877\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__41877\,
            I => \N__41874\
        );

    \I__8861\ : Span4Mux_v
    port map (
            O => \N__41874\,
            I => \N__41871\
        );

    \I__8860\ : Odrv4
    port map (
            O => \N__41871\,
            I => \sDAC_mem_38Z0Z_7\
        );

    \I__8859\ : CEMux
    port map (
            O => \N__41868\,
            I => \N__41863\
        );

    \I__8858\ : CEMux
    port map (
            O => \N__41867\,
            I => \N__41860\
        );

    \I__8857\ : CEMux
    port map (
            O => \N__41866\,
            I => \N__41857\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__41863\,
            I => \N__41854\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__41860\,
            I => \N__41851\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__41857\,
            I => \N__41848\
        );

    \I__8853\ : Span4Mux_h
    port map (
            O => \N__41854\,
            I => \N__41845\
        );

    \I__8852\ : Span4Mux_v
    port map (
            O => \N__41851\,
            I => \N__41842\
        );

    \I__8851\ : Span4Mux_v
    port map (
            O => \N__41848\,
            I => \N__41839\
        );

    \I__8850\ : Odrv4
    port map (
            O => \N__41845\,
            I => \sDAC_mem_38_1_sqmuxa\
        );

    \I__8849\ : Odrv4
    port map (
            O => \N__41842\,
            I => \sDAC_mem_38_1_sqmuxa\
        );

    \I__8848\ : Odrv4
    port map (
            O => \N__41839\,
            I => \sDAC_mem_38_1_sqmuxa\
        );

    \I__8847\ : InMux
    port map (
            O => \N__41832\,
            I => \N__41829\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__41829\,
            I => \N__41826\
        );

    \I__8845\ : Span4Mux_h
    port map (
            O => \N__41826\,
            I => \N__41823\
        );

    \I__8844\ : Odrv4
    port map (
            O => \N__41823\,
            I => \sDAC_mem_40Z0Z_2\
        );

    \I__8843\ : InMux
    port map (
            O => \N__41820\,
            I => \N__41817\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__41817\,
            I => \N__41814\
        );

    \I__8841\ : Span4Mux_v
    port map (
            O => \N__41814\,
            I => \N__41811\
        );

    \I__8840\ : Odrv4
    port map (
            O => \N__41811\,
            I => \sDAC_mem_40Z0Z_3\
        );

    \I__8839\ : InMux
    port map (
            O => \N__41808\,
            I => \N__41805\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__41805\,
            I => \N__41802\
        );

    \I__8837\ : Span4Mux_h
    port map (
            O => \N__41802\,
            I => \N__41799\
        );

    \I__8836\ : Odrv4
    port map (
            O => \N__41799\,
            I => \sDAC_mem_40Z0Z_4\
        );

    \I__8835\ : InMux
    port map (
            O => \N__41796\,
            I => \N__41793\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__41793\,
            I => \N__41790\
        );

    \I__8833\ : Span4Mux_h
    port map (
            O => \N__41790\,
            I => \N__41787\
        );

    \I__8832\ : Odrv4
    port map (
            O => \N__41787\,
            I => \sDAC_mem_40Z0Z_6\
        );

    \I__8831\ : InMux
    port map (
            O => \N__41784\,
            I => \N__41781\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__41781\,
            I => \sDAC_mem_28Z0Z_7\
        );

    \I__8829\ : CEMux
    port map (
            O => \N__41778\,
            I => \N__41773\
        );

    \I__8828\ : CEMux
    port map (
            O => \N__41777\,
            I => \N__41769\
        );

    \I__8827\ : CEMux
    port map (
            O => \N__41776\,
            I => \N__41766\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__41773\,
            I => \N__41763\
        );

    \I__8825\ : CEMux
    port map (
            O => \N__41772\,
            I => \N__41760\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__41769\,
            I => \N__41757\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__41766\,
            I => \N__41754\
        );

    \I__8822\ : Span4Mux_v
    port map (
            O => \N__41763\,
            I => \N__41751\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__41760\,
            I => \N__41748\
        );

    \I__8820\ : Span4Mux_v
    port map (
            O => \N__41757\,
            I => \N__41745\
        );

    \I__8819\ : Odrv4
    port map (
            O => \N__41754\,
            I => \sDAC_mem_28_1_sqmuxa\
        );

    \I__8818\ : Odrv4
    port map (
            O => \N__41751\,
            I => \sDAC_mem_28_1_sqmuxa\
        );

    \I__8817\ : Odrv4
    port map (
            O => \N__41748\,
            I => \sDAC_mem_28_1_sqmuxa\
        );

    \I__8816\ : Odrv4
    port map (
            O => \N__41745\,
            I => \sDAC_mem_28_1_sqmuxa\
        );

    \I__8815\ : InMux
    port map (
            O => \N__41736\,
            I => \N__41733\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__41733\,
            I => \N__41730\
        );

    \I__8813\ : Odrv4
    port map (
            O => \N__41730\,
            I => \sDAC_mem_25Z0Z_1\
        );

    \I__8812\ : CEMux
    port map (
            O => \N__41727\,
            I => \N__41724\
        );

    \I__8811\ : LocalMux
    port map (
            O => \N__41724\,
            I => \N__41720\
        );

    \I__8810\ : CEMux
    port map (
            O => \N__41723\,
            I => \N__41717\
        );

    \I__8809\ : Span4Mux_v
    port map (
            O => \N__41720\,
            I => \N__41713\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__41717\,
            I => \N__41710\
        );

    \I__8807\ : CEMux
    port map (
            O => \N__41716\,
            I => \N__41707\
        );

    \I__8806\ : Span4Mux_h
    port map (
            O => \N__41713\,
            I => \N__41702\
        );

    \I__8805\ : Span4Mux_v
    port map (
            O => \N__41710\,
            I => \N__41702\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__41707\,
            I => \N__41699\
        );

    \I__8803\ : Odrv4
    port map (
            O => \N__41702\,
            I => \sDAC_mem_25_1_sqmuxa\
        );

    \I__8802\ : Odrv4
    port map (
            O => \N__41699\,
            I => \sDAC_mem_25_1_sqmuxa\
        );

    \I__8801\ : InMux
    port map (
            O => \N__41694\,
            I => \N__41691\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__41691\,
            I => \N__41688\
        );

    \I__8799\ : Span4Mux_v
    port map (
            O => \N__41688\,
            I => \N__41685\
        );

    \I__8798\ : Span4Mux_h
    port map (
            O => \N__41685\,
            I => \N__41682\
        );

    \I__8797\ : Span4Mux_v
    port map (
            O => \N__41682\,
            I => \N__41679\
        );

    \I__8796\ : Odrv4
    port map (
            O => \N__41679\,
            I => \sDAC_mem_17Z0Z_1\
        );

    \I__8795\ : CascadeMux
    port map (
            O => \N__41676\,
            I => \N__41673\
        );

    \I__8794\ : InMux
    port map (
            O => \N__41673\,
            I => \N__41670\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__41670\,
            I => \N__41667\
        );

    \I__8792\ : Span12Mux_s11_h
    port map (
            O => \N__41667\,
            I => \N__41664\
        );

    \I__8791\ : Odrv12
    port map (
            O => \N__41664\,
            I => \sDAC_data_RNO_29Z0Z_4\
        );

    \I__8790\ : InMux
    port map (
            O => \N__41661\,
            I => \N__41658\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__41658\,
            I => \N__41655\
        );

    \I__8788\ : Span4Mux_v
    port map (
            O => \N__41655\,
            I => \N__41652\
        );

    \I__8787\ : Span4Mux_h
    port map (
            O => \N__41652\,
            I => \N__41649\
        );

    \I__8786\ : Odrv4
    port map (
            O => \N__41649\,
            I => \sDAC_mem_38Z0Z_0\
        );

    \I__8785\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41643\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__41643\,
            I => \N__41640\
        );

    \I__8783\ : Span4Mux_h
    port map (
            O => \N__41640\,
            I => \N__41637\
        );

    \I__8782\ : Odrv4
    port map (
            O => \N__41637\,
            I => \sDAC_mem_38Z0Z_2\
        );

    \I__8781\ : InMux
    port map (
            O => \N__41634\,
            I => \N__41631\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__41631\,
            I => \N__41628\
        );

    \I__8779\ : Odrv4
    port map (
            O => \N__41628\,
            I => \sDAC_mem_38Z0Z_3\
        );

    \I__8778\ : InMux
    port map (
            O => \N__41625\,
            I => \N__41622\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__41622\,
            I => \N__41619\
        );

    \I__8776\ : Span4Mux_h
    port map (
            O => \N__41619\,
            I => \N__41616\
        );

    \I__8775\ : Odrv4
    port map (
            O => \N__41616\,
            I => \sDAC_mem_38Z0Z_4\
        );

    \I__8774\ : InMux
    port map (
            O => \N__41613\,
            I => \N__41610\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__41610\,
            I => \sDAC_mem_28Z0Z_0\
        );

    \I__8772\ : InMux
    port map (
            O => \N__41607\,
            I => \N__41604\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__41604\,
            I => \N__41601\
        );

    \I__8770\ : Span4Mux_h
    port map (
            O => \N__41601\,
            I => \N__41598\
        );

    \I__8769\ : Odrv4
    port map (
            O => \N__41598\,
            I => \sDAC_mem_24Z0Z_1\
        );

    \I__8768\ : CascadeMux
    port map (
            O => \N__41595\,
            I => \sDAC_data_RNO_31Z0Z_4_cascade_\
        );

    \I__8767\ : InMux
    port map (
            O => \N__41592\,
            I => \N__41589\
        );

    \I__8766\ : LocalMux
    port map (
            O => \N__41589\,
            I => \sDAC_data_RNO_24Z0Z_4\
        );

    \I__8765\ : CascadeMux
    port map (
            O => \N__41586\,
            I => \sDAC_data_2_39_ns_1_4_cascade_\
        );

    \I__8764\ : InMux
    port map (
            O => \N__41583\,
            I => \N__41580\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__41580\,
            I => \sDAC_data_RNO_23Z0Z_4\
        );

    \I__8762\ : InMux
    port map (
            O => \N__41577\,
            I => \N__41574\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__41574\,
            I => \N__41571\
        );

    \I__8760\ : Odrv12
    port map (
            O => \N__41571\,
            I => \sDAC_data_RNO_11Z0Z_4\
        );

    \I__8759\ : InMux
    port map (
            O => \N__41568\,
            I => \N__41565\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__41565\,
            I => \N__41562\
        );

    \I__8757\ : Span4Mux_v
    port map (
            O => \N__41562\,
            I => \N__41559\
        );

    \I__8756\ : Odrv4
    port map (
            O => \N__41559\,
            I => \sDAC_mem_26Z0Z_1\
        );

    \I__8755\ : InMux
    port map (
            O => \N__41556\,
            I => \N__41553\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__41553\,
            I => \N__41550\
        );

    \I__8753\ : Odrv4
    port map (
            O => \N__41550\,
            I => \sDAC_mem_27Z0Z_1\
        );

    \I__8752\ : InMux
    port map (
            O => \N__41547\,
            I => \N__41544\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__41544\,
            I => \sDAC_data_RNO_32Z0Z_4\
        );

    \I__8750\ : InMux
    port map (
            O => \N__41541\,
            I => \N__41538\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__41538\,
            I => \sDAC_mem_28Z0Z_1\
        );

    \I__8748\ : InMux
    port map (
            O => \N__41535\,
            I => \N__41532\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__41532\,
            I => \N__41529\
        );

    \I__8746\ : Span4Mux_h
    port map (
            O => \N__41529\,
            I => \N__41526\
        );

    \I__8745\ : Odrv4
    port map (
            O => \N__41526\,
            I => \sDAC_mem_28Z0Z_2\
        );

    \I__8744\ : InMux
    port map (
            O => \N__41523\,
            I => \N__41520\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__41520\,
            I => \N__41517\
        );

    \I__8742\ : Span4Mux_v
    port map (
            O => \N__41517\,
            I => \N__41514\
        );

    \I__8741\ : Odrv4
    port map (
            O => \N__41514\,
            I => \sDAC_mem_28Z0Z_4\
        );

    \I__8740\ : InMux
    port map (
            O => \N__41511\,
            I => \N__41508\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__41508\,
            I => \N__41505\
        );

    \I__8738\ : Span4Mux_h
    port map (
            O => \N__41505\,
            I => \N__41502\
        );

    \I__8737\ : Odrv4
    port map (
            O => \N__41502\,
            I => \sDAC_mem_28Z0Z_5\
        );

    \I__8736\ : InMux
    port map (
            O => \N__41499\,
            I => \N__41496\
        );

    \I__8735\ : LocalMux
    port map (
            O => \N__41496\,
            I => \N__41493\
        );

    \I__8734\ : Span4Mux_h
    port map (
            O => \N__41493\,
            I => \N__41490\
        );

    \I__8733\ : Odrv4
    port map (
            O => \N__41490\,
            I => \sDAC_mem_27Z0Z_5\
        );

    \I__8732\ : InMux
    port map (
            O => \N__41487\,
            I => \N__41484\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__41484\,
            I => \N__41481\
        );

    \I__8730\ : Span4Mux_v
    port map (
            O => \N__41481\,
            I => \N__41478\
        );

    \I__8729\ : Span4Mux_h
    port map (
            O => \N__41478\,
            I => \N__41475\
        );

    \I__8728\ : Odrv4
    port map (
            O => \N__41475\,
            I => \sDAC_mem_27Z0Z_6\
        );

    \I__8727\ : CascadeMux
    port map (
            O => \N__41472\,
            I => \N__41469\
        );

    \I__8726\ : InMux
    port map (
            O => \N__41469\,
            I => \N__41466\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__41466\,
            I => \N__41463\
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__41463\,
            I => \sDAC_mem_27Z0Z_7\
        );

    \I__8723\ : InMux
    port map (
            O => \N__41460\,
            I => \N__41457\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__41457\,
            I => \N__41454\
        );

    \I__8721\ : Odrv12
    port map (
            O => \N__41454\,
            I => \sEEADC_freqZ0Z_0\
        );

    \I__8720\ : InMux
    port map (
            O => \N__41451\,
            I => \N__41448\
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__41448\,
            I => \N__41445\
        );

    \I__8718\ : Odrv12
    port map (
            O => \N__41445\,
            I => \sEEADC_freqZ0Z_6\
        );

    \I__8717\ : CascadeMux
    port map (
            O => \N__41442\,
            I => \N__41439\
        );

    \I__8716\ : InMux
    port map (
            O => \N__41439\,
            I => \N__41436\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__41436\,
            I => \N__41433\
        );

    \I__8714\ : Span4Mux_h
    port map (
            O => \N__41433\,
            I => \N__41430\
        );

    \I__8713\ : Odrv4
    port map (
            O => \N__41430\,
            I => \sEEADC_freqZ0Z_7\
        );

    \I__8712\ : InMux
    port map (
            O => \N__41427\,
            I => \N__41424\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__41424\,
            I => \N__41421\
        );

    \I__8710\ : Span4Mux_h
    port map (
            O => \N__41421\,
            I => \N__41418\
        );

    \I__8709\ : Odrv4
    port map (
            O => \N__41418\,
            I => \sDAC_mem_31Z0Z_0\
        );

    \I__8708\ : InMux
    port map (
            O => \N__41415\,
            I => \N__41412\
        );

    \I__8707\ : LocalMux
    port map (
            O => \N__41412\,
            I => \sDAC_mem_30Z0Z_0\
        );

    \I__8706\ : InMux
    port map (
            O => \N__41409\,
            I => \N__41406\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__41406\,
            I => \N__41403\
        );

    \I__8704\ : Odrv4
    port map (
            O => \N__41403\,
            I => \sDAC_mem_29Z0Z_0\
        );

    \I__8703\ : InMux
    port map (
            O => \N__41400\,
            I => \N__41397\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__41397\,
            I => \sDAC_data_RNO_24Z0Z_3\
        );

    \I__8701\ : CascadeMux
    port map (
            O => \N__41394\,
            I => \sDAC_data_RNO_23Z0Z_3_cascade_\
        );

    \I__8700\ : InMux
    port map (
            O => \N__41391\,
            I => \N__41388\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__41388\,
            I => \sDAC_data_2_39_ns_1_3\
        );

    \I__8698\ : InMux
    port map (
            O => \N__41385\,
            I => \N__41382\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__41382\,
            I => \N__41379\
        );

    \I__8696\ : Span4Mux_h
    port map (
            O => \N__41379\,
            I => \N__41376\
        );

    \I__8695\ : Odrv4
    port map (
            O => \N__41376\,
            I => \sDAC_data_RNO_11Z0Z_3\
        );

    \I__8694\ : CascadeMux
    port map (
            O => \N__41373\,
            I => \sDAC_data_2_3_cascade_\
        );

    \I__8693\ : InMux
    port map (
            O => \N__41370\,
            I => \N__41367\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__41367\,
            I => \N__41364\
        );

    \I__8691\ : Span4Mux_v
    port map (
            O => \N__41364\,
            I => \N__41361\
        );

    \I__8690\ : Span4Mux_h
    port map (
            O => \N__41361\,
            I => \N__41358\
        );

    \I__8689\ : Span4Mux_v
    port map (
            O => \N__41358\,
            I => \N__41355\
        );

    \I__8688\ : Odrv4
    port map (
            O => \N__41355\,
            I => \sDAC_dataZ0Z_3\
        );

    \I__8687\ : InMux
    port map (
            O => \N__41352\,
            I => \N__41349\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__41349\,
            I => \N__41346\
        );

    \I__8685\ : Span4Mux_v
    port map (
            O => \N__41346\,
            I => \N__41343\
        );

    \I__8684\ : Span4Mux_h
    port map (
            O => \N__41343\,
            I => \N__41340\
        );

    \I__8683\ : Odrv4
    port map (
            O => \N__41340\,
            I => \sDAC_mem_16Z0Z_7\
        );

    \I__8682\ : InMux
    port map (
            O => \N__41337\,
            I => \N__41334\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__41334\,
            I => \N__41331\
        );

    \I__8680\ : Span4Mux_h
    port map (
            O => \N__41331\,
            I => \N__41328\
        );

    \I__8679\ : Span4Mux_v
    port map (
            O => \N__41328\,
            I => \N__41325\
        );

    \I__8678\ : Odrv4
    port map (
            O => \N__41325\,
            I => \sDAC_mem_17Z0Z_7\
        );

    \I__8677\ : InMux
    port map (
            O => \N__41322\,
            I => \N__41319\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__41319\,
            I => \sDAC_data_RNO_29Z0Z_10\
        );

    \I__8675\ : InMux
    port map (
            O => \N__41316\,
            I => \N__41313\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__41313\,
            I => \N__41310\
        );

    \I__8673\ : Span4Mux_h
    port map (
            O => \N__41310\,
            I => \N__41307\
        );

    \I__8672\ : Odrv4
    port map (
            O => \N__41307\,
            I => \sDAC_mem_19Z0Z_3\
        );

    \I__8671\ : InMux
    port map (
            O => \N__41304\,
            I => \N__41301\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__41301\,
            I => \N__41298\
        );

    \I__8669\ : Odrv12
    port map (
            O => \N__41298\,
            I => \sDAC_mem_18Z0Z_3\
        );

    \I__8668\ : InMux
    port map (
            O => \N__41295\,
            I => \N__41292\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__41292\,
            I => \N__41289\
        );

    \I__8666\ : Span4Mux_v
    port map (
            O => \N__41289\,
            I => \N__41286\
        );

    \I__8665\ : Span4Mux_h
    port map (
            O => \N__41286\,
            I => \N__41283\
        );

    \I__8664\ : Odrv4
    port map (
            O => \N__41283\,
            I => \sDAC_mem_23Z0Z_1\
        );

    \I__8663\ : InMux
    port map (
            O => \N__41280\,
            I => \N__41277\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__41277\,
            I => \N__41274\
        );

    \I__8661\ : Span4Mux_h
    port map (
            O => \N__41274\,
            I => \N__41271\
        );

    \I__8660\ : Span4Mux_v
    port map (
            O => \N__41271\,
            I => \N__41268\
        );

    \I__8659\ : Odrv4
    port map (
            O => \N__41268\,
            I => \sDAC_mem_22Z0Z_1\
        );

    \I__8658\ : InMux
    port map (
            O => \N__41265\,
            I => \N__41262\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__41262\,
            I => \N__41259\
        );

    \I__8656\ : Odrv12
    port map (
            O => \N__41259\,
            I => \sDAC_data_RNO_21Z0Z_4\
        );

    \I__8655\ : InMux
    port map (
            O => \N__41256\,
            I => \N__41253\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__41253\,
            I => \N__41250\
        );

    \I__8653\ : Span4Mux_v
    port map (
            O => \N__41250\,
            I => \N__41247\
        );

    \I__8652\ : Span4Mux_h
    port map (
            O => \N__41247\,
            I => \N__41244\
        );

    \I__8651\ : Odrv4
    port map (
            O => \N__41244\,
            I => \sDAC_mem_27Z0Z_2\
        );

    \I__8650\ : InMux
    port map (
            O => \N__41241\,
            I => \N__41238\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__41238\,
            I => \N__41235\
        );

    \I__8648\ : Span4Mux_h
    port map (
            O => \N__41235\,
            I => \N__41232\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__41232\,
            I => \N__41229\
        );

    \I__8646\ : Odrv4
    port map (
            O => \N__41229\,
            I => \sDAC_mem_27Z0Z_3\
        );

    \I__8645\ : InMux
    port map (
            O => \N__41226\,
            I => \N__41223\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__41223\,
            I => \N__41220\
        );

    \I__8643\ : Span4Mux_h
    port map (
            O => \N__41220\,
            I => \N__41217\
        );

    \I__8642\ : Odrv4
    port map (
            O => \N__41217\,
            I => \sDAC_mem_27Z0Z_4\
        );

    \I__8641\ : CascadeMux
    port map (
            O => \N__41214\,
            I => \sDAC_data_RNO_1Z0Z_4_cascade_\
        );

    \I__8640\ : InMux
    port map (
            O => \N__41211\,
            I => \N__41208\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__41208\,
            I => \sDAC_data_2_41_ns_1_4\
        );

    \I__8638\ : CascadeMux
    port map (
            O => \N__41205\,
            I => \sDAC_data_2_4_cascade_\
        );

    \I__8637\ : InMux
    port map (
            O => \N__41202\,
            I => \N__41199\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__41199\,
            I => \N__41196\
        );

    \I__8635\ : Span12Mux_h
    port map (
            O => \N__41196\,
            I => \N__41193\
        );

    \I__8634\ : Odrv12
    port map (
            O => \N__41193\,
            I => \sDAC_dataZ0Z_4\
        );

    \I__8633\ : InMux
    port map (
            O => \N__41190\,
            I => \N__41187\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__41187\,
            I => \N__41184\
        );

    \I__8631\ : Span4Mux_v
    port map (
            O => \N__41184\,
            I => \N__41181\
        );

    \I__8630\ : Odrv4
    port map (
            O => \N__41181\,
            I => \sDAC_data_RNO_21Z0Z_3\
        );

    \I__8629\ : CascadeMux
    port map (
            O => \N__41178\,
            I => \sDAC_data_RNO_10Z0Z_3_cascade_\
        );

    \I__8628\ : InMux
    port map (
            O => \N__41175\,
            I => \N__41172\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__41172\,
            I => \N__41169\
        );

    \I__8626\ : Odrv4
    port map (
            O => \N__41169\,
            I => \sDAC_data_RNO_30Z0Z_3\
        );

    \I__8625\ : InMux
    port map (
            O => \N__41166\,
            I => \N__41163\
        );

    \I__8624\ : LocalMux
    port map (
            O => \N__41163\,
            I => \sDAC_data_2_32_ns_1_3\
        );

    \I__8623\ : CascadeMux
    port map (
            O => \N__41160\,
            I => \N__41157\
        );

    \I__8622\ : InMux
    port map (
            O => \N__41157\,
            I => \N__41154\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__41154\,
            I => \N__41151\
        );

    \I__8620\ : Span4Mux_h
    port map (
            O => \N__41151\,
            I => \N__41148\
        );

    \I__8619\ : Sp12to4
    port map (
            O => \N__41148\,
            I => \N__41145\
        );

    \I__8618\ : Odrv12
    port map (
            O => \N__41145\,
            I => \sDAC_data_RNO_15Z0Z_3\
        );

    \I__8617\ : InMux
    port map (
            O => \N__41142\,
            I => \N__41139\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__41139\,
            I => \sDAC_data_RNO_14Z0Z_3\
        );

    \I__8615\ : InMux
    port map (
            O => \N__41136\,
            I => \N__41133\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__41133\,
            I => \N__41130\
        );

    \I__8613\ : Span4Mux_v
    port map (
            O => \N__41130\,
            I => \N__41127\
        );

    \I__8612\ : Span4Mux_v
    port map (
            O => \N__41127\,
            I => \N__41124\
        );

    \I__8611\ : Odrv4
    port map (
            O => \N__41124\,
            I => \sDAC_data_RNO_5Z0Z_3\
        );

    \I__8610\ : CascadeMux
    port map (
            O => \N__41121\,
            I => \sDAC_data_2_14_ns_1_3_cascade_\
        );

    \I__8609\ : InMux
    port map (
            O => \N__41118\,
            I => \N__41115\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__41115\,
            I => \sDAC_data_RNO_4Z0Z_3\
        );

    \I__8607\ : CascadeMux
    port map (
            O => \N__41112\,
            I => \sDAC_data_RNO_1Z0Z_3_cascade_\
        );

    \I__8606\ : InMux
    port map (
            O => \N__41109\,
            I => \N__41106\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__41106\,
            I => \sDAC_data_2_41_ns_1_3\
        );

    \I__8604\ : CascadeMux
    port map (
            O => \N__41103\,
            I => \sDAC_data_RNO_17Z0Z_6_cascade_\
        );

    \I__8603\ : InMux
    port map (
            O => \N__41100\,
            I => \N__41097\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__41097\,
            I => \N__41094\
        );

    \I__8601\ : Span4Mux_v
    port map (
            O => \N__41094\,
            I => \N__41091\
        );

    \I__8600\ : Odrv4
    port map (
            O => \N__41091\,
            I => \sDAC_mem_8Z0Z_3\
        );

    \I__8599\ : CascadeMux
    port map (
            O => \N__41088\,
            I => \sDAC_data_2_20_am_1_6_cascade_\
        );

    \I__8598\ : InMux
    port map (
            O => \N__41085\,
            I => \N__41082\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__41082\,
            I => \N__41079\
        );

    \I__8596\ : Span4Mux_v
    port map (
            O => \N__41079\,
            I => \N__41076\
        );

    \I__8595\ : Odrv4
    port map (
            O => \N__41076\,
            I => \sDAC_data_2_24_ns_1_6\
        );

    \I__8594\ : CascadeMux
    port map (
            O => \N__41073\,
            I => \sDAC_data_RNO_7Z0Z_6_cascade_\
        );

    \I__8593\ : InMux
    port map (
            O => \N__41070\,
            I => \N__41067\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__41067\,
            I => \sDAC_data_RNO_8Z0Z_6\
        );

    \I__8591\ : CascadeMux
    port map (
            O => \N__41064\,
            I => \sDAC_data_RNO_10Z0Z_4_cascade_\
        );

    \I__8590\ : InMux
    port map (
            O => \N__41061\,
            I => \N__41058\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__41058\,
            I => \N__41055\
        );

    \I__8588\ : Span4Mux_h
    port map (
            O => \N__41055\,
            I => \N__41052\
        );

    \I__8587\ : Odrv4
    port map (
            O => \N__41052\,
            I => \sDAC_data_RNO_30Z0Z_4\
        );

    \I__8586\ : InMux
    port map (
            O => \N__41049\,
            I => \N__41046\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__41046\,
            I => \sDAC_data_2_32_ns_1_4\
        );

    \I__8584\ : CascadeMux
    port map (
            O => \N__41043\,
            I => \N__41040\
        );

    \I__8583\ : InMux
    port map (
            O => \N__41040\,
            I => \N__41037\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__41037\,
            I => \N__41034\
        );

    \I__8581\ : Odrv12
    port map (
            O => \N__41034\,
            I => \sDAC_data_RNO_15Z0Z_4\
        );

    \I__8580\ : InMux
    port map (
            O => \N__41031\,
            I => \N__41028\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__41028\,
            I => \N__41025\
        );

    \I__8578\ : Span4Mux_v
    port map (
            O => \N__41025\,
            I => \N__41022\
        );

    \I__8577\ : Odrv4
    port map (
            O => \N__41022\,
            I => \sDAC_data_RNO_14Z0Z_4\
        );

    \I__8576\ : InMux
    port map (
            O => \N__41019\,
            I => \N__41016\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__41016\,
            I => \N__41013\
        );

    \I__8574\ : Span4Mux_h
    port map (
            O => \N__41013\,
            I => \N__41010\
        );

    \I__8573\ : Span4Mux_v
    port map (
            O => \N__41010\,
            I => \N__41007\
        );

    \I__8572\ : Odrv4
    port map (
            O => \N__41007\,
            I => \sDAC_data_RNO_5Z0Z_4\
        );

    \I__8571\ : CascadeMux
    port map (
            O => \N__41004\,
            I => \sDAC_data_2_14_ns_1_4_cascade_\
        );

    \I__8570\ : InMux
    port map (
            O => \N__41001\,
            I => \N__40998\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__40998\,
            I => \N__40995\
        );

    \I__8568\ : Span4Mux_h
    port map (
            O => \N__40995\,
            I => \N__40992\
        );

    \I__8567\ : Odrv4
    port map (
            O => \N__40992\,
            I => \sDAC_data_RNO_4Z0Z_4\
        );

    \I__8566\ : CascadeMux
    port map (
            O => \N__40989\,
            I => \N__40986\
        );

    \I__8565\ : InMux
    port map (
            O => \N__40986\,
            I => \N__40983\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__40983\,
            I => \N__40980\
        );

    \I__8563\ : Odrv4
    port map (
            O => \N__40980\,
            I => \sDAC_data_RNO_15Z0Z_8\
        );

    \I__8562\ : InMux
    port map (
            O => \N__40977\,
            I => \N__40974\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__40974\,
            I => \N__40971\
        );

    \I__8560\ : Odrv4
    port map (
            O => \N__40971\,
            I => \sDAC_data_RNO_14Z0Z_8\
        );

    \I__8559\ : InMux
    port map (
            O => \N__40968\,
            I => \N__40965\
        );

    \I__8558\ : LocalMux
    port map (
            O => \N__40965\,
            I => \sDAC_data_RNO_5Z0Z_8\
        );

    \I__8557\ : CascadeMux
    port map (
            O => \N__40962\,
            I => \sDAC_data_2_14_ns_1_8_cascade_\
        );

    \I__8556\ : InMux
    port map (
            O => \N__40959\,
            I => \N__40956\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__40956\,
            I => \sDAC_data_RNO_4Z0Z_8\
        );

    \I__8554\ : InMux
    port map (
            O => \N__40953\,
            I => \N__40950\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__40950\,
            I => \sDAC_data_RNO_10Z0Z_8\
        );

    \I__8552\ : CascadeMux
    port map (
            O => \N__40947\,
            I => \N__40944\
        );

    \I__8551\ : InMux
    port map (
            O => \N__40944\,
            I => \N__40941\
        );

    \I__8550\ : LocalMux
    port map (
            O => \N__40941\,
            I => \N__40938\
        );

    \I__8549\ : Span4Mux_h
    port map (
            O => \N__40938\,
            I => \N__40935\
        );

    \I__8548\ : Span4Mux_h
    port map (
            O => \N__40935\,
            I => \N__40932\
        );

    \I__8547\ : Odrv4
    port map (
            O => \N__40932\,
            I => \sDAC_data_RNO_11Z0Z_8\
        );

    \I__8546\ : CascadeMux
    port map (
            O => \N__40929\,
            I => \sDAC_data_2_41_ns_1_8_cascade_\
        );

    \I__8545\ : InMux
    port map (
            O => \N__40926\,
            I => \N__40923\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__40923\,
            I => \sDAC_data_RNO_1Z0Z_8\
        );

    \I__8543\ : CascadeMux
    port map (
            O => \N__40920\,
            I => \sDAC_data_2_8_cascade_\
        );

    \I__8542\ : InMux
    port map (
            O => \N__40917\,
            I => \N__40914\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__40914\,
            I => \N__40911\
        );

    \I__8540\ : Span4Mux_h
    port map (
            O => \N__40911\,
            I => \N__40908\
        );

    \I__8539\ : Span4Mux_h
    port map (
            O => \N__40908\,
            I => \N__40905\
        );

    \I__8538\ : Sp12to4
    port map (
            O => \N__40905\,
            I => \N__40902\
        );

    \I__8537\ : Odrv12
    port map (
            O => \N__40902\,
            I => \sDAC_dataZ0Z_8\
        );

    \I__8536\ : CascadeMux
    port map (
            O => \N__40899\,
            I => \N__40896\
        );

    \I__8535\ : InMux
    port map (
            O => \N__40896\,
            I => \N__40893\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__40893\,
            I => \N__40890\
        );

    \I__8533\ : Span4Mux_v
    port map (
            O => \N__40890\,
            I => \N__40887\
        );

    \I__8532\ : Odrv4
    port map (
            O => \N__40887\,
            I => \sDAC_mem_2Z0Z_1\
        );

    \I__8531\ : InMux
    port map (
            O => \N__40884\,
            I => \N__40881\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__40881\,
            I => \N__40878\
        );

    \I__8529\ : Odrv12
    port map (
            O => \N__40878\,
            I => \sDAC_mem_34Z0Z_1\
        );

    \I__8528\ : InMux
    port map (
            O => \N__40875\,
            I => \N__40872\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__40872\,
            I => \N__40869\
        );

    \I__8526\ : Odrv12
    port map (
            O => \N__40869\,
            I => \sDAC_mem_35Z0Z_1\
        );

    \I__8525\ : CascadeMux
    port map (
            O => \N__40866\,
            I => \sDAC_data_2_6_bm_1_4_cascade_\
        );

    \I__8524\ : InMux
    port map (
            O => \N__40863\,
            I => \N__40860\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__40860\,
            I => \sDAC_mem_3Z0Z_1\
        );

    \I__8522\ : InMux
    port map (
            O => \N__40857\,
            I => \N__40854\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__40854\,
            I => \N__40851\
        );

    \I__8520\ : Span4Mux_v
    port map (
            O => \N__40851\,
            I => \N__40848\
        );

    \I__8519\ : Odrv4
    port map (
            O => \N__40848\,
            I => \sDAC_mem_7Z0Z_3\
        );

    \I__8518\ : CascadeMux
    port map (
            O => \N__40845\,
            I => \sDAC_data_2_13_bm_1_6_cascade_\
        );

    \I__8517\ : InMux
    port map (
            O => \N__40842\,
            I => \N__40839\
        );

    \I__8516\ : LocalMux
    port map (
            O => \N__40839\,
            I => \N__40836\
        );

    \I__8515\ : Span4Mux_v
    port map (
            O => \N__40836\,
            I => \N__40833\
        );

    \I__8514\ : Odrv4
    port map (
            O => \N__40833\,
            I => \sDAC_mem_39Z0Z_3\
        );

    \I__8513\ : InMux
    port map (
            O => \N__40830\,
            I => \N__40827\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__40827\,
            I => \sDAC_mem_6Z0Z_3\
        );

    \I__8511\ : InMux
    port map (
            O => \N__40824\,
            I => \N__40821\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__40821\,
            I => \sDAC_mem_6Z0Z_4\
        );

    \I__8509\ : InMux
    port map (
            O => \N__40818\,
            I => \N__40815\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__40815\,
            I => \N__40812\
        );

    \I__8507\ : Span4Mux_v
    port map (
            O => \N__40812\,
            I => \N__40809\
        );

    \I__8506\ : Odrv4
    port map (
            O => \N__40809\,
            I => \sDAC_mem_6Z0Z_5\
        );

    \I__8505\ : InMux
    port map (
            O => \N__40806\,
            I => \N__40803\
        );

    \I__8504\ : LocalMux
    port map (
            O => \N__40803\,
            I => \N__40800\
        );

    \I__8503\ : Span4Mux_v
    port map (
            O => \N__40800\,
            I => \N__40797\
        );

    \I__8502\ : Odrv4
    port map (
            O => \N__40797\,
            I => \sDAC_mem_7Z0Z_5\
        );

    \I__8501\ : CascadeMux
    port map (
            O => \N__40794\,
            I => \sDAC_data_2_13_bm_1_8_cascade_\
        );

    \I__8500\ : InMux
    port map (
            O => \N__40791\,
            I => \N__40788\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__40788\,
            I => \N__40785\
        );

    \I__8498\ : Span4Mux_v
    port map (
            O => \N__40785\,
            I => \N__40782\
        );

    \I__8497\ : Odrv4
    port map (
            O => \N__40782\,
            I => \sDAC_mem_39Z0Z_5\
        );

    \I__8496\ : InMux
    port map (
            O => \N__40779\,
            I => \N__40776\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__40776\,
            I => \N__40773\
        );

    \I__8494\ : Span4Mux_v
    port map (
            O => \N__40773\,
            I => \N__40770\
        );

    \I__8493\ : Odrv4
    port map (
            O => \N__40770\,
            I => \sDAC_data_RNO_21Z0Z_8\
        );

    \I__8492\ : InMux
    port map (
            O => \N__40767\,
            I => \N__40764\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__40764\,
            I => \N__40761\
        );

    \I__8490\ : Odrv4
    port map (
            O => \N__40761\,
            I => \sDAC_data_RNO_20Z0Z_8\
        );

    \I__8489\ : CascadeMux
    port map (
            O => \N__40758\,
            I => \N__40755\
        );

    \I__8488\ : InMux
    port map (
            O => \N__40755\,
            I => \N__40752\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__40752\,
            I => \N__40749\
        );

    \I__8486\ : Odrv12
    port map (
            O => \N__40749\,
            I => \sDAC_data_RNO_29Z0Z_8\
        );

    \I__8485\ : InMux
    port map (
            O => \N__40746\,
            I => \N__40743\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__40743\,
            I => \N__40740\
        );

    \I__8483\ : Span4Mux_h
    port map (
            O => \N__40740\,
            I => \N__40737\
        );

    \I__8482\ : Odrv4
    port map (
            O => \N__40737\,
            I => \sDAC_data_RNO_30Z0Z_8\
        );

    \I__8481\ : CascadeMux
    port map (
            O => \N__40734\,
            I => \N__40731\
        );

    \I__8480\ : InMux
    port map (
            O => \N__40731\,
            I => \N__40728\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__40728\,
            I => \N__40725\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__40725\,
            I => \sDAC_data_2_32_ns_1_8\
        );

    \I__8477\ : InMux
    port map (
            O => \N__40722\,
            I => \N__40719\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__40719\,
            I => \N__40716\
        );

    \I__8475\ : Span4Mux_v
    port map (
            O => \N__40716\,
            I => \N__40713\
        );

    \I__8474\ : Odrv4
    port map (
            O => \N__40713\,
            I => \sDAC_mem_35Z0Z_6\
        );

    \I__8473\ : CEMux
    port map (
            O => \N__40710\,
            I => \N__40707\
        );

    \I__8472\ : LocalMux
    port map (
            O => \N__40707\,
            I => \sDAC_mem_35_1_sqmuxa\
        );

    \I__8471\ : InMux
    port map (
            O => \N__40704\,
            I => \N__40701\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__40701\,
            I => \sDAC_mem_21Z0Z_4\
        );

    \I__8469\ : InMux
    port map (
            O => \N__40698\,
            I => \N__40695\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__40695\,
            I => \sDAC_mem_21Z0Z_5\
        );

    \I__8467\ : InMux
    port map (
            O => \N__40692\,
            I => \N__40689\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__40689\,
            I => \sDAC_mem_21Z0Z_6\
        );

    \I__8465\ : InMux
    port map (
            O => \N__40686\,
            I => \N__40683\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__40683\,
            I => \N__40680\
        );

    \I__8463\ : Span4Mux_v
    port map (
            O => \N__40680\,
            I => \N__40677\
        );

    \I__8462\ : Odrv4
    port map (
            O => \N__40677\,
            I => \sDAC_mem_21Z0Z_7\
        );

    \I__8461\ : CEMux
    port map (
            O => \N__40674\,
            I => \N__40671\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__40671\,
            I => \N__40668\
        );

    \I__8459\ : Span4Mux_h
    port map (
            O => \N__40668\,
            I => \N__40665\
        );

    \I__8458\ : Span4Mux_v
    port map (
            O => \N__40665\,
            I => \N__40662\
        );

    \I__8457\ : Span4Mux_h
    port map (
            O => \N__40662\,
            I => \N__40659\
        );

    \I__8456\ : Odrv4
    port map (
            O => \N__40659\,
            I => \sDAC_mem_21_1_sqmuxa\
        );

    \I__8455\ : CEMux
    port map (
            O => \N__40656\,
            I => \N__40653\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__40653\,
            I => \N__40650\
        );

    \I__8453\ : Span4Mux_h
    port map (
            O => \N__40650\,
            I => \N__40647\
        );

    \I__8452\ : Span4Mux_h
    port map (
            O => \N__40647\,
            I => \N__40644\
        );

    \I__8451\ : Odrv4
    port map (
            O => \N__40644\,
            I => \sDAC_mem_36_1_sqmuxa\
        );

    \I__8450\ : InMux
    port map (
            O => \N__40641\,
            I => \N__40638\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__40638\,
            I => \N__40630\
        );

    \I__8448\ : InMux
    port map (
            O => \N__40637\,
            I => \N__40619\
        );

    \I__8447\ : InMux
    port map (
            O => \N__40636\,
            I => \N__40619\
        );

    \I__8446\ : InMux
    port map (
            O => \N__40635\,
            I => \N__40619\
        );

    \I__8445\ : InMux
    port map (
            O => \N__40634\,
            I => \N__40619\
        );

    \I__8444\ : InMux
    port map (
            O => \N__40633\,
            I => \N__40619\
        );

    \I__8443\ : Odrv4
    port map (
            O => \N__40630\,
            I => \N_288\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__40619\,
            I => \N_288\
        );

    \I__8441\ : CascadeMux
    port map (
            O => \N__40614\,
            I => \N__40605\
        );

    \I__8440\ : InMux
    port map (
            O => \N__40613\,
            I => \N__40600\
        );

    \I__8439\ : InMux
    port map (
            O => \N__40612\,
            I => \N__40587\
        );

    \I__8438\ : InMux
    port map (
            O => \N__40611\,
            I => \N__40587\
        );

    \I__8437\ : InMux
    port map (
            O => \N__40610\,
            I => \N__40587\
        );

    \I__8436\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40587\
        );

    \I__8435\ : InMux
    port map (
            O => \N__40608\,
            I => \N__40587\
        );

    \I__8434\ : InMux
    port map (
            O => \N__40605\,
            I => \N__40587\
        );

    \I__8433\ : CascadeMux
    port map (
            O => \N__40604\,
            I => \N__40579\
        );

    \I__8432\ : CascadeMux
    port map (
            O => \N__40603\,
            I => \N__40576\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__40600\,
            I => \N__40572\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__40587\,
            I => \N__40569\
        );

    \I__8429\ : InMux
    port map (
            O => \N__40586\,
            I => \N__40556\
        );

    \I__8428\ : InMux
    port map (
            O => \N__40585\,
            I => \N__40556\
        );

    \I__8427\ : InMux
    port map (
            O => \N__40584\,
            I => \N__40556\
        );

    \I__8426\ : InMux
    port map (
            O => \N__40583\,
            I => \N__40556\
        );

    \I__8425\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40556\
        );

    \I__8424\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40556\
        );

    \I__8423\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40552\
        );

    \I__8422\ : InMux
    port map (
            O => \N__40575\,
            I => \N__40549\
        );

    \I__8421\ : Span4Mux_v
    port map (
            O => \N__40572\,
            I => \N__40542\
        );

    \I__8420\ : Span4Mux_h
    port map (
            O => \N__40569\,
            I => \N__40542\
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__40556\,
            I => \N__40542\
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__40555\,
            I => \N__40535\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__40552\,
            I => \N__40526\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__40549\,
            I => \N__40526\
        );

    \I__8415\ : Span4Mux_v
    port map (
            O => \N__40542\,
            I => \N__40523\
        );

    \I__8414\ : InMux
    port map (
            O => \N__40541\,
            I => \N__40520\
        );

    \I__8413\ : CascadeMux
    port map (
            O => \N__40540\,
            I => \N__40513\
        );

    \I__8412\ : CascadeMux
    port map (
            O => \N__40539\,
            I => \N__40508\
        );

    \I__8411\ : CascadeMux
    port map (
            O => \N__40538\,
            I => \N__40505\
        );

    \I__8410\ : InMux
    port map (
            O => \N__40535\,
            I => \N__40502\
        );

    \I__8409\ : InMux
    port map (
            O => \N__40534\,
            I => \N__40499\
        );

    \I__8408\ : CascadeMux
    port map (
            O => \N__40533\,
            I => \N__40496\
        );

    \I__8407\ : InMux
    port map (
            O => \N__40532\,
            I => \N__40490\
        );

    \I__8406\ : InMux
    port map (
            O => \N__40531\,
            I => \N__40490\
        );

    \I__8405\ : Span4Mux_v
    port map (
            O => \N__40526\,
            I => \N__40485\
        );

    \I__8404\ : Span4Mux_h
    port map (
            O => \N__40523\,
            I => \N__40485\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__40520\,
            I => \N__40482\
        );

    \I__8402\ : InMux
    port map (
            O => \N__40519\,
            I => \N__40479\
        );

    \I__8401\ : InMux
    port map (
            O => \N__40518\,
            I => \N__40472\
        );

    \I__8400\ : InMux
    port map (
            O => \N__40517\,
            I => \N__40472\
        );

    \I__8399\ : InMux
    port map (
            O => \N__40516\,
            I => \N__40472\
        );

    \I__8398\ : InMux
    port map (
            O => \N__40513\,
            I => \N__40465\
        );

    \I__8397\ : InMux
    port map (
            O => \N__40512\,
            I => \N__40465\
        );

    \I__8396\ : InMux
    port map (
            O => \N__40511\,
            I => \N__40465\
        );

    \I__8395\ : InMux
    port map (
            O => \N__40508\,
            I => \N__40462\
        );

    \I__8394\ : InMux
    port map (
            O => \N__40505\,
            I => \N__40459\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__40502\,
            I => \N__40454\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__40499\,
            I => \N__40454\
        );

    \I__8391\ : InMux
    port map (
            O => \N__40496\,
            I => \N__40449\
        );

    \I__8390\ : InMux
    port map (
            O => \N__40495\,
            I => \N__40449\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__40490\,
            I => \N__40444\
        );

    \I__8388\ : Span4Mux_h
    port map (
            O => \N__40485\,
            I => \N__40444\
        );

    \I__8387\ : Span4Mux_h
    port map (
            O => \N__40482\,
            I => \N__40441\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__40479\,
            I => \sAddressZ0Z_3\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__40472\,
            I => \sAddressZ0Z_3\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__40465\,
            I => \sAddressZ0Z_3\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__40462\,
            I => \sAddressZ0Z_3\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__40459\,
            I => \sAddressZ0Z_3\
        );

    \I__8381\ : Odrv4
    port map (
            O => \N__40454\,
            I => \sAddressZ0Z_3\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__40449\,
            I => \sAddressZ0Z_3\
        );

    \I__8379\ : Odrv4
    port map (
            O => \N__40444\,
            I => \sAddressZ0Z_3\
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__40441\,
            I => \sAddressZ0Z_3\
        );

    \I__8377\ : CascadeMux
    port map (
            O => \N__40422\,
            I => \N_288_cascade_\
        );

    \I__8376\ : CascadeMux
    port map (
            O => \N__40419\,
            I => \N__40413\
        );

    \I__8375\ : CascadeMux
    port map (
            O => \N__40418\,
            I => \N__40409\
        );

    \I__8374\ : InMux
    port map (
            O => \N__40417\,
            I => \N__40403\
        );

    \I__8373\ : InMux
    port map (
            O => \N__40416\,
            I => \N__40392\
        );

    \I__8372\ : InMux
    port map (
            O => \N__40413\,
            I => \N__40379\
        );

    \I__8371\ : InMux
    port map (
            O => \N__40412\,
            I => \N__40379\
        );

    \I__8370\ : InMux
    port map (
            O => \N__40409\,
            I => \N__40379\
        );

    \I__8369\ : InMux
    port map (
            O => \N__40408\,
            I => \N__40379\
        );

    \I__8368\ : InMux
    port map (
            O => \N__40407\,
            I => \N__40379\
        );

    \I__8367\ : InMux
    port map (
            O => \N__40406\,
            I => \N__40379\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__40403\,
            I => \N__40376\
        );

    \I__8365\ : InMux
    port map (
            O => \N__40402\,
            I => \N__40367\
        );

    \I__8364\ : InMux
    port map (
            O => \N__40401\,
            I => \N__40367\
        );

    \I__8363\ : InMux
    port map (
            O => \N__40400\,
            I => \N__40367\
        );

    \I__8362\ : InMux
    port map (
            O => \N__40399\,
            I => \N__40367\
        );

    \I__8361\ : InMux
    port map (
            O => \N__40398\,
            I => \N__40360\
        );

    \I__8360\ : InMux
    port map (
            O => \N__40397\,
            I => \N__40360\
        );

    \I__8359\ : InMux
    port map (
            O => \N__40396\,
            I => \N__40360\
        );

    \I__8358\ : InMux
    port map (
            O => \N__40395\,
            I => \N__40356\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__40392\,
            I => \N__40352\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__40379\,
            I => \N__40349\
        );

    \I__8355\ : Span4Mux_v
    port map (
            O => \N__40376\,
            I => \N__40340\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__40367\,
            I => \N__40340\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__40360\,
            I => \N__40340\
        );

    \I__8352\ : InMux
    port map (
            O => \N__40359\,
            I => \N__40337\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__40356\,
            I => \N__40330\
        );

    \I__8350\ : CascadeMux
    port map (
            O => \N__40355\,
            I => \N__40320\
        );

    \I__8349\ : Span4Mux_v
    port map (
            O => \N__40352\,
            I => \N__40315\
        );

    \I__8348\ : Span4Mux_v
    port map (
            O => \N__40349\,
            I => \N__40315\
        );

    \I__8347\ : InMux
    port map (
            O => \N__40348\,
            I => \N__40310\
        );

    \I__8346\ : InMux
    port map (
            O => \N__40347\,
            I => \N__40310\
        );

    \I__8345\ : Span4Mux_h
    port map (
            O => \N__40340\,
            I => \N__40307\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__40337\,
            I => \N__40301\
        );

    \I__8343\ : InMux
    port map (
            O => \N__40336\,
            I => \N__40296\
        );

    \I__8342\ : InMux
    port map (
            O => \N__40335\,
            I => \N__40296\
        );

    \I__8341\ : InMux
    port map (
            O => \N__40334\,
            I => \N__40291\
        );

    \I__8340\ : InMux
    port map (
            O => \N__40333\,
            I => \N__40291\
        );

    \I__8339\ : Span4Mux_h
    port map (
            O => \N__40330\,
            I => \N__40288\
        );

    \I__8338\ : InMux
    port map (
            O => \N__40329\,
            I => \N__40283\
        );

    \I__8337\ : InMux
    port map (
            O => \N__40328\,
            I => \N__40283\
        );

    \I__8336\ : InMux
    port map (
            O => \N__40327\,
            I => \N__40278\
        );

    \I__8335\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40278\
        );

    \I__8334\ : InMux
    port map (
            O => \N__40325\,
            I => \N__40269\
        );

    \I__8333\ : InMux
    port map (
            O => \N__40324\,
            I => \N__40269\
        );

    \I__8332\ : InMux
    port map (
            O => \N__40323\,
            I => \N__40269\
        );

    \I__8331\ : InMux
    port map (
            O => \N__40320\,
            I => \N__40269\
        );

    \I__8330\ : Span4Mux_h
    port map (
            O => \N__40315\,
            I => \N__40264\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__40310\,
            I => \N__40264\
        );

    \I__8328\ : Span4Mux_v
    port map (
            O => \N__40307\,
            I => \N__40261\
        );

    \I__8327\ : InMux
    port map (
            O => \N__40306\,
            I => \N__40254\
        );

    \I__8326\ : InMux
    port map (
            O => \N__40305\,
            I => \N__40254\
        );

    \I__8325\ : InMux
    port map (
            O => \N__40304\,
            I => \N__40254\
        );

    \I__8324\ : Span12Mux_h
    port map (
            O => \N__40301\,
            I => \N__40251\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__40296\,
            I => \sAddressZ0Z_0\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__40291\,
            I => \sAddressZ0Z_0\
        );

    \I__8321\ : Odrv4
    port map (
            O => \N__40288\,
            I => \sAddressZ0Z_0\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__40283\,
            I => \sAddressZ0Z_0\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__40278\,
            I => \sAddressZ0Z_0\
        );

    \I__8318\ : LocalMux
    port map (
            O => \N__40269\,
            I => \sAddressZ0Z_0\
        );

    \I__8317\ : Odrv4
    port map (
            O => \N__40264\,
            I => \sAddressZ0Z_0\
        );

    \I__8316\ : Odrv4
    port map (
            O => \N__40261\,
            I => \sAddressZ0Z_0\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__40254\,
            I => \sAddressZ0Z_0\
        );

    \I__8314\ : Odrv12
    port map (
            O => \N__40251\,
            I => \sAddressZ0Z_0\
        );

    \I__8313\ : InMux
    port map (
            O => \N__40230\,
            I => \N__40227\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__40227\,
            I => \N__40224\
        );

    \I__8311\ : Odrv12
    port map (
            O => \N__40224\,
            I => \sDAC_mem_35Z0Z_0\
        );

    \I__8310\ : InMux
    port map (
            O => \N__40221\,
            I => \N__40218\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__40218\,
            I => \N__40215\
        );

    \I__8308\ : Span4Mux_v
    port map (
            O => \N__40215\,
            I => \N__40212\
        );

    \I__8307\ : Odrv4
    port map (
            O => \N__40212\,
            I => \sDAC_mem_35Z0Z_2\
        );

    \I__8306\ : InMux
    port map (
            O => \N__40209\,
            I => \N__40206\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__40206\,
            I => \N__40203\
        );

    \I__8304\ : Span4Mux_v
    port map (
            O => \N__40203\,
            I => \N__40200\
        );

    \I__8303\ : Span4Mux_h
    port map (
            O => \N__40200\,
            I => \N__40197\
        );

    \I__8302\ : Odrv4
    port map (
            O => \N__40197\,
            I => \sDAC_mem_35Z0Z_4\
        );

    \I__8301\ : InMux
    port map (
            O => \N__40194\,
            I => \N__40191\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__40191\,
            I => \N__40188\
        );

    \I__8299\ : Span4Mux_v
    port map (
            O => \N__40188\,
            I => \N__40185\
        );

    \I__8298\ : Odrv4
    port map (
            O => \N__40185\,
            I => \sDAC_mem_35Z0Z_5\
        );

    \I__8297\ : InMux
    port map (
            O => \N__40182\,
            I => \N__40179\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__40179\,
            I => \N__40176\
        );

    \I__8295\ : Odrv4
    port map (
            O => \N__40176\,
            I => \sDAC_mem_39Z0Z_2\
        );

    \I__8294\ : InMux
    port map (
            O => \N__40173\,
            I => \N__40170\
        );

    \I__8293\ : LocalMux
    port map (
            O => \N__40170\,
            I => \N__40167\
        );

    \I__8292\ : Span4Mux_v
    port map (
            O => \N__40167\,
            I => \N__40164\
        );

    \I__8291\ : Odrv4
    port map (
            O => \N__40164\,
            I => \sDAC_mem_39Z0Z_4\
        );

    \I__8290\ : InMux
    port map (
            O => \N__40161\,
            I => \N__40158\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__40158\,
            I => \N__40155\
        );

    \I__8288\ : Span4Mux_v
    port map (
            O => \N__40155\,
            I => \N__40152\
        );

    \I__8287\ : Odrv4
    port map (
            O => \N__40152\,
            I => \sDAC_mem_39Z0Z_7\
        );

    \I__8286\ : CEMux
    port map (
            O => \N__40149\,
            I => \N__40146\
        );

    \I__8285\ : LocalMux
    port map (
            O => \N__40146\,
            I => \N__40143\
        );

    \I__8284\ : Odrv4
    port map (
            O => \N__40143\,
            I => \sDAC_mem_37_1_sqmuxa\
        );

    \I__8283\ : CEMux
    port map (
            O => \N__40140\,
            I => \N__40137\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__40137\,
            I => \sDAC_mem_39_1_sqmuxa\
        );

    \I__8281\ : InMux
    port map (
            O => \N__40134\,
            I => \N__40131\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__40131\,
            I => \sDAC_mem_25Z0Z_2\
        );

    \I__8279\ : InMux
    port map (
            O => \N__40128\,
            I => \N__40125\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__40125\,
            I => \N__40122\
        );

    \I__8277\ : Span4Mux_v
    port map (
            O => \N__40122\,
            I => \N__40119\
        );

    \I__8276\ : Span4Mux_v
    port map (
            O => \N__40119\,
            I => \N__40116\
        );

    \I__8275\ : Odrv4
    port map (
            O => \N__40116\,
            I => \sDAC_mem_25Z0Z_5\
        );

    \I__8274\ : InMux
    port map (
            O => \N__40113\,
            I => \N__40110\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__40110\,
            I => \sDAC_mem_25Z0Z_0\
        );

    \I__8272\ : InMux
    port map (
            O => \N__40107\,
            I => \N__40104\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__40104\,
            I => \N__40101\
        );

    \I__8270\ : Odrv4
    port map (
            O => \N__40101\,
            I => \sDAC_mem_25Z0Z_6\
        );

    \I__8269\ : InMux
    port map (
            O => \N__40098\,
            I => \N__40095\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__40095\,
            I => \N__40092\
        );

    \I__8267\ : Odrv4
    port map (
            O => \N__40092\,
            I => \sDAC_mem_25Z0Z_3\
        );

    \I__8266\ : CEMux
    port map (
            O => \N__40089\,
            I => \N__40085\
        );

    \I__8265\ : CEMux
    port map (
            O => \N__40088\,
            I => \N__40082\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__40085\,
            I => \N__40079\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__40082\,
            I => \N__40076\
        );

    \I__8262\ : Span4Mux_v
    port map (
            O => \N__40079\,
            I => \N__40073\
        );

    \I__8261\ : Odrv12
    port map (
            O => \N__40076\,
            I => \sDAC_mem_34_1_sqmuxa\
        );

    \I__8260\ : Odrv4
    port map (
            O => \N__40073\,
            I => \sDAC_mem_34_1_sqmuxa\
        );

    \I__8259\ : InMux
    port map (
            O => \N__40068\,
            I => \N__40065\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__40065\,
            I => \N__40062\
        );

    \I__8257\ : Odrv12
    port map (
            O => \N__40062\,
            I => \sDAC_mem_39Z0Z_0\
        );

    \I__8256\ : InMux
    port map (
            O => \N__40059\,
            I => \N__40056\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__40056\,
            I => \N__40053\
        );

    \I__8254\ : Span4Mux_h
    port map (
            O => \N__40053\,
            I => \N__40050\
        );

    \I__8253\ : Odrv4
    port map (
            O => \N__40050\,
            I => \sDAC_mem_39Z0Z_1\
        );

    \I__8252\ : CascadeMux
    port map (
            O => \N__40047\,
            I => \sDAC_data_2_39_ns_1_10_cascade_\
        );

    \I__8251\ : CascadeMux
    port map (
            O => \N__40044\,
            I => \N__40041\
        );

    \I__8250\ : InMux
    port map (
            O => \N__40041\,
            I => \N__40038\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__40038\,
            I => \N__40035\
        );

    \I__8248\ : Odrv12
    port map (
            O => \N__40035\,
            I => \sDAC_data_RNO_11Z0Z_10\
        );

    \I__8247\ : InMux
    port map (
            O => \N__40032\,
            I => \N__40029\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__40029\,
            I => \N__40026\
        );

    \I__8245\ : Odrv4
    port map (
            O => \N__40026\,
            I => \sDAC_mem_26Z0Z_7\
        );

    \I__8244\ : InMux
    port map (
            O => \N__40023\,
            I => \N__40020\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__40020\,
            I => \sDAC_data_RNO_32Z0Z_10\
        );

    \I__8242\ : InMux
    port map (
            O => \N__40017\,
            I => \N__40014\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__40014\,
            I => \sDAC_mem_29Z0Z_7\
        );

    \I__8240\ : InMux
    port map (
            O => \N__40011\,
            I => \N__40008\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__40008\,
            I => \sDAC_data_RNO_23Z0Z_10\
        );

    \I__8238\ : InMux
    port map (
            O => \N__40005\,
            I => \N__40002\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__40002\,
            I => \N__39999\
        );

    \I__8236\ : Span4Mux_v
    port map (
            O => \N__39999\,
            I => \N__39996\
        );

    \I__8235\ : Odrv4
    port map (
            O => \N__39996\,
            I => \sDAC_mem_31Z0Z_7\
        );

    \I__8234\ : InMux
    port map (
            O => \N__39993\,
            I => \N__39990\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__39990\,
            I => \N__39987\
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__39987\,
            I => \sDAC_mem_30Z0Z_7\
        );

    \I__8231\ : InMux
    port map (
            O => \N__39984\,
            I => \N__39981\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__39981\,
            I => \sDAC_data_RNO_24Z0Z_10\
        );

    \I__8229\ : InMux
    port map (
            O => \N__39978\,
            I => \N__39975\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__39975\,
            I => \sDAC_mem_24Z0Z_7\
        );

    \I__8227\ : CEMux
    port map (
            O => \N__39972\,
            I => \N__39968\
        );

    \I__8226\ : CEMux
    port map (
            O => \N__39971\,
            I => \N__39964\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__39968\,
            I => \N__39961\
        );

    \I__8224\ : CEMux
    port map (
            O => \N__39967\,
            I => \N__39958\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__39964\,
            I => \N__39955\
        );

    \I__8222\ : Span4Mux_h
    port map (
            O => \N__39961\,
            I => \N__39951\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__39958\,
            I => \N__39948\
        );

    \I__8220\ : Span4Mux_h
    port map (
            O => \N__39955\,
            I => \N__39945\
        );

    \I__8219\ : CEMux
    port map (
            O => \N__39954\,
            I => \N__39942\
        );

    \I__8218\ : Span4Mux_h
    port map (
            O => \N__39951\,
            I => \N__39939\
        );

    \I__8217\ : Span4Mux_h
    port map (
            O => \N__39948\,
            I => \N__39932\
        );

    \I__8216\ : Span4Mux_h
    port map (
            O => \N__39945\,
            I => \N__39932\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__39942\,
            I => \N__39932\
        );

    \I__8214\ : Span4Mux_v
    port map (
            O => \N__39939\,
            I => \N__39929\
        );

    \I__8213\ : Span4Mux_v
    port map (
            O => \N__39932\,
            I => \N__39926\
        );

    \I__8212\ : Odrv4
    port map (
            O => \N__39929\,
            I => \sDAC_mem_24_1_sqmuxa\
        );

    \I__8211\ : Odrv4
    port map (
            O => \N__39926\,
            I => \sDAC_mem_24_1_sqmuxa\
        );

    \I__8210\ : CascadeMux
    port map (
            O => \N__39921\,
            I => \N__39918\
        );

    \I__8209\ : InMux
    port map (
            O => \N__39918\,
            I => \N__39915\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__39915\,
            I => \N__39912\
        );

    \I__8207\ : Span4Mux_h
    port map (
            O => \N__39912\,
            I => \N__39909\
        );

    \I__8206\ : Odrv4
    port map (
            O => \N__39909\,
            I => \sDAC_data_RNO_32Z0Z_3\
        );

    \I__8205\ : InMux
    port map (
            O => \N__39906\,
            I => \N__39903\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__39903\,
            I => \N__39900\
        );

    \I__8203\ : Odrv4
    port map (
            O => \N__39900\,
            I => \sDAC_data_RNO_31Z0Z_3\
        );

    \I__8202\ : InMux
    port map (
            O => \N__39897\,
            I => \N__39894\
        );

    \I__8201\ : LocalMux
    port map (
            O => \N__39894\,
            I => \sDAC_mem_25Z0Z_4\
        );

    \I__8200\ : InMux
    port map (
            O => \N__39891\,
            I => \N__39888\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__39888\,
            I => \sDAC_mem_25Z0Z_7\
        );

    \I__8198\ : InMux
    port map (
            O => \N__39885\,
            I => \N__39882\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__39882\,
            I => \N__39879\
        );

    \I__8196\ : Span4Mux_v
    port map (
            O => \N__39879\,
            I => \N__39876\
        );

    \I__8195\ : Span4Mux_h
    port map (
            O => \N__39876\,
            I => \N__39873\
        );

    \I__8194\ : Span4Mux_v
    port map (
            O => \N__39873\,
            I => \N__39870\
        );

    \I__8193\ : Odrv4
    port map (
            O => \N__39870\,
            I => \sDAC_mem_23Z0Z_5\
        );

    \I__8192\ : InMux
    port map (
            O => \N__39867\,
            I => \N__39864\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__39864\,
            I => \sDAC_mem_22Z0Z_5\
        );

    \I__8190\ : InMux
    port map (
            O => \N__39861\,
            I => \N__39858\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__39858\,
            I => \N__39855\
        );

    \I__8188\ : Span4Mux_v
    port map (
            O => \N__39855\,
            I => \N__39852\
        );

    \I__8187\ : Span4Mux_h
    port map (
            O => \N__39852\,
            I => \N__39849\
        );

    \I__8186\ : Span4Mux_v
    port map (
            O => \N__39849\,
            I => \N__39846\
        );

    \I__8185\ : Odrv4
    port map (
            O => \N__39846\,
            I => \sDAC_mem_23Z0Z_6\
        );

    \I__8184\ : InMux
    port map (
            O => \N__39843\,
            I => \N__39840\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__39840\,
            I => \N__39837\
        );

    \I__8182\ : Span4Mux_v
    port map (
            O => \N__39837\,
            I => \N__39834\
        );

    \I__8181\ : Odrv4
    port map (
            O => \N__39834\,
            I => \sDAC_data_RNO_21Z0Z_9\
        );

    \I__8180\ : InMux
    port map (
            O => \N__39831\,
            I => \N__39828\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__39828\,
            I => \sDAC_mem_22Z0Z_6\
        );

    \I__8178\ : CEMux
    port map (
            O => \N__39825\,
            I => \N__39821\
        );

    \I__8177\ : CEMux
    port map (
            O => \N__39824\,
            I => \N__39818\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__39821\,
            I => \N__39814\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__39818\,
            I => \N__39811\
        );

    \I__8174\ : CEMux
    port map (
            O => \N__39817\,
            I => \N__39808\
        );

    \I__8173\ : Span4Mux_v
    port map (
            O => \N__39814\,
            I => \N__39805\
        );

    \I__8172\ : Span4Mux_v
    port map (
            O => \N__39811\,
            I => \N__39802\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__39808\,
            I => \N__39799\
        );

    \I__8170\ : Span4Mux_h
    port map (
            O => \N__39805\,
            I => \N__39794\
        );

    \I__8169\ : Span4Mux_h
    port map (
            O => \N__39802\,
            I => \N__39794\
        );

    \I__8168\ : Span4Mux_h
    port map (
            O => \N__39799\,
            I => \N__39791\
        );

    \I__8167\ : Odrv4
    port map (
            O => \N__39794\,
            I => \sDAC_mem_22_1_sqmuxa\
        );

    \I__8166\ : Odrv4
    port map (
            O => \N__39791\,
            I => \sDAC_mem_22_1_sqmuxa\
        );

    \I__8165\ : InMux
    port map (
            O => \N__39786\,
            I => \N__39783\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__39783\,
            I => \sDAC_mem_29Z0Z_1\
        );

    \I__8163\ : InMux
    port map (
            O => \N__39780\,
            I => \N__39777\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__39777\,
            I => \sDAC_mem_30Z0Z_1\
        );

    \I__8161\ : InMux
    port map (
            O => \N__39774\,
            I => \N__39771\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__39771\,
            I => \N__39768\
        );

    \I__8159\ : Span4Mux_h
    port map (
            O => \N__39768\,
            I => \N__39765\
        );

    \I__8158\ : Odrv4
    port map (
            O => \N__39765\,
            I => \sDAC_mem_31Z0Z_1\
        );

    \I__8157\ : InMux
    port map (
            O => \N__39762\,
            I => \N__39759\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__39759\,
            I => \N__39756\
        );

    \I__8155\ : Span4Mux_h
    port map (
            O => \N__39756\,
            I => \N__39753\
        );

    \I__8154\ : Odrv4
    port map (
            O => \N__39753\,
            I => \sDAC_mem_31Z0Z_4\
        );

    \I__8153\ : InMux
    port map (
            O => \N__39750\,
            I => \N__39747\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__39747\,
            I => \sDAC_mem_30Z0Z_4\
        );

    \I__8151\ : InMux
    port map (
            O => \N__39744\,
            I => \N__39741\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__39741\,
            I => \N__39738\
        );

    \I__8149\ : Odrv4
    port map (
            O => \N__39738\,
            I => \sDAC_data_RNO_24Z0Z_7\
        );

    \I__8148\ : CascadeMux
    port map (
            O => \N__39735\,
            I => \sDAC_data_RNO_31Z0Z_10_cascade_\
        );

    \I__8147\ : CascadeMux
    port map (
            O => \N__39732\,
            I => \N_142_cascade_\
        );

    \I__8146\ : InMux
    port map (
            O => \N__39729\,
            I => \N__39726\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__39726\,
            I => \N__39723\
        );

    \I__8144\ : Odrv4
    port map (
            O => \N__39723\,
            I => \sDAC_mem_30Z0Z_2\
        );

    \I__8143\ : InMux
    port map (
            O => \N__39720\,
            I => \N__39717\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__39717\,
            I => \N__39714\
        );

    \I__8141\ : Span4Mux_v
    port map (
            O => \N__39714\,
            I => \N__39711\
        );

    \I__8140\ : Odrv4
    port map (
            O => \N__39711\,
            I => \sDAC_mem_30Z0Z_3\
        );

    \I__8139\ : InMux
    port map (
            O => \N__39708\,
            I => \N__39705\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__39705\,
            I => \N__39702\
        );

    \I__8137\ : Odrv4
    port map (
            O => \N__39702\,
            I => \sDAC_mem_30Z0Z_5\
        );

    \I__8136\ : InMux
    port map (
            O => \N__39699\,
            I => \N__39696\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__39696\,
            I => \sDAC_mem_30Z0Z_6\
        );

    \I__8134\ : CEMux
    port map (
            O => \N__39693\,
            I => \N__39690\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__39690\,
            I => \sDAC_mem_30_1_sqmuxa\
        );

    \I__8132\ : InMux
    port map (
            O => \N__39687\,
            I => \N__39684\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__39684\,
            I => \N__39681\
        );

    \I__8130\ : Span12Mux_v
    port map (
            O => \N__39681\,
            I => \N__39678\
        );

    \I__8129\ : Odrv12
    port map (
            O => \N__39678\,
            I => \sDAC_mem_36Z0Z_0\
        );

    \I__8128\ : InMux
    port map (
            O => \N__39675\,
            I => \N__39672\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__39672\,
            I => \N__39669\
        );

    \I__8126\ : Span4Mux_v
    port map (
            O => \N__39669\,
            I => \N__39666\
        );

    \I__8125\ : Span4Mux_v
    port map (
            O => \N__39666\,
            I => \N__39663\
        );

    \I__8124\ : Odrv4
    port map (
            O => \N__39663\,
            I => \sDAC_mem_37Z0Z_0\
        );

    \I__8123\ : CascadeMux
    port map (
            O => \N__39660\,
            I => \sDAC_data_2_13_am_1_3_cascade_\
        );

    \I__8122\ : InMux
    port map (
            O => \N__39657\,
            I => \N__39654\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__39654\,
            I => \N__39651\
        );

    \I__8120\ : Span12Mux_h
    port map (
            O => \N__39651\,
            I => \N__39648\
        );

    \I__8119\ : Odrv12
    port map (
            O => \N__39648\,
            I => \sDAC_mem_5Z0Z_0\
        );

    \I__8118\ : InMux
    port map (
            O => \N__39645\,
            I => \N__39642\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__39642\,
            I => \sDAC_mem_4Z0Z_0\
        );

    \I__8116\ : CEMux
    port map (
            O => \N__39639\,
            I => \N__39636\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__39636\,
            I => \N__39632\
        );

    \I__8114\ : CEMux
    port map (
            O => \N__39635\,
            I => \N__39628\
        );

    \I__8113\ : Span4Mux_v
    port map (
            O => \N__39632\,
            I => \N__39624\
        );

    \I__8112\ : CEMux
    port map (
            O => \N__39631\,
            I => \N__39621\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__39628\,
            I => \N__39618\
        );

    \I__8110\ : CEMux
    port map (
            O => \N__39627\,
            I => \N__39615\
        );

    \I__8109\ : Span4Mux_h
    port map (
            O => \N__39624\,
            I => \N__39610\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__39621\,
            I => \N__39610\
        );

    \I__8107\ : Span4Mux_h
    port map (
            O => \N__39618\,
            I => \N__39607\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__39615\,
            I => \N__39604\
        );

    \I__8105\ : Odrv4
    port map (
            O => \N__39610\,
            I => \sDAC_mem_4_1_sqmuxa\
        );

    \I__8104\ : Odrv4
    port map (
            O => \N__39607\,
            I => \sDAC_mem_4_1_sqmuxa\
        );

    \I__8103\ : Odrv4
    port map (
            O => \N__39604\,
            I => \sDAC_mem_4_1_sqmuxa\
        );

    \I__8102\ : InMux
    port map (
            O => \N__39597\,
            I => \N__39594\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__39594\,
            I => \N__39591\
        );

    \I__8100\ : Odrv12
    port map (
            O => \N__39591\,
            I => \sDAC_mem_36Z0Z_1\
        );

    \I__8099\ : InMux
    port map (
            O => \N__39588\,
            I => \N__39585\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__39585\,
            I => \N__39582\
        );

    \I__8097\ : Span4Mux_v
    port map (
            O => \N__39582\,
            I => \N__39579\
        );

    \I__8096\ : Span4Mux_h
    port map (
            O => \N__39579\,
            I => \N__39576\
        );

    \I__8095\ : Span4Mux_v
    port map (
            O => \N__39576\,
            I => \N__39573\
        );

    \I__8094\ : Odrv4
    port map (
            O => \N__39573\,
            I => \sDAC_mem_4Z0Z_1\
        );

    \I__8093\ : InMux
    port map (
            O => \N__39570\,
            I => \N__39567\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__39567\,
            I => \N__39564\
        );

    \I__8091\ : Span4Mux_v
    port map (
            O => \N__39564\,
            I => \N__39561\
        );

    \I__8090\ : Span4Mux_v
    port map (
            O => \N__39561\,
            I => \N__39558\
        );

    \I__8089\ : Odrv4
    port map (
            O => \N__39558\,
            I => \sDAC_mem_37Z0Z_1\
        );

    \I__8088\ : CascadeMux
    port map (
            O => \N__39555\,
            I => \sDAC_data_2_13_am_1_4_cascade_\
        );

    \I__8087\ : InMux
    port map (
            O => \N__39552\,
            I => \N__39549\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__39549\,
            I => \N__39546\
        );

    \I__8085\ : Span4Mux_v
    port map (
            O => \N__39546\,
            I => \N__39543\
        );

    \I__8084\ : Span4Mux_v
    port map (
            O => \N__39543\,
            I => \N__39540\
        );

    \I__8083\ : Odrv4
    port map (
            O => \N__39540\,
            I => \sDAC_mem_5Z0Z_1\
        );

    \I__8082\ : InMux
    port map (
            O => \N__39537\,
            I => \N__39534\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__39534\,
            I => \N__39531\
        );

    \I__8080\ : Odrv4
    port map (
            O => \N__39531\,
            I => \sDAC_data_RNO_20Z0Z_10\
        );

    \I__8079\ : CEMux
    port map (
            O => \N__39528\,
            I => \N__39525\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__39525\,
            I => \N__39522\
        );

    \I__8077\ : Span4Mux_h
    port map (
            O => \N__39522\,
            I => \N__39519\
        );

    \I__8076\ : Span4Mux_h
    port map (
            O => \N__39519\,
            I => \N__39516\
        );

    \I__8075\ : Odrv4
    port map (
            O => \N__39516\,
            I => \sDAC_mem_26_1_sqmuxa\
        );

    \I__8074\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39510\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__39510\,
            I => \N__39507\
        );

    \I__8072\ : Odrv4
    port map (
            O => \N__39507\,
            I => \sDAC_data_RNO_14Z0Z_10\
        );

    \I__8071\ : InMux
    port map (
            O => \N__39504\,
            I => \N__39501\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__39501\,
            I => \N__39498\
        );

    \I__8069\ : Odrv4
    port map (
            O => \N__39498\,
            I => \sDAC_data_RNO_5Z0Z_10\
        );

    \I__8068\ : CascadeMux
    port map (
            O => \N__39495\,
            I => \sDAC_data_2_14_ns_1_10_cascade_\
        );

    \I__8067\ : InMux
    port map (
            O => \N__39492\,
            I => \N__39489\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__39489\,
            I => \sDAC_data_RNO_10Z0Z_10\
        );

    \I__8065\ : InMux
    port map (
            O => \N__39486\,
            I => \N__39483\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__39483\,
            I => \sDAC_data_RNO_2Z0Z_10\
        );

    \I__8063\ : CascadeMux
    port map (
            O => \N__39480\,
            I => \sDAC_data_2_41_ns_1_10_cascade_\
        );

    \I__8062\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39474\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__39474\,
            I => \sDAC_data_RNO_1Z0Z_10\
        );

    \I__8060\ : CascadeMux
    port map (
            O => \N__39471\,
            I => \sDAC_data_2_10_cascade_\
        );

    \I__8059\ : InMux
    port map (
            O => \N__39468\,
            I => \N__39465\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__39465\,
            I => \N__39462\
        );

    \I__8057\ : Span4Mux_v
    port map (
            O => \N__39462\,
            I => \N__39459\
        );

    \I__8056\ : Span4Mux_h
    port map (
            O => \N__39459\,
            I => \N__39456\
        );

    \I__8055\ : Sp12to4
    port map (
            O => \N__39456\,
            I => \N__39453\
        );

    \I__8054\ : Odrv12
    port map (
            O => \N__39453\,
            I => \sDAC_dataZ0Z_10\
        );

    \I__8053\ : InMux
    port map (
            O => \N__39450\,
            I => \N__39447\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__39447\,
            I => \N__39444\
        );

    \I__8051\ : Span12Mux_v
    port map (
            O => \N__39444\,
            I => \N__39441\
        );

    \I__8050\ : Odrv12
    port map (
            O => \N__39441\,
            I => \sDAC_mem_36Z0Z_7\
        );

    \I__8049\ : InMux
    port map (
            O => \N__39438\,
            I => \N__39435\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__39435\,
            I => \N__39432\
        );

    \I__8047\ : Sp12to4
    port map (
            O => \N__39432\,
            I => \N__39429\
        );

    \I__8046\ : Odrv12
    port map (
            O => \N__39429\,
            I => \sDAC_mem_37Z0Z_7\
        );

    \I__8045\ : CascadeMux
    port map (
            O => \N__39426\,
            I => \sDAC_data_2_13_am_1_10_cascade_\
        );

    \I__8044\ : InMux
    port map (
            O => \N__39423\,
            I => \N__39420\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__39420\,
            I => \N__39417\
        );

    \I__8042\ : Span12Mux_v
    port map (
            O => \N__39417\,
            I => \N__39414\
        );

    \I__8041\ : Odrv12
    port map (
            O => \N__39414\,
            I => \sDAC_mem_5Z0Z_7\
        );

    \I__8040\ : InMux
    port map (
            O => \N__39411\,
            I => \N__39408\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__39408\,
            I => \sDAC_data_RNO_4Z0Z_10\
        );

    \I__8038\ : InMux
    port map (
            O => \N__39405\,
            I => \N__39402\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__39402\,
            I => \sDAC_mem_4Z0Z_7\
        );

    \I__8036\ : CascadeMux
    port map (
            O => \N__39399\,
            I => \N__39396\
        );

    \I__8035\ : InMux
    port map (
            O => \N__39396\,
            I => \N__39393\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__39393\,
            I => \N__39390\
        );

    \I__8033\ : Span12Mux_h
    port map (
            O => \N__39390\,
            I => \N__39387\
        );

    \I__8032\ : Odrv12
    port map (
            O => \N__39387\,
            I => \sDAC_mem_2Z0Z_5\
        );

    \I__8031\ : InMux
    port map (
            O => \N__39384\,
            I => \N__39381\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__39381\,
            I => \N__39378\
        );

    \I__8029\ : Span4Mux_v
    port map (
            O => \N__39378\,
            I => \N__39375\
        );

    \I__8028\ : Span4Mux_v
    port map (
            O => \N__39375\,
            I => \N__39372\
        );

    \I__8027\ : Odrv4
    port map (
            O => \N__39372\,
            I => \sDAC_mem_34Z0Z_5\
        );

    \I__8026\ : CascadeMux
    port map (
            O => \N__39369\,
            I => \sDAC_data_2_6_bm_1_8_cascade_\
        );

    \I__8025\ : InMux
    port map (
            O => \N__39366\,
            I => \N__39363\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__39363\,
            I => \sDAC_mem_3Z0Z_5\
        );

    \I__8023\ : InMux
    port map (
            O => \N__39360\,
            I => \N__39357\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__39357\,
            I => \N__39354\
        );

    \I__8021\ : Span4Mux_h
    port map (
            O => \N__39354\,
            I => \N__39351\
        );

    \I__8020\ : Span4Mux_h
    port map (
            O => \N__39351\,
            I => \N__39348\
        );

    \I__8019\ : Odrv4
    port map (
            O => \N__39348\,
            I => \sDAC_mem_33Z0Z_7\
        );

    \I__8018\ : CascadeMux
    port map (
            O => \N__39345\,
            I => \sDAC_data_RNO_26Z0Z_10_cascade_\
        );

    \I__8017\ : CascadeMux
    port map (
            O => \N__39342\,
            I => \N__39338\
        );

    \I__8016\ : CascadeMux
    port map (
            O => \N__39341\,
            I => \N__39335\
        );

    \I__8015\ : InMux
    port map (
            O => \N__39338\,
            I => \N__39330\
        );

    \I__8014\ : InMux
    port map (
            O => \N__39335\,
            I => \N__39330\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__39330\,
            I => \N__39327\
        );

    \I__8012\ : Span4Mux_v
    port map (
            O => \N__39327\,
            I => \N__39324\
        );

    \I__8011\ : Odrv4
    port map (
            O => \N__39324\,
            I => \sDAC_mem_1Z0Z_7\
        );

    \I__8010\ : InMux
    port map (
            O => \N__39321\,
            I => \N__39315\
        );

    \I__8009\ : InMux
    port map (
            O => \N__39320\,
            I => \N__39315\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__39315\,
            I => \N__39312\
        );

    \I__8007\ : Span4Mux_h
    port map (
            O => \N__39312\,
            I => \N__39309\
        );

    \I__8006\ : Odrv4
    port map (
            O => \N__39309\,
            I => \sDAC_mem_32Z0Z_7\
        );

    \I__8005\ : InMux
    port map (
            O => \N__39306\,
            I => \N__39303\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__39303\,
            I => \sDAC_data_RNO_27Z0Z_10\
        );

    \I__8003\ : CascadeMux
    port map (
            O => \N__39300\,
            I => \N__39297\
        );

    \I__8002\ : InMux
    port map (
            O => \N__39297\,
            I => \N__39293\
        );

    \I__8001\ : CascadeMux
    port map (
            O => \N__39296\,
            I => \N__39290\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__39293\,
            I => \N__39287\
        );

    \I__7999\ : InMux
    port map (
            O => \N__39290\,
            I => \N__39284\
        );

    \I__7998\ : Span4Mux_h
    port map (
            O => \N__39287\,
            I => \N__39279\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__39284\,
            I => \N__39279\
        );

    \I__7996\ : Span4Mux_h
    port map (
            O => \N__39279\,
            I => \N__39276\
        );

    \I__7995\ : Span4Mux_h
    port map (
            O => \N__39276\,
            I => \N__39273\
        );

    \I__7994\ : Odrv4
    port map (
            O => \N__39273\,
            I => \sDAC_mem_1Z0Z_0\
        );

    \I__7993\ : InMux
    port map (
            O => \N__39270\,
            I => \N__39267\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__39267\,
            I => \N__39264\
        );

    \I__7991\ : Span4Mux_h
    port map (
            O => \N__39264\,
            I => \N__39260\
        );

    \I__7990\ : InMux
    port map (
            O => \N__39263\,
            I => \N__39257\
        );

    \I__7989\ : Odrv4
    port map (
            O => \N__39260\,
            I => \sDAC_mem_32Z0Z_0\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__39257\,
            I => \sDAC_mem_32Z0Z_0\
        );

    \I__7987\ : InMux
    port map (
            O => \N__39252\,
            I => \N__39249\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__39249\,
            I => \N__39246\
        );

    \I__7985\ : Span4Mux_v
    port map (
            O => \N__39246\,
            I => \N__39243\
        );

    \I__7984\ : Span4Mux_h
    port map (
            O => \N__39243\,
            I => \N__39240\
        );

    \I__7983\ : Odrv4
    port map (
            O => \N__39240\,
            I => \sDAC_mem_33Z0Z_0\
        );

    \I__7982\ : CascadeMux
    port map (
            O => \N__39237\,
            I => \sDAC_data_RNO_26Z0Z_3_cascade_\
        );

    \I__7981\ : InMux
    port map (
            O => \N__39234\,
            I => \N__39231\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__39231\,
            I => \N__39228\
        );

    \I__7979\ : Odrv4
    port map (
            O => \N__39228\,
            I => \sDAC_data_RNO_27Z0Z_3\
        );

    \I__7978\ : InMux
    port map (
            O => \N__39225\,
            I => \N__39222\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__39222\,
            I => \N__39219\
        );

    \I__7976\ : Span4Mux_v
    port map (
            O => \N__39219\,
            I => \N__39216\
        );

    \I__7975\ : Odrv4
    port map (
            O => \N__39216\,
            I => \sDAC_data_RNO_21Z0Z_10\
        );

    \I__7974\ : CascadeMux
    port map (
            O => \N__39213\,
            I => \N__39210\
        );

    \I__7973\ : InMux
    port map (
            O => \N__39210\,
            I => \N__39207\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__39207\,
            I => \N__39204\
        );

    \I__7971\ : Odrv12
    port map (
            O => \N__39204\,
            I => \sDAC_data_RNO_30Z0Z_10\
        );

    \I__7970\ : InMux
    port map (
            O => \N__39201\,
            I => \N__39198\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__39198\,
            I => \sDAC_data_2_32_ns_1_10\
        );

    \I__7968\ : InMux
    port map (
            O => \N__39195\,
            I => \N__39192\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__39192\,
            I => \sDAC_data_RNO_4Z0Z_9\
        );

    \I__7966\ : InMux
    port map (
            O => \N__39189\,
            I => \N__39186\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__39186\,
            I => \N__39183\
        );

    \I__7964\ : Span4Mux_v
    port map (
            O => \N__39183\,
            I => \N__39180\
        );

    \I__7963\ : Odrv4
    port map (
            O => \N__39180\,
            I => \sDAC_data_RNO_2Z0Z_9\
        );

    \I__7962\ : CascadeMux
    port map (
            O => \N__39177\,
            I => \sDAC_data_RNO_1Z0Z_9_cascade_\
        );

    \I__7961\ : CascadeMux
    port map (
            O => \N__39174\,
            I => \sDAC_data_2_9_cascade_\
        );

    \I__7960\ : InMux
    port map (
            O => \N__39171\,
            I => \N__39168\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__39168\,
            I => \N__39165\
        );

    \I__7958\ : Span4Mux_v
    port map (
            O => \N__39165\,
            I => \N__39162\
        );

    \I__7957\ : Span4Mux_h
    port map (
            O => \N__39162\,
            I => \N__39159\
        );

    \I__7956\ : Odrv4
    port map (
            O => \N__39159\,
            I => \sDAC_dataZ0Z_9\
        );

    \I__7955\ : CascadeMux
    port map (
            O => \N__39156\,
            I => \N__39153\
        );

    \I__7954\ : InMux
    port map (
            O => \N__39153\,
            I => \N__39150\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__39150\,
            I => \N__39147\
        );

    \I__7952\ : Odrv4
    port map (
            O => \N__39147\,
            I => \sDAC_data_RNO_15Z0Z_9\
        );

    \I__7951\ : InMux
    port map (
            O => \N__39144\,
            I => \N__39141\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__39141\,
            I => \N__39138\
        );

    \I__7949\ : Span4Mux_v
    port map (
            O => \N__39138\,
            I => \N__39135\
        );

    \I__7948\ : Odrv4
    port map (
            O => \N__39135\,
            I => \sDAC_data_RNO_14Z0Z_9\
        );

    \I__7947\ : InMux
    port map (
            O => \N__39132\,
            I => \N__39129\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__39129\,
            I => \sDAC_data_2_14_ns_1_9\
        );

    \I__7945\ : InMux
    port map (
            O => \N__39126\,
            I => \N__39123\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__39123\,
            I => \sDAC_data_RNO_29Z0Z_9\
        );

    \I__7943\ : InMux
    port map (
            O => \N__39120\,
            I => \N__39117\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__39117\,
            I => \N__39114\
        );

    \I__7941\ : Span4Mux_h
    port map (
            O => \N__39114\,
            I => \N__39111\
        );

    \I__7940\ : Odrv4
    port map (
            O => \N__39111\,
            I => \sDAC_data_RNO_30Z0Z_9\
        );

    \I__7939\ : CascadeMux
    port map (
            O => \N__39108\,
            I => \sDAC_data_2_32_ns_1_9_cascade_\
        );

    \I__7938\ : InMux
    port map (
            O => \N__39105\,
            I => \N__39102\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__39102\,
            I => \N__39099\
        );

    \I__7936\ : Odrv4
    port map (
            O => \N__39099\,
            I => \sDAC_data_RNO_20Z0Z_9\
        );

    \I__7935\ : CascadeMux
    port map (
            O => \N__39096\,
            I => \sDAC_data_RNO_10Z0Z_9_cascade_\
        );

    \I__7934\ : InMux
    port map (
            O => \N__39093\,
            I => \N__39090\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__39090\,
            I => \sDAC_data_RNO_11Z0Z_9\
        );

    \I__7932\ : InMux
    port map (
            O => \N__39087\,
            I => \N__39084\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__39084\,
            I => \sDAC_data_2_41_ns_1_9\
        );

    \I__7930\ : InMux
    port map (
            O => \N__39081\,
            I => \N__39078\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__39078\,
            I => \sDAC_mem_3Z0Z_4\
        );

    \I__7928\ : CascadeMux
    port map (
            O => \N__39075\,
            I => \sDAC_data_2_6_bm_1_7_cascade_\
        );

    \I__7927\ : InMux
    port map (
            O => \N__39072\,
            I => \N__39069\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__39069\,
            I => \sDAC_data_RNO_15Z0Z_7\
        );

    \I__7925\ : InMux
    port map (
            O => \N__39066\,
            I => \N__39063\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__39063\,
            I => \N__39060\
        );

    \I__7923\ : Odrv12
    port map (
            O => \N__39060\,
            I => \sDAC_mem_36Z0Z_5\
        );

    \I__7922\ : InMux
    port map (
            O => \N__39057\,
            I => \N__39054\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__39054\,
            I => \N__39051\
        );

    \I__7920\ : Odrv12
    port map (
            O => \N__39051\,
            I => \sDAC_mem_37Z0Z_5\
        );

    \I__7919\ : CascadeMux
    port map (
            O => \N__39048\,
            I => \sDAC_data_2_13_am_1_8_cascade_\
        );

    \I__7918\ : InMux
    port map (
            O => \N__39045\,
            I => \N__39042\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__39042\,
            I => \N__39039\
        );

    \I__7916\ : Span4Mux_v
    port map (
            O => \N__39039\,
            I => \N__39036\
        );

    \I__7915\ : Odrv4
    port map (
            O => \N__39036\,
            I => \sDAC_mem_5Z0Z_5\
        );

    \I__7914\ : InMux
    port map (
            O => \N__39033\,
            I => \N__39030\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__39030\,
            I => \sDAC_mem_4Z0Z_5\
        );

    \I__7912\ : InMux
    port map (
            O => \N__39027\,
            I => \N__39024\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__39024\,
            I => \N__39021\
        );

    \I__7910\ : Odrv12
    port map (
            O => \N__39021\,
            I => \sDAC_mem_36Z0Z_6\
        );

    \I__7909\ : InMux
    port map (
            O => \N__39018\,
            I => \N__39015\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__39015\,
            I => \N__39012\
        );

    \I__7907\ : Odrv12
    port map (
            O => \N__39012\,
            I => \sDAC_mem_37Z0Z_6\
        );

    \I__7906\ : CascadeMux
    port map (
            O => \N__39009\,
            I => \sDAC_data_2_13_am_1_9_cascade_\
        );

    \I__7905\ : InMux
    port map (
            O => \N__39006\,
            I => \N__39003\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__39003\,
            I => \N__39000\
        );

    \I__7903\ : Span4Mux_v
    port map (
            O => \N__39000\,
            I => \N__38997\
        );

    \I__7902\ : Odrv4
    port map (
            O => \N__38997\,
            I => \sDAC_mem_5Z0Z_6\
        );

    \I__7901\ : InMux
    port map (
            O => \N__38994\,
            I => \N__38991\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__38991\,
            I => \sDAC_mem_4Z0Z_6\
        );

    \I__7899\ : InMux
    port map (
            O => \N__38988\,
            I => \N__38985\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__38985\,
            I => \N__38982\
        );

    \I__7897\ : Span4Mux_v
    port map (
            O => \N__38982\,
            I => \N__38979\
        );

    \I__7896\ : Odrv4
    port map (
            O => \N__38979\,
            I => \sDAC_mem_6Z0Z_7\
        );

    \I__7895\ : CascadeMux
    port map (
            O => \N__38976\,
            I => \sDAC_data_2_13_bm_1_10_cascade_\
        );

    \I__7894\ : InMux
    port map (
            O => \N__38973\,
            I => \N__38970\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__38970\,
            I => \N__38967\
        );

    \I__7892\ : Span4Mux_v
    port map (
            O => \N__38967\,
            I => \N__38964\
        );

    \I__7891\ : Odrv4
    port map (
            O => \N__38964\,
            I => \sDAC_mem_7Z0Z_7\
        );

    \I__7890\ : InMux
    port map (
            O => \N__38961\,
            I => \N__38958\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__38958\,
            I => \sDAC_mem_20Z0Z_6\
        );

    \I__7888\ : InMux
    port map (
            O => \N__38955\,
            I => \N__38952\
        );

    \I__7887\ : LocalMux
    port map (
            O => \N__38952\,
            I => \N__38949\
        );

    \I__7886\ : Odrv12
    port map (
            O => \N__38949\,
            I => \sDAC_mem_23Z0Z_7\
        );

    \I__7885\ : InMux
    port map (
            O => \N__38946\,
            I => \N__38943\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__38943\,
            I => \N__38940\
        );

    \I__7883\ : Span4Mux_h
    port map (
            O => \N__38940\,
            I => \N__38937\
        );

    \I__7882\ : Span4Mux_h
    port map (
            O => \N__38937\,
            I => \N__38934\
        );

    \I__7881\ : Odrv4
    port map (
            O => \N__38934\,
            I => \sDAC_mem_22Z0Z_7\
        );

    \I__7880\ : InMux
    port map (
            O => \N__38931\,
            I => \N__38928\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__38928\,
            I => \N__38925\
        );

    \I__7878\ : Odrv12
    port map (
            O => \N__38925\,
            I => \sDAC_mem_23Z0Z_0\
        );

    \I__7877\ : InMux
    port map (
            O => \N__38922\,
            I => \N__38919\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__38919\,
            I => \N__38916\
        );

    \I__7875\ : Span4Mux_h
    port map (
            O => \N__38916\,
            I => \N__38913\
        );

    \I__7874\ : Span4Mux_h
    port map (
            O => \N__38913\,
            I => \N__38910\
        );

    \I__7873\ : Odrv4
    port map (
            O => \N__38910\,
            I => \sDAC_mem_22Z0Z_0\
        );

    \I__7872\ : CascadeMux
    port map (
            O => \N__38907\,
            I => \sDAC_data_2_13_bm_1_7_cascade_\
        );

    \I__7871\ : InMux
    port map (
            O => \N__38904\,
            I => \N__38901\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__38901\,
            I => \N__38898\
        );

    \I__7869\ : Span4Mux_v
    port map (
            O => \N__38898\,
            I => \N__38895\
        );

    \I__7868\ : Odrv4
    port map (
            O => \N__38895\,
            I => \sDAC_mem_7Z0Z_4\
        );

    \I__7867\ : InMux
    port map (
            O => \N__38892\,
            I => \N__38889\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__38889\,
            I => \sDAC_data_RNO_5Z0Z_7\
        );

    \I__7865\ : CascadeMux
    port map (
            O => \N__38886\,
            I => \N__38883\
        );

    \I__7864\ : InMux
    port map (
            O => \N__38883\,
            I => \N__38880\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__38880\,
            I => \N__38877\
        );

    \I__7862\ : Span4Mux_h
    port map (
            O => \N__38877\,
            I => \N__38874\
        );

    \I__7861\ : Span4Mux_v
    port map (
            O => \N__38874\,
            I => \N__38871\
        );

    \I__7860\ : Odrv4
    port map (
            O => \N__38871\,
            I => \sDAC_data_RNO_30Z0Z_7\
        );

    \I__7859\ : InMux
    port map (
            O => \N__38868\,
            I => \N__38865\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__38865\,
            I => \sDAC_data_RNO_29Z0Z_7\
        );

    \I__7857\ : InMux
    port map (
            O => \N__38862\,
            I => \N__38859\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__38859\,
            I => \sDAC_data_2_32_ns_1_7\
        );

    \I__7855\ : CascadeMux
    port map (
            O => \N__38856\,
            I => \N__38853\
        );

    \I__7854\ : InMux
    port map (
            O => \N__38853\,
            I => \N__38850\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__38850\,
            I => \N__38847\
        );

    \I__7852\ : Span4Mux_v
    port map (
            O => \N__38847\,
            I => \N__38844\
        );

    \I__7851\ : Odrv4
    port map (
            O => \N__38844\,
            I => \sDAC_mem_34Z0Z_4\
        );

    \I__7850\ : InMux
    port map (
            O => \N__38841\,
            I => \N__38838\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__38838\,
            I => \N__38835\
        );

    \I__7848\ : Span4Mux_h
    port map (
            O => \N__38835\,
            I => \N__38832\
        );

    \I__7847\ : Odrv4
    port map (
            O => \N__38832\,
            I => \sDAC_mem_2Z0Z_4\
        );

    \I__7846\ : InMux
    port map (
            O => \N__38829\,
            I => \N__38826\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__38826\,
            I => \N__38823\
        );

    \I__7844\ : Span4Mux_h
    port map (
            O => \N__38823\,
            I => \N__38820\
        );

    \I__7843\ : Odrv4
    port map (
            O => \N__38820\,
            I => \sDAC_mem_8Z0Z_4\
        );

    \I__7842\ : InMux
    port map (
            O => \N__38817\,
            I => \N__38814\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__38814\,
            I => \N__38811\
        );

    \I__7840\ : Odrv4
    port map (
            O => \N__38811\,
            I => \sDAC_mem_8Z0Z_6\
        );

    \I__7839\ : InMux
    port map (
            O => \N__38808\,
            I => \N__38805\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__38805\,
            I => \N__38802\
        );

    \I__7837\ : Span4Mux_v
    port map (
            O => \N__38802\,
            I => \N__38799\
        );

    \I__7836\ : Odrv4
    port map (
            O => \N__38799\,
            I => \sDAC_mem_8Z0Z_7\
        );

    \I__7835\ : CEMux
    port map (
            O => \N__38796\,
            I => \N__38793\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__38793\,
            I => \sDAC_mem_8_1_sqmuxa\
        );

    \I__7833\ : InMux
    port map (
            O => \N__38790\,
            I => \N__38787\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__38787\,
            I => \N__38784\
        );

    \I__7831\ : Odrv4
    port map (
            O => \N__38784\,
            I => \sDAC_data_RNO_20Z0Z_7\
        );

    \I__7830\ : InMux
    port map (
            O => \N__38781\,
            I => \N__38778\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__38778\,
            I => \sDAC_mem_20Z0Z_4\
        );

    \I__7828\ : InMux
    port map (
            O => \N__38775\,
            I => \N__38772\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__38772\,
            I => \sDAC_mem_20Z0Z_5\
        );

    \I__7826\ : InMux
    port map (
            O => \N__38769\,
            I => \N__38766\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__38766\,
            I => \N__38763\
        );

    \I__7824\ : Odrv4
    port map (
            O => \N__38763\,
            I => \sDAC_mem_37Z0Z_2\
        );

    \I__7823\ : InMux
    port map (
            O => \N__38760\,
            I => \N__38757\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__38757\,
            I => \N__38754\
        );

    \I__7821\ : Odrv4
    port map (
            O => \N__38754\,
            I => \sDAC_mem_37Z0Z_3\
        );

    \I__7820\ : InMux
    port map (
            O => \N__38751\,
            I => \N__38748\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__38748\,
            I => \N__38745\
        );

    \I__7818\ : Odrv4
    port map (
            O => \N__38745\,
            I => \sDAC_mem_37Z0Z_4\
        );

    \I__7817\ : InMux
    port map (
            O => \N__38742\,
            I => \N__38739\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__38739\,
            I => \N__38736\
        );

    \I__7815\ : Odrv4
    port map (
            O => \N__38736\,
            I => \sDAC_mem_8Z0Z_2\
        );

    \I__7814\ : InMux
    port map (
            O => \N__38733\,
            I => \N__38730\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__38730\,
            I => \N__38727\
        );

    \I__7812\ : Span4Mux_h
    port map (
            O => \N__38727\,
            I => \N__38724\
        );

    \I__7811\ : Odrv4
    port map (
            O => \N__38724\,
            I => \sDAC_mem_36Z0Z_2\
        );

    \I__7810\ : InMux
    port map (
            O => \N__38721\,
            I => \N__38718\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__38718\,
            I => \N__38715\
        );

    \I__7808\ : Span4Mux_h
    port map (
            O => \N__38715\,
            I => \N__38712\
        );

    \I__7807\ : Odrv4
    port map (
            O => \N__38712\,
            I => \sDAC_mem_36Z0Z_3\
        );

    \I__7806\ : InMux
    port map (
            O => \N__38709\,
            I => \N__38706\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__38706\,
            I => \N__38703\
        );

    \I__7804\ : Span4Mux_v
    port map (
            O => \N__38703\,
            I => \N__38700\
        );

    \I__7803\ : Odrv4
    port map (
            O => \N__38700\,
            I => \sDAC_mem_36Z0Z_4\
        );

    \I__7802\ : InMux
    port map (
            O => \N__38697\,
            I => \N__38694\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__38694\,
            I => \N__38691\
        );

    \I__7800\ : Span4Mux_v
    port map (
            O => \N__38691\,
            I => \N__38688\
        );

    \I__7799\ : Odrv4
    port map (
            O => \N__38688\,
            I => \sDAC_mem_31Z0Z_2\
        );

    \I__7798\ : InMux
    port map (
            O => \N__38685\,
            I => \N__38682\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__38682\,
            I => \sDAC_data_RNO_24Z0Z_5\
        );

    \I__7796\ : InMux
    port map (
            O => \N__38679\,
            I => \N__38676\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__38676\,
            I => \sDAC_mem_24Z0Z_2\
        );

    \I__7794\ : CascadeMux
    port map (
            O => \N__38673\,
            I => \N__38670\
        );

    \I__7793\ : InMux
    port map (
            O => \N__38670\,
            I => \N__38667\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__38667\,
            I => \sDAC_data_RNO_31Z0Z_6\
        );

    \I__7791\ : InMux
    port map (
            O => \N__38664\,
            I => \N__38661\
        );

    \I__7790\ : LocalMux
    port map (
            O => \N__38661\,
            I => \sDAC_data_2_39_ns_1_6\
        );

    \I__7789\ : InMux
    port map (
            O => \N__38658\,
            I => \N__38655\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__38655\,
            I => \N__38652\
        );

    \I__7787\ : Odrv4
    port map (
            O => \N__38652\,
            I => \sDAC_mem_29Z0Z_4\
        );

    \I__7786\ : InMux
    port map (
            O => \N__38649\,
            I => \N__38646\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__38646\,
            I => \N__38643\
        );

    \I__7784\ : Odrv4
    port map (
            O => \N__38643\,
            I => \sDAC_data_RNO_23Z0Z_7\
        );

    \I__7783\ : InMux
    port map (
            O => \N__38640\,
            I => \N__38637\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__38637\,
            I => \N__38634\
        );

    \I__7781\ : Odrv12
    port map (
            O => \N__38634\,
            I => \sDAC_mem_26Z0Z_3\
        );

    \I__7780\ : InMux
    port map (
            O => \N__38631\,
            I => \N__38628\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__38628\,
            I => \sDAC_data_RNO_32Z0Z_6\
        );

    \I__7778\ : InMux
    port map (
            O => \N__38625\,
            I => \N__38622\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__38622\,
            I => \N__38619\
        );

    \I__7776\ : Span4Mux_h
    port map (
            O => \N__38619\,
            I => \N__38616\
        );

    \I__7775\ : Span4Mux_v
    port map (
            O => \N__38616\,
            I => \N__38613\
        );

    \I__7774\ : Odrv4
    port map (
            O => \N__38613\,
            I => \sDAC_mem_24Z0Z_0\
        );

    \I__7773\ : InMux
    port map (
            O => \N__38610\,
            I => \N__38607\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__38607\,
            I => \N__38604\
        );

    \I__7771\ : Span4Mux_h
    port map (
            O => \N__38604\,
            I => \N__38601\
        );

    \I__7770\ : Sp12to4
    port map (
            O => \N__38601\,
            I => \N__38598\
        );

    \I__7769\ : Odrv12
    port map (
            O => \N__38598\,
            I => \sDAC_mem_17Z0Z_3\
        );

    \I__7768\ : InMux
    port map (
            O => \N__38595\,
            I => \N__38591\
        );

    \I__7767\ : InMux
    port map (
            O => \N__38594\,
            I => \N__38588\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__38591\,
            I => \N__38585\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__38588\,
            I => \N__38582\
        );

    \I__7764\ : Span4Mux_v
    port map (
            O => \N__38585\,
            I => \N__38579\
        );

    \I__7763\ : Span4Mux_v
    port map (
            O => \N__38582\,
            I => \N__38576\
        );

    \I__7762\ : Span4Mux_h
    port map (
            O => \N__38579\,
            I => \N__38573\
        );

    \I__7761\ : Span4Mux_h
    port map (
            O => \N__38576\,
            I => \N__38570\
        );

    \I__7760\ : Odrv4
    port map (
            O => \N__38573\,
            I => \spi_slave_inst.spi_miso\
        );

    \I__7759\ : Odrv4
    port map (
            O => \N__38570\,
            I => \spi_slave_inst.spi_miso\
        );

    \I__7758\ : InMux
    port map (
            O => \N__38565\,
            I => \N__38558\
        );

    \I__7757\ : InMux
    port map (
            O => \N__38564\,
            I => \N__38558\
        );

    \I__7756\ : InMux
    port map (
            O => \N__38563\,
            I => \N__38555\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__38558\,
            I => \N__38549\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__38555\,
            I => \N__38546\
        );

    \I__7753\ : InMux
    port map (
            O => \N__38554\,
            I => \N__38541\
        );

    \I__7752\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38541\
        );

    \I__7751\ : InMux
    port map (
            O => \N__38552\,
            I => \N__38538\
        );

    \I__7750\ : Span4Mux_v
    port map (
            O => \N__38549\,
            I => \N__38535\
        );

    \I__7749\ : Span4Mux_h
    port map (
            O => \N__38546\,
            I => \N__38528\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__38541\,
            I => \N__38528\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__38538\,
            I => \N__38528\
        );

    \I__7746\ : Span4Mux_v
    port map (
            O => \N__38535\,
            I => \N__38522\
        );

    \I__7745\ : Span4Mux_h
    port map (
            O => \N__38528\,
            I => \N__38519\
        );

    \I__7744\ : InMux
    port map (
            O => \N__38527\,
            I => \N__38512\
        );

    \I__7743\ : InMux
    port map (
            O => \N__38526\,
            I => \N__38512\
        );

    \I__7742\ : InMux
    port map (
            O => \N__38525\,
            I => \N__38512\
        );

    \I__7741\ : Sp12to4
    port map (
            O => \N__38522\,
            I => \N__38509\
        );

    \I__7740\ : Span4Mux_v
    port map (
            O => \N__38519\,
            I => \N__38506\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__38512\,
            I => \N__38503\
        );

    \I__7738\ : Span12Mux_h
    port map (
            O => \N__38509\,
            I => \N__38496\
        );

    \I__7737\ : Sp12to4
    port map (
            O => \N__38506\,
            I => \N__38496\
        );

    \I__7736\ : Span12Mux_s11_v
    port map (
            O => \N__38503\,
            I => \N__38496\
        );

    \I__7735\ : Span12Mux_h
    port map (
            O => \N__38496\,
            I => \N__38493\
        );

    \I__7734\ : Odrv12
    port map (
            O => \N__38493\,
            I => spi_select_c
        );

    \I__7733\ : IoInMux
    port map (
            O => \N__38490\,
            I => \N__38487\
        );

    \I__7732\ : LocalMux
    port map (
            O => \N__38487\,
            I => \N__38484\
        );

    \I__7731\ : Span4Mux_s3_v
    port map (
            O => \N__38484\,
            I => \N__38481\
        );

    \I__7730\ : Span4Mux_h
    port map (
            O => \N__38481\,
            I => \N__38478\
        );

    \I__7729\ : Span4Mux_h
    port map (
            O => \N__38478\,
            I => \N__38475\
        );

    \I__7728\ : Odrv4
    port map (
            O => \N__38475\,
            I => spi_miso_ft_c
        );

    \I__7727\ : CascadeMux
    port map (
            O => \N__38472\,
            I => \sDAC_data_2_39_ns_1_7_cascade_\
        );

    \I__7726\ : InMux
    port map (
            O => \N__38469\,
            I => \N__38466\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__38466\,
            I => \N__38463\
        );

    \I__7724\ : Span12Mux_v
    port map (
            O => \N__38463\,
            I => \N__38460\
        );

    \I__7723\ : Odrv12
    port map (
            O => \N__38460\,
            I => \sDAC_data_RNO_11Z0Z_7\
        );

    \I__7722\ : InMux
    port map (
            O => \N__38457\,
            I => \N__38454\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__38454\,
            I => \sDAC_mem_28Z0Z_3\
        );

    \I__7720\ : InMux
    port map (
            O => \N__38451\,
            I => \N__38448\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__38448\,
            I => \N__38445\
        );

    \I__7718\ : Odrv4
    port map (
            O => \N__38445\,
            I => \sDAC_mem_26Z0Z_4\
        );

    \I__7717\ : InMux
    port map (
            O => \N__38442\,
            I => \N__38439\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__38439\,
            I => \sDAC_data_RNO_32Z0Z_7\
        );

    \I__7715\ : InMux
    port map (
            O => \N__38436\,
            I => \N__38433\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__38433\,
            I => \N__38430\
        );

    \I__7713\ : Span4Mux_v
    port map (
            O => \N__38430\,
            I => \N__38427\
        );

    \I__7712\ : Odrv4
    port map (
            O => \N__38427\,
            I => \sDAC_mem_31Z0Z_3\
        );

    \I__7711\ : InMux
    port map (
            O => \N__38424\,
            I => \N__38421\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__38421\,
            I => \sDAC_data_RNO_24Z0Z_6\
        );

    \I__7709\ : CascadeMux
    port map (
            O => \N__38418\,
            I => \sDAC_data_RNO_31Z0Z_5_cascade_\
        );

    \I__7708\ : CascadeMux
    port map (
            O => \N__38415\,
            I => \sDAC_data_2_39_ns_1_5_cascade_\
        );

    \I__7707\ : InMux
    port map (
            O => \N__38412\,
            I => \N__38409\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__38409\,
            I => \N__38406\
        );

    \I__7705\ : Span4Mux_v
    port map (
            O => \N__38406\,
            I => \N__38403\
        );

    \I__7704\ : Span4Mux_v
    port map (
            O => \N__38403\,
            I => \N__38400\
        );

    \I__7703\ : Odrv4
    port map (
            O => \N__38400\,
            I => \sDAC_data_RNO_11Z0Z_5\
        );

    \I__7702\ : InMux
    port map (
            O => \N__38397\,
            I => \N__38394\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__38394\,
            I => \N__38391\
        );

    \I__7700\ : Odrv12
    port map (
            O => \N__38391\,
            I => \sDAC_mem_26Z0Z_2\
        );

    \I__7699\ : InMux
    port map (
            O => \N__38388\,
            I => \N__38385\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__38385\,
            I => \N__38382\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__38382\,
            I => \sDAC_data_RNO_32Z0Z_5\
        );

    \I__7696\ : InMux
    port map (
            O => \N__38379\,
            I => \N__38376\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__38376\,
            I => \N__38373\
        );

    \I__7694\ : Odrv4
    port map (
            O => \N__38373\,
            I => \sDAC_mem_29Z0Z_2\
        );

    \I__7693\ : InMux
    port map (
            O => \N__38370\,
            I => \N__38367\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__38367\,
            I => \sDAC_data_RNO_23Z0Z_5\
        );

    \I__7691\ : InMux
    port map (
            O => \N__38364\,
            I => \N__38361\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__38361\,
            I => \N__38358\
        );

    \I__7689\ : Odrv12
    port map (
            O => \N__38358\,
            I => \sDAC_mem_29Z0Z_5\
        );

    \I__7688\ : InMux
    port map (
            O => \N__38355\,
            I => \N__38352\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__38352\,
            I => \N__38349\
        );

    \I__7686\ : Odrv12
    port map (
            O => \N__38349\,
            I => \sDAC_mem_29Z0Z_6\
        );

    \I__7685\ : CEMux
    port map (
            O => \N__38346\,
            I => \N__38343\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__38343\,
            I => \N__38340\
        );

    \I__7683\ : Span4Mux_h
    port map (
            O => \N__38340\,
            I => \N__38337\
        );

    \I__7682\ : Span4Mux_v
    port map (
            O => \N__38337\,
            I => \N__38334\
        );

    \I__7681\ : Odrv4
    port map (
            O => \N__38334\,
            I => \sDAC_mem_29_1_sqmuxa\
        );

    \I__7680\ : InMux
    port map (
            O => \N__38331\,
            I => \N__38328\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__38328\,
            I => \sDAC_mem_29Z0Z_3\
        );

    \I__7678\ : InMux
    port map (
            O => \N__38325\,
            I => \N__38322\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__38322\,
            I => \sDAC_data_RNO_23Z0Z_6\
        );

    \I__7676\ : InMux
    port map (
            O => \N__38319\,
            I => \N__38316\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__38316\,
            I => \N__38313\
        );

    \I__7674\ : Span4Mux_h
    port map (
            O => \N__38313\,
            I => \N__38310\
        );

    \I__7673\ : Odrv4
    port map (
            O => \N__38310\,
            I => \sDAC_mem_24Z0Z_4\
        );

    \I__7672\ : CascadeMux
    port map (
            O => \N__38307\,
            I => \sDAC_data_RNO_31Z0Z_7_cascade_\
        );

    \I__7671\ : CascadeMux
    port map (
            O => \N__38304\,
            I => \sDAC_data_RNO_18Z0Z_9_cascade_\
        );

    \I__7670\ : InMux
    port map (
            O => \N__38301\,
            I => \N__38298\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__38298\,
            I => \sDAC_data_RNO_19Z0Z_9\
        );

    \I__7668\ : InMux
    port map (
            O => \N__38295\,
            I => \N__38292\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__38292\,
            I => \N__38289\
        );

    \I__7666\ : Span4Mux_v
    port map (
            O => \N__38289\,
            I => \N__38286\
        );

    \I__7665\ : Odrv4
    port map (
            O => \N__38286\,
            I => \sDAC_data_2_24_ns_1_9\
        );

    \I__7664\ : InMux
    port map (
            O => \N__38283\,
            I => \N__38279\
        );

    \I__7663\ : InMux
    port map (
            O => \N__38282\,
            I => \N__38276\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__38279\,
            I => \N__38273\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__38276\,
            I => \sCounterADCZ0Z_1\
        );

    \I__7660\ : Odrv12
    port map (
            O => \N__38273\,
            I => \sCounterADCZ0Z_1\
        );

    \I__7659\ : InMux
    port map (
            O => \N__38268\,
            I => \N__38264\
        );

    \I__7658\ : InMux
    port map (
            O => \N__38267\,
            I => \N__38261\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__38264\,
            I => \N__38258\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__38261\,
            I => \sCounterADCZ0Z_0\
        );

    \I__7655\ : Odrv4
    port map (
            O => \N__38258\,
            I => \sCounterADCZ0Z_0\
        );

    \I__7654\ : InMux
    port map (
            O => \N__38253\,
            I => \N__38250\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__38250\,
            I => \un11_sacqtime_NE_3\
        );

    \I__7652\ : InMux
    port map (
            O => \N__38247\,
            I => \N__38244\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__38244\,
            I => \un11_sacqtime_NE_2\
        );

    \I__7650\ : CascadeMux
    port map (
            O => \N__38241\,
            I => \un11_sacqtime_NE_0_0_cascade_\
        );

    \I__7649\ : InMux
    port map (
            O => \N__38238\,
            I => \N__38235\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__38235\,
            I => \N__38232\
        );

    \I__7647\ : Odrv4
    port map (
            O => \N__38232\,
            I => \un11_sacqtime_NE_1\
        );

    \I__7646\ : CascadeMux
    port map (
            O => \N__38229\,
            I => \N__38222\
        );

    \I__7645\ : InMux
    port map (
            O => \N__38228\,
            I => \N__38213\
        );

    \I__7644\ : InMux
    port map (
            O => \N__38227\,
            I => \N__38213\
        );

    \I__7643\ : InMux
    port map (
            O => \N__38226\,
            I => \N__38213\
        );

    \I__7642\ : InMux
    port map (
            O => \N__38225\,
            I => \N__38213\
        );

    \I__7641\ : InMux
    port map (
            O => \N__38222\,
            I => \N__38210\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__38213\,
            I => \N__38207\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__38210\,
            I => \N__38200\
        );

    \I__7638\ : Span4Mux_h
    port map (
            O => \N__38207\,
            I => \N__38197\
        );

    \I__7637\ : InMux
    port map (
            O => \N__38206\,
            I => \N__38188\
        );

    \I__7636\ : InMux
    port map (
            O => \N__38205\,
            I => \N__38188\
        );

    \I__7635\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38188\
        );

    \I__7634\ : InMux
    port map (
            O => \N__38203\,
            I => \N__38188\
        );

    \I__7633\ : Span4Mux_v
    port map (
            O => \N__38200\,
            I => \N__38185\
        );

    \I__7632\ : Span4Mux_h
    port map (
            O => \N__38197\,
            I => \N__38178\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__38188\,
            I => \N__38178\
        );

    \I__7630\ : Span4Mux_h
    port map (
            O => \N__38185\,
            I => \N__38178\
        );

    \I__7629\ : Odrv4
    port map (
            O => \N__38178\,
            I => \un11_sacqtime_NE_0\
        );

    \I__7628\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38172\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__38172\,
            I => \sDAC_mem_31Z0Z_6\
        );

    \I__7626\ : InMux
    port map (
            O => \N__38169\,
            I => \N__38166\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__38166\,
            I => \N__38163\
        );

    \I__7624\ : Span4Mux_v
    port map (
            O => \N__38163\,
            I => \N__38160\
        );

    \I__7623\ : Odrv4
    port map (
            O => \N__38160\,
            I => \sDAC_data_RNO_24Z0Z_9\
        );

    \I__7622\ : InMux
    port map (
            O => \N__38157\,
            I => \N__38154\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__38154\,
            I => \sDAC_mem_24Z0Z_5\
        );

    \I__7620\ : CascadeMux
    port map (
            O => \N__38151\,
            I => \N__38148\
        );

    \I__7619\ : InMux
    port map (
            O => \N__38148\,
            I => \N__38145\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__38145\,
            I => \N__38142\
        );

    \I__7617\ : Span4Mux_h
    port map (
            O => \N__38142\,
            I => \N__38139\
        );

    \I__7616\ : Span4Mux_v
    port map (
            O => \N__38139\,
            I => \N__38136\
        );

    \I__7615\ : Odrv4
    port map (
            O => \N__38136\,
            I => \sDAC_data_RNO_31Z0Z_9\
        );

    \I__7614\ : InMux
    port map (
            O => \N__38133\,
            I => \N__38130\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__38130\,
            I => \N__38127\
        );

    \I__7612\ : Span4Mux_v
    port map (
            O => \N__38127\,
            I => \N__38124\
        );

    \I__7611\ : Odrv4
    port map (
            O => \N__38124\,
            I => \sDAC_data_RNO_32Z0Z_9\
        );

    \I__7610\ : InMux
    port map (
            O => \N__38121\,
            I => \N__38118\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__38118\,
            I => \N__38115\
        );

    \I__7608\ : Odrv4
    port map (
            O => \N__38115\,
            I => \sDAC_data_2_39_ns_1_9\
        );

    \I__7607\ : InMux
    port map (
            O => \N__38112\,
            I => \N__38109\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__38109\,
            I => \N__38106\
        );

    \I__7605\ : Span4Mux_v
    port map (
            O => \N__38106\,
            I => \N__38103\
        );

    \I__7604\ : Odrv4
    port map (
            O => \N__38103\,
            I => \sDAC_mem_26Z0Z_0\
        );

    \I__7603\ : InMux
    port map (
            O => \N__38100\,
            I => \N__38097\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__38097\,
            I => \sDAC_mem_26Z0Z_5\
        );

    \I__7601\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38091\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__38091\,
            I => \N__38088\
        );

    \I__7599\ : Span4Mux_v
    port map (
            O => \N__38088\,
            I => \N__38085\
        );

    \I__7598\ : Odrv4
    port map (
            O => \N__38085\,
            I => \sDAC_mem_26Z0Z_6\
        );

    \I__7597\ : CascadeMux
    port map (
            O => \N__38082\,
            I => \N__38065\
        );

    \I__7596\ : CascadeMux
    port map (
            O => \N__38081\,
            I => \N__38062\
        );

    \I__7595\ : CascadeMux
    port map (
            O => \N__38080\,
            I => \N__38059\
        );

    \I__7594\ : CascadeMux
    port map (
            O => \N__38079\,
            I => \N__38056\
        );

    \I__7593\ : CascadeMux
    port map (
            O => \N__38078\,
            I => \N__38053\
        );

    \I__7592\ : CascadeMux
    port map (
            O => \N__38077\,
            I => \N__38050\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__38076\,
            I => \N__38047\
        );

    \I__7590\ : CascadeMux
    port map (
            O => \N__38075\,
            I => \N__38044\
        );

    \I__7589\ : CascadeMux
    port map (
            O => \N__38074\,
            I => \N__38040\
        );

    \I__7588\ : CascadeMux
    port map (
            O => \N__38073\,
            I => \N__38037\
        );

    \I__7587\ : CascadeMux
    port map (
            O => \N__38072\,
            I => \N__38034\
        );

    \I__7586\ : CascadeMux
    port map (
            O => \N__38071\,
            I => \N__38030\
        );

    \I__7585\ : CascadeMux
    port map (
            O => \N__38070\,
            I => \N__38027\
        );

    \I__7584\ : CascadeMux
    port map (
            O => \N__38069\,
            I => \N__38024\
        );

    \I__7583\ : CascadeMux
    port map (
            O => \N__38068\,
            I => \N__38021\
        );

    \I__7582\ : InMux
    port map (
            O => \N__38065\,
            I => \N__38009\
        );

    \I__7581\ : InMux
    port map (
            O => \N__38062\,
            I => \N__38009\
        );

    \I__7580\ : InMux
    port map (
            O => \N__38059\,
            I => \N__38009\
        );

    \I__7579\ : InMux
    port map (
            O => \N__38056\,
            I => \N__38009\
        );

    \I__7578\ : InMux
    port map (
            O => \N__38053\,
            I => \N__38000\
        );

    \I__7577\ : InMux
    port map (
            O => \N__38050\,
            I => \N__38000\
        );

    \I__7576\ : InMux
    port map (
            O => \N__38047\,
            I => \N__38000\
        );

    \I__7575\ : InMux
    port map (
            O => \N__38044\,
            I => \N__38000\
        );

    \I__7574\ : InMux
    port map (
            O => \N__38043\,
            I => \N__37991\
        );

    \I__7573\ : InMux
    port map (
            O => \N__38040\,
            I => \N__37991\
        );

    \I__7572\ : InMux
    port map (
            O => \N__38037\,
            I => \N__37991\
        );

    \I__7571\ : InMux
    port map (
            O => \N__38034\,
            I => \N__37991\
        );

    \I__7570\ : InMux
    port map (
            O => \N__38033\,
            I => \N__37982\
        );

    \I__7569\ : InMux
    port map (
            O => \N__38030\,
            I => \N__37982\
        );

    \I__7568\ : InMux
    port map (
            O => \N__38027\,
            I => \N__37982\
        );

    \I__7567\ : InMux
    port map (
            O => \N__38024\,
            I => \N__37982\
        );

    \I__7566\ : InMux
    port map (
            O => \N__38021\,
            I => \N__37977\
        );

    \I__7565\ : InMux
    port map (
            O => \N__38020\,
            I => \N__37977\
        );

    \I__7564\ : InMux
    port map (
            O => \N__38019\,
            I => \N__37972\
        );

    \I__7563\ : InMux
    port map (
            O => \N__38018\,
            I => \N__37972\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__38009\,
            I => \N__37959\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__38000\,
            I => \N__37959\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__37991\,
            I => \N__37954\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__37982\,
            I => \N__37954\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__37977\,
            I => \N__37951\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__37972\,
            I => \N__37948\
        );

    \I__7556\ : CascadeMux
    port map (
            O => \N__37971\,
            I => \N__37945\
        );

    \I__7555\ : CascadeMux
    port map (
            O => \N__37970\,
            I => \N__37941\
        );

    \I__7554\ : CascadeMux
    port map (
            O => \N__37969\,
            I => \N__37937\
        );

    \I__7553\ : CascadeMux
    port map (
            O => \N__37968\,
            I => \N__37933\
        );

    \I__7552\ : CascadeMux
    port map (
            O => \N__37967\,
            I => \N__37925\
        );

    \I__7551\ : CascadeMux
    port map (
            O => \N__37966\,
            I => \N__37921\
        );

    \I__7550\ : CascadeMux
    port map (
            O => \N__37965\,
            I => \N__37917\
        );

    \I__7549\ : CascadeMux
    port map (
            O => \N__37964\,
            I => \N__37913\
        );

    \I__7548\ : Span4Mux_v
    port map (
            O => \N__37959\,
            I => \N__37904\
        );

    \I__7547\ : Span4Mux_v
    port map (
            O => \N__37954\,
            I => \N__37898\
        );

    \I__7546\ : Span4Mux_v
    port map (
            O => \N__37951\,
            I => \N__37898\
        );

    \I__7545\ : Span4Mux_h
    port map (
            O => \N__37948\,
            I => \N__37895\
        );

    \I__7544\ : InMux
    port map (
            O => \N__37945\,
            I => \N__37878\
        );

    \I__7543\ : InMux
    port map (
            O => \N__37944\,
            I => \N__37878\
        );

    \I__7542\ : InMux
    port map (
            O => \N__37941\,
            I => \N__37878\
        );

    \I__7541\ : InMux
    port map (
            O => \N__37940\,
            I => \N__37878\
        );

    \I__7540\ : InMux
    port map (
            O => \N__37937\,
            I => \N__37878\
        );

    \I__7539\ : InMux
    port map (
            O => \N__37936\,
            I => \N__37878\
        );

    \I__7538\ : InMux
    port map (
            O => \N__37933\,
            I => \N__37878\
        );

    \I__7537\ : InMux
    port map (
            O => \N__37932\,
            I => \N__37878\
        );

    \I__7536\ : CascadeMux
    port map (
            O => \N__37931\,
            I => \N__37875\
        );

    \I__7535\ : CascadeMux
    port map (
            O => \N__37930\,
            I => \N__37870\
        );

    \I__7534\ : CascadeMux
    port map (
            O => \N__37929\,
            I => \N__37866\
        );

    \I__7533\ : CascadeMux
    port map (
            O => \N__37928\,
            I => \N__37862\
        );

    \I__7532\ : InMux
    port map (
            O => \N__37925\,
            I => \N__37845\
        );

    \I__7531\ : InMux
    port map (
            O => \N__37924\,
            I => \N__37845\
        );

    \I__7530\ : InMux
    port map (
            O => \N__37921\,
            I => \N__37845\
        );

    \I__7529\ : InMux
    port map (
            O => \N__37920\,
            I => \N__37845\
        );

    \I__7528\ : InMux
    port map (
            O => \N__37917\,
            I => \N__37845\
        );

    \I__7527\ : InMux
    port map (
            O => \N__37916\,
            I => \N__37845\
        );

    \I__7526\ : InMux
    port map (
            O => \N__37913\,
            I => \N__37845\
        );

    \I__7525\ : InMux
    port map (
            O => \N__37912\,
            I => \N__37845\
        );

    \I__7524\ : CascadeMux
    port map (
            O => \N__37911\,
            I => \N__37842\
        );

    \I__7523\ : CascadeMux
    port map (
            O => \N__37910\,
            I => \N__37838\
        );

    \I__7522\ : CascadeMux
    port map (
            O => \N__37909\,
            I => \N__37834\
        );

    \I__7521\ : CascadeMux
    port map (
            O => \N__37908\,
            I => \N__37830\
        );

    \I__7520\ : CascadeMux
    port map (
            O => \N__37907\,
            I => \N__37825\
        );

    \I__7519\ : Sp12to4
    port map (
            O => \N__37904\,
            I => \N__37821\
        );

    \I__7518\ : InMux
    port map (
            O => \N__37903\,
            I => \N__37818\
        );

    \I__7517\ : Span4Mux_v
    port map (
            O => \N__37898\,
            I => \N__37811\
        );

    \I__7516\ : Span4Mux_h
    port map (
            O => \N__37895\,
            I => \N__37811\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__37878\,
            I => \N__37811\
        );

    \I__7514\ : InMux
    port map (
            O => \N__37875\,
            I => \N__37794\
        );

    \I__7513\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37794\
        );

    \I__7512\ : InMux
    port map (
            O => \N__37873\,
            I => \N__37794\
        );

    \I__7511\ : InMux
    port map (
            O => \N__37870\,
            I => \N__37794\
        );

    \I__7510\ : InMux
    port map (
            O => \N__37869\,
            I => \N__37794\
        );

    \I__7509\ : InMux
    port map (
            O => \N__37866\,
            I => \N__37794\
        );

    \I__7508\ : InMux
    port map (
            O => \N__37865\,
            I => \N__37794\
        );

    \I__7507\ : InMux
    port map (
            O => \N__37862\,
            I => \N__37794\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__37845\,
            I => \N__37791\
        );

    \I__7505\ : InMux
    port map (
            O => \N__37842\,
            I => \N__37774\
        );

    \I__7504\ : InMux
    port map (
            O => \N__37841\,
            I => \N__37774\
        );

    \I__7503\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37774\
        );

    \I__7502\ : InMux
    port map (
            O => \N__37837\,
            I => \N__37774\
        );

    \I__7501\ : InMux
    port map (
            O => \N__37834\,
            I => \N__37774\
        );

    \I__7500\ : InMux
    port map (
            O => \N__37833\,
            I => \N__37774\
        );

    \I__7499\ : InMux
    port map (
            O => \N__37830\,
            I => \N__37774\
        );

    \I__7498\ : InMux
    port map (
            O => \N__37829\,
            I => \N__37774\
        );

    \I__7497\ : InMux
    port map (
            O => \N__37828\,
            I => \N__37767\
        );

    \I__7496\ : InMux
    port map (
            O => \N__37825\,
            I => \N__37767\
        );

    \I__7495\ : InMux
    port map (
            O => \N__37824\,
            I => \N__37767\
        );

    \I__7494\ : Span12Mux_h
    port map (
            O => \N__37821\,
            I => \N__37762\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__37818\,
            I => \N__37762\
        );

    \I__7492\ : Span4Mux_h
    port map (
            O => \N__37811\,
            I => \N__37757\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__37794\,
            I => \N__37757\
        );

    \I__7490\ : Span4Mux_v
    port map (
            O => \N__37791\,
            I => \N__37752\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__37774\,
            I => \N__37752\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__37767\,
            I => \N__37749\
        );

    \I__7487\ : Span12Mux_v
    port map (
            O => \N__37762\,
            I => \N__37746\
        );

    \I__7486\ : Span4Mux_v
    port map (
            O => \N__37757\,
            I => \N__37743\
        );

    \I__7485\ : Span4Mux_h
    port map (
            O => \N__37752\,
            I => \N__37738\
        );

    \I__7484\ : Span4Mux_v
    port map (
            O => \N__37749\,
            I => \N__37738\
        );

    \I__7483\ : Odrv12
    port map (
            O => \N__37746\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7482\ : Odrv4
    port map (
            O => \N__37743\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7481\ : Odrv4
    port map (
            O => \N__37738\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7480\ : InMux
    port map (
            O => \N__37731\,
            I => \N__37728\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__37728\,
            I => \N__37725\
        );

    \I__7478\ : Span12Mux_h
    port map (
            O => \N__37725\,
            I => \N__37722\
        );

    \I__7477\ : Odrv12
    port map (
            O => \N__37722\,
            I => \sDAC_dataZ0Z_13\
        );

    \I__7476\ : InMux
    port map (
            O => \N__37719\,
            I => \N__37716\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__37716\,
            I => \N__37713\
        );

    \I__7474\ : Span4Mux_h
    port map (
            O => \N__37713\,
            I => \N__37710\
        );

    \I__7473\ : Span4Mux_v
    port map (
            O => \N__37710\,
            I => \N__37707\
        );

    \I__7472\ : Span4Mux_h
    port map (
            O => \N__37707\,
            I => \N__37704\
        );

    \I__7471\ : Odrv4
    port map (
            O => \N__37704\,
            I => \sDAC_dataZ0Z_14\
        );

    \I__7470\ : InMux
    port map (
            O => \N__37701\,
            I => \N__37698\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__37698\,
            I => \N__37695\
        );

    \I__7468\ : Span4Mux_h
    port map (
            O => \N__37695\,
            I => \N__37692\
        );

    \I__7467\ : Span4Mux_v
    port map (
            O => \N__37692\,
            I => \N__37689\
        );

    \I__7466\ : Span4Mux_h
    port map (
            O => \N__37689\,
            I => \N__37686\
        );

    \I__7465\ : Odrv4
    port map (
            O => \N__37686\,
            I => \sDAC_dataZ0Z_15\
        );

    \I__7464\ : CascadeMux
    port map (
            O => \N__37683\,
            I => \sDAC_data_RNO_31Z0Z_8_cascade_\
        );

    \I__7463\ : CascadeMux
    port map (
            O => \N__37680\,
            I => \sDAC_data_2_39_ns_1_8_cascade_\
        );

    \I__7462\ : InMux
    port map (
            O => \N__37677\,
            I => \N__37674\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__37674\,
            I => \sDAC_data_RNO_32Z0Z_8\
        );

    \I__7460\ : InMux
    port map (
            O => \N__37671\,
            I => \N__37668\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__37668\,
            I => \sDAC_data_RNO_23Z0Z_8\
        );

    \I__7458\ : InMux
    port map (
            O => \N__37665\,
            I => \N__37662\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__37662\,
            I => \sDAC_mem_31Z0Z_5\
        );

    \I__7456\ : InMux
    port map (
            O => \N__37659\,
            I => \N__37656\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__37656\,
            I => \sDAC_data_RNO_24Z0Z_8\
        );

    \I__7454\ : InMux
    port map (
            O => \N__37653\,
            I => \N__37650\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__37650\,
            I => \sDAC_data_RNO_17Z0Z_10\
        );

    \I__7452\ : InMux
    port map (
            O => \N__37647\,
            I => \N__37644\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__37644\,
            I => \sDAC_data_2_24_ns_1_10\
        );

    \I__7450\ : CascadeMux
    port map (
            O => \N__37641\,
            I => \sDAC_data_RNO_8Z0Z_10_cascade_\
        );

    \I__7449\ : CascadeMux
    port map (
            O => \N__37638\,
            I => \sDAC_data_2_20_am_1_10_cascade_\
        );

    \I__7448\ : InMux
    port map (
            O => \N__37635\,
            I => \N__37632\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__37632\,
            I => \sDAC_data_RNO_7Z0Z_10\
        );

    \I__7446\ : InMux
    port map (
            O => \N__37629\,
            I => \N__37626\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__37626\,
            I => \sDAC_mem_28Z0Z_6\
        );

    \I__7444\ : InMux
    port map (
            O => \N__37623\,
            I => \N__37620\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__37620\,
            I => \N__37617\
        );

    \I__7442\ : Span4Mux_h
    port map (
            O => \N__37617\,
            I => \N__37614\
        );

    \I__7441\ : Span4Mux_h
    port map (
            O => \N__37614\,
            I => \N__37611\
        );

    \I__7440\ : Span4Mux_v
    port map (
            O => \N__37611\,
            I => \N__37608\
        );

    \I__7439\ : Odrv4
    port map (
            O => \N__37608\,
            I => \sDAC_dataZ0Z_1\
        );

    \I__7438\ : InMux
    port map (
            O => \N__37605\,
            I => \N__37602\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__37602\,
            I => \N__37599\
        );

    \I__7436\ : Span4Mux_v
    port map (
            O => \N__37599\,
            I => \N__37596\
        );

    \I__7435\ : Span4Mux_v
    port map (
            O => \N__37596\,
            I => \N__37593\
        );

    \I__7434\ : Span4Mux_h
    port map (
            O => \N__37593\,
            I => \N__37590\
        );

    \I__7433\ : Odrv4
    port map (
            O => \N__37590\,
            I => \sDAC_dataZ0Z_11\
        );

    \I__7432\ : InMux
    port map (
            O => \N__37587\,
            I => \N__37584\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__37584\,
            I => \N__37581\
        );

    \I__7430\ : Span4Mux_v
    port map (
            O => \N__37581\,
            I => \N__37578\
        );

    \I__7429\ : Span4Mux_v
    port map (
            O => \N__37578\,
            I => \N__37575\
        );

    \I__7428\ : Span4Mux_h
    port map (
            O => \N__37575\,
            I => \N__37572\
        );

    \I__7427\ : Odrv4
    port map (
            O => \N__37572\,
            I => \sDAC_dataZ0Z_12\
        );

    \I__7426\ : InMux
    port map (
            O => \N__37569\,
            I => \N__37566\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__37566\,
            I => \N__37563\
        );

    \I__7424\ : Odrv4
    port map (
            O => \N__37563\,
            I => \sDAC_mem_17Z0Z_6\
        );

    \I__7423\ : InMux
    port map (
            O => \N__37560\,
            I => \N__37557\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__37557\,
            I => \sDAC_mem_16Z0Z_6\
        );

    \I__7421\ : InMux
    port map (
            O => \N__37554\,
            I => \sDAC_mem_pointer_0_cry_1\
        );

    \I__7420\ : InMux
    port map (
            O => \N__37551\,
            I => \sDAC_mem_pointer_0_cry_2\
        );

    \I__7419\ : InMux
    port map (
            O => \N__37548\,
            I => \sDAC_mem_pointer_0_cry_3\
        );

    \I__7418\ : InMux
    port map (
            O => \N__37545\,
            I => \sDAC_mem_pointer_0_cry_4\
        );

    \I__7417\ : CascadeMux
    port map (
            O => \N__37542\,
            I => \sDAC_data_RNO_23Z0Z_9_cascade_\
        );

    \I__7416\ : CascadeMux
    port map (
            O => \N__37539\,
            I => \sDAC_data_RNO_17Z0Z_9_cascade_\
        );

    \I__7415\ : CascadeMux
    port map (
            O => \N__37536\,
            I => \sDAC_data_RNO_8Z0Z_9_cascade_\
        );

    \I__7414\ : CascadeMux
    port map (
            O => \N__37533\,
            I => \sDAC_data_2_20_am_1_9_cascade_\
        );

    \I__7413\ : InMux
    port map (
            O => \N__37530\,
            I => \N__37527\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__37527\,
            I => \sDAC_data_RNO_7Z0Z_9\
        );

    \I__7411\ : InMux
    port map (
            O => \N__37524\,
            I => \N__37521\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__37521\,
            I => \N__37518\
        );

    \I__7409\ : Odrv4
    port map (
            O => \N__37518\,
            I => \sDAC_mem_17Z0Z_4\
        );

    \I__7408\ : InMux
    port map (
            O => \N__37515\,
            I => \N__37512\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__37512\,
            I => \sDAC_mem_16Z0Z_4\
        );

    \I__7406\ : InMux
    port map (
            O => \N__37509\,
            I => \N__37506\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__37506\,
            I => \N__37503\
        );

    \I__7404\ : Odrv12
    port map (
            O => \N__37503\,
            I => \sDAC_mem_17Z0Z_5\
        );

    \I__7403\ : InMux
    port map (
            O => \N__37500\,
            I => \N__37497\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__37497\,
            I => \sDAC_mem_16Z0Z_5\
        );

    \I__7401\ : InMux
    port map (
            O => \N__37494\,
            I => \N__37476\
        );

    \I__7400\ : InMux
    port map (
            O => \N__37493\,
            I => \N__37476\
        );

    \I__7399\ : InMux
    port map (
            O => \N__37492\,
            I => \N__37476\
        );

    \I__7398\ : InMux
    port map (
            O => \N__37491\,
            I => \N__37476\
        );

    \I__7397\ : InMux
    port map (
            O => \N__37490\,
            I => \N__37476\
        );

    \I__7396\ : InMux
    port map (
            O => \N__37489\,
            I => \N__37476\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__37476\,
            I => \N_279\
        );

    \I__7394\ : CascadeMux
    port map (
            O => \N__37473\,
            I => \N_279_cascade_\
        );

    \I__7393\ : InMux
    port map (
            O => \N__37470\,
            I => \N__37467\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__37467\,
            I => \N__37464\
        );

    \I__7391\ : Odrv4
    port map (
            O => \N__37464\,
            I => \sDAC_data_RNO_21Z0Z_7\
        );

    \I__7390\ : CascadeMux
    port map (
            O => \N__37461\,
            I => \sDAC_data_2_14_ns_1_7_cascade_\
        );

    \I__7389\ : InMux
    port map (
            O => \N__37458\,
            I => \N__37455\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__37455\,
            I => \N__37452\
        );

    \I__7387\ : Odrv4
    port map (
            O => \N__37452\,
            I => \sDAC_data_RNO_4Z0Z_7\
        );

    \I__7386\ : InMux
    port map (
            O => \N__37449\,
            I => \N__37446\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__37446\,
            I => \sDAC_data_RNO_10Z0Z_7\
        );

    \I__7384\ : InMux
    port map (
            O => \N__37443\,
            I => \N__37440\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__37440\,
            I => \sDAC_data_RNO_2Z0Z_7\
        );

    \I__7382\ : CascadeMux
    port map (
            O => \N__37437\,
            I => \sDAC_data_2_41_ns_1_7_cascade_\
        );

    \I__7381\ : InMux
    port map (
            O => \N__37434\,
            I => \N__37431\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__37431\,
            I => \sDAC_data_RNO_1Z0Z_7\
        );

    \I__7379\ : CascadeMux
    port map (
            O => \N__37428\,
            I => \sDAC_data_2_7_cascade_\
        );

    \I__7378\ : InMux
    port map (
            O => \N__37425\,
            I => \N__37422\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__37422\,
            I => \N__37419\
        );

    \I__7376\ : Span4Mux_h
    port map (
            O => \N__37419\,
            I => \N__37416\
        );

    \I__7375\ : Odrv4
    port map (
            O => \N__37416\,
            I => \sDAC_dataZ0Z_7\
        );

    \I__7374\ : InMux
    port map (
            O => \N__37413\,
            I => \N__37410\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__37410\,
            I => \sDAC_mem_5Z0Z_4\
        );

    \I__7372\ : CEMux
    port map (
            O => \N__37407\,
            I => \N__37404\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__37404\,
            I => \N__37401\
        );

    \I__7370\ : Span4Mux_h
    port map (
            O => \N__37401\,
            I => \N__37398\
        );

    \I__7369\ : Odrv4
    port map (
            O => \N__37398\,
            I => \sDAC_mem_2_1_sqmuxa\
        );

    \I__7368\ : CEMux
    port map (
            O => \N__37395\,
            I => \N__37392\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__37392\,
            I => \N__37389\
        );

    \I__7366\ : Span4Mux_v
    port map (
            O => \N__37389\,
            I => \N__37386\
        );

    \I__7365\ : Odrv4
    port map (
            O => \N__37386\,
            I => \sDAC_mem_5_1_sqmuxa\
        );

    \I__7364\ : CEMux
    port map (
            O => \N__37383\,
            I => \N__37380\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__37380\,
            I => \N__37377\
        );

    \I__7362\ : Span4Mux_v
    port map (
            O => \N__37377\,
            I => \N__37374\
        );

    \I__7361\ : Span4Mux_h
    port map (
            O => \N__37374\,
            I => \N__37371\
        );

    \I__7360\ : Odrv4
    port map (
            O => \N__37371\,
            I => \sDAC_mem_7_1_sqmuxa\
        );

    \I__7359\ : InMux
    port map (
            O => \N__37368\,
            I => \N__37365\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__37365\,
            I => \N__37362\
        );

    \I__7357\ : Odrv4
    port map (
            O => \N__37362\,
            I => \sDAC_mem_7Z0Z_2\
        );

    \I__7356\ : InMux
    port map (
            O => \N__37359\,
            I => \N__37356\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__37356\,
            I => \sDAC_mem_5Z0Z_2\
        );

    \I__7354\ : InMux
    port map (
            O => \N__37353\,
            I => \N__37350\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__37350\,
            I => \sDAC_mem_5Z0Z_3\
        );

    \I__7352\ : InMux
    port map (
            O => \N__37347\,
            I => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4\
        );

    \I__7351\ : InMux
    port map (
            O => \N__37344\,
            I => \N__37340\
        );

    \I__7350\ : InMux
    port map (
            O => \N__37343\,
            I => \N__37337\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__37340\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__37337\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__7347\ : InMux
    port map (
            O => \N__37332\,
            I => \N__37329\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__37329\,
            I => \N__37326\
        );

    \I__7345\ : Span4Mux_v
    port map (
            O => \N__37326\,
            I => \N__37323\
        );

    \I__7344\ : Odrv4
    port map (
            O => \N__37323\,
            I => \sDAC_mem_34Z0Z_0\
        );

    \I__7343\ : InMux
    port map (
            O => \N__37320\,
            I => \N__37317\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__37317\,
            I => \N__37314\
        );

    \I__7341\ : Span4Mux_v
    port map (
            O => \N__37314\,
            I => \N__37311\
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__37311\,
            I => \sDAC_mem_34Z0Z_2\
        );

    \I__7339\ : InMux
    port map (
            O => \N__37308\,
            I => \N__37305\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__37305\,
            I => \N__37302\
        );

    \I__7337\ : Span4Mux_v
    port map (
            O => \N__37302\,
            I => \N__37299\
        );

    \I__7336\ : Odrv4
    port map (
            O => \N__37299\,
            I => \sDAC_mem_34Z0Z_6\
        );

    \I__7335\ : InMux
    port map (
            O => \N__37296\,
            I => \N__37293\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__37293\,
            I => \sDAC_mem_7Z0Z_0\
        );

    \I__7333\ : InMux
    port map (
            O => \N__37290\,
            I => \N__37287\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__37287\,
            I => \sDAC_mem_7Z0Z_1\
        );

    \I__7331\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37281\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__37281\,
            I => \sDAC_mem_16Z0Z_2\
        );

    \I__7329\ : InMux
    port map (
            O => \N__37278\,
            I => \N__37275\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__37275\,
            I => \sDAC_mem_pointerZ0Z_6\
        );

    \I__7327\ : InMux
    port map (
            O => \N__37272\,
            I => \N__37269\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__37269\,
            I => \sDAC_mem_pointerZ0Z_7\
        );

    \I__7325\ : CascadeMux
    port map (
            O => \N__37266\,
            I => \N__37262\
        );

    \I__7324\ : InMux
    port map (
            O => \N__37265\,
            I => \N__37259\
        );

    \I__7323\ : InMux
    port map (
            O => \N__37262\,
            I => \N__37256\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__37259\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__37256\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1\
        );

    \I__7320\ : InMux
    port map (
            O => \N__37251\,
            I => \N__37248\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__37248\,
            I => \N__37245\
        );

    \I__7318\ : Span4Mux_h
    port map (
            O => \N__37245\,
            I => \N__37241\
        );

    \I__7317\ : CascadeMux
    port map (
            O => \N__37244\,
            I => \N__37237\
        );

    \I__7316\ : Span4Mux_v
    port map (
            O => \N__37241\,
            I => \N__37234\
        );

    \I__7315\ : InMux
    port map (
            O => \N__37240\,
            I => \N__37231\
        );

    \I__7314\ : InMux
    port map (
            O => \N__37237\,
            I => \N__37228\
        );

    \I__7313\ : Odrv4
    port map (
            O => \N__37234\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__37231\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__37228\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__7310\ : InMux
    port map (
            O => \N__37221\,
            I => \N__37215\
        );

    \I__7309\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37215\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__37215\,
            I => \N__37212\
        );

    \I__7307\ : Span4Mux_h
    port map (
            O => \N__37212\,
            I => \N__37209\
        );

    \I__7306\ : Span4Mux_v
    port map (
            O => \N__37209\,
            I => \N__37204\
        );

    \I__7305\ : InMux
    port map (
            O => \N__37208\,
            I => \N__37201\
        );

    \I__7304\ : InMux
    port map (
            O => \N__37207\,
            I => \N__37198\
        );

    \I__7303\ : Odrv4
    port map (
            O => \N__37204\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__37201\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__37198\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__7300\ : InMux
    port map (
            O => \N__37191\,
            I => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0\
        );

    \I__7299\ : CascadeMux
    port map (
            O => \N__37188\,
            I => \N__37182\
        );

    \I__7298\ : InMux
    port map (
            O => \N__37187\,
            I => \N__37177\
        );

    \I__7297\ : InMux
    port map (
            O => \N__37186\,
            I => \N__37177\
        );

    \I__7296\ : InMux
    port map (
            O => \N__37185\,
            I => \N__37174\
        );

    \I__7295\ : InMux
    port map (
            O => \N__37182\,
            I => \N__37171\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__37177\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_i6\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__37174\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_i6\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__37171\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_i6\
        );

    \I__7291\ : InMux
    port map (
            O => \N__37164\,
            I => \N__37157\
        );

    \I__7290\ : InMux
    port map (
            O => \N__37163\,
            I => \N__37157\
        );

    \I__7289\ : InMux
    port map (
            O => \N__37162\,
            I => \N__37154\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__37157\,
            I => \N__37148\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__37154\,
            I => \N__37148\
        );

    \I__7286\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37145\
        );

    \I__7285\ : Span4Mux_v
    port map (
            O => \N__37148\,
            I => \N__37140\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__37145\,
            I => \N__37140\
        );

    \I__7283\ : Span4Mux_h
    port map (
            O => \N__37140\,
            I => \N__37135\
        );

    \I__7282\ : InMux
    port map (
            O => \N__37139\,
            I => \N__37132\
        );

    \I__7281\ : InMux
    port map (
            O => \N__37138\,
            I => \N__37129\
        );

    \I__7280\ : Odrv4
    port map (
            O => \N__37135\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__37132\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__37129\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__7277\ : InMux
    port map (
            O => \N__37122\,
            I => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1\
        );

    \I__7276\ : InMux
    port map (
            O => \N__37119\,
            I => \N__37115\
        );

    \I__7275\ : InMux
    port map (
            O => \N__37118\,
            I => \N__37112\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__37115\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__37112\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__7272\ : InMux
    port map (
            O => \N__37107\,
            I => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2\
        );

    \I__7271\ : InMux
    port map (
            O => \N__37104\,
            I => \N__37100\
        );

    \I__7270\ : InMux
    port map (
            O => \N__37103\,
            I => \N__37097\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__37100\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__37097\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__7267\ : InMux
    port map (
            O => \N__37092\,
            I => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3\
        );

    \I__7266\ : CascadeMux
    port map (
            O => \N__37089\,
            I => \N__37084\
        );

    \I__7265\ : InMux
    port map (
            O => \N__37088\,
            I => \N__37080\
        );

    \I__7264\ : InMux
    port map (
            O => \N__37087\,
            I => \N__37076\
        );

    \I__7263\ : InMux
    port map (
            O => \N__37084\,
            I => \N__37071\
        );

    \I__7262\ : CascadeMux
    port map (
            O => \N__37083\,
            I => \N__37068\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__37080\,
            I => \N__37065\
        );

    \I__7260\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37062\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__37076\,
            I => \N__37059\
        );

    \I__7258\ : InMux
    port map (
            O => \N__37075\,
            I => \N__37055\
        );

    \I__7257\ : InMux
    port map (
            O => \N__37074\,
            I => \N__37050\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__37071\,
            I => \N__37047\
        );

    \I__7255\ : InMux
    port map (
            O => \N__37068\,
            I => \N__37044\
        );

    \I__7254\ : Span4Mux_h
    port map (
            O => \N__37065\,
            I => \N__37039\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__37062\,
            I => \N__37039\
        );

    \I__7252\ : Span4Mux_v
    port map (
            O => \N__37059\,
            I => \N__37036\
        );

    \I__7251\ : InMux
    port map (
            O => \N__37058\,
            I => \N__37033\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__37055\,
            I => \N__37030\
        );

    \I__7249\ : InMux
    port map (
            O => \N__37054\,
            I => \N__37027\
        );

    \I__7248\ : InMux
    port map (
            O => \N__37053\,
            I => \N__37024\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__37050\,
            I => \N__37021\
        );

    \I__7246\ : Span4Mux_v
    port map (
            O => \N__37047\,
            I => \N__37016\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__37044\,
            I => \N__37016\
        );

    \I__7244\ : Span4Mux_v
    port map (
            O => \N__37039\,
            I => \N__37009\
        );

    \I__7243\ : Span4Mux_h
    port map (
            O => \N__37036\,
            I => \N__37009\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__37033\,
            I => \N__37009\
        );

    \I__7241\ : Span4Mux_h
    port map (
            O => \N__37030\,
            I => \N__37006\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__37027\,
            I => un7_spon_23
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__37024\,
            I => un7_spon_23
        );

    \I__7238\ : Odrv12
    port map (
            O => \N__37021\,
            I => un7_spon_23
        );

    \I__7237\ : Odrv4
    port map (
            O => \N__37016\,
            I => un7_spon_23
        );

    \I__7236\ : Odrv4
    port map (
            O => \N__37009\,
            I => un7_spon_23
        );

    \I__7235\ : Odrv4
    port map (
            O => \N__37006\,
            I => un7_spon_23
        );

    \I__7234\ : InMux
    port map (
            O => \N__36993\,
            I => \N__36990\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__36990\,
            I => \N__36987\
        );

    \I__7232\ : Span4Mux_v
    port map (
            O => \N__36987\,
            I => \N__36984\
        );

    \I__7231\ : Span4Mux_v
    port map (
            O => \N__36984\,
            I => \N__36981\
        );

    \I__7230\ : Odrv4
    port map (
            O => \N__36981\,
            I => un17_sdacdyn_1
        );

    \I__7229\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36975\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__36975\,
            I => \N__36969\
        );

    \I__7227\ : InMux
    port map (
            O => \N__36974\,
            I => \N__36964\
        );

    \I__7226\ : InMux
    port map (
            O => \N__36973\,
            I => \N__36964\
        );

    \I__7225\ : InMux
    port map (
            O => \N__36972\,
            I => \N__36961\
        );

    \I__7224\ : Span4Mux_h
    port map (
            O => \N__36969\,
            I => \N__36952\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__36964\,
            I => \N__36949\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__36961\,
            I => \N__36946\
        );

    \I__7221\ : InMux
    port map (
            O => \N__36960\,
            I => \N__36941\
        );

    \I__7220\ : InMux
    port map (
            O => \N__36959\,
            I => \N__36941\
        );

    \I__7219\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36938\
        );

    \I__7218\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36935\
        );

    \I__7217\ : InMux
    port map (
            O => \N__36956\,
            I => \N__36931\
        );

    \I__7216\ : InMux
    port map (
            O => \N__36955\,
            I => \N__36928\
        );

    \I__7215\ : Span4Mux_h
    port map (
            O => \N__36952\,
            I => \N__36925\
        );

    \I__7214\ : Span4Mux_h
    port map (
            O => \N__36949\,
            I => \N__36922\
        );

    \I__7213\ : Span4Mux_v
    port map (
            O => \N__36946\,
            I => \N__36917\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__36941\,
            I => \N__36917\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__36938\,
            I => \N__36914\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__36935\,
            I => \N__36911\
        );

    \I__7209\ : InMux
    port map (
            O => \N__36934\,
            I => \N__36908\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__36931\,
            I => \N__36901\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__36928\,
            I => \N__36901\
        );

    \I__7206\ : Span4Mux_v
    port map (
            O => \N__36925\,
            I => \N__36901\
        );

    \I__7205\ : Odrv4
    port map (
            O => \N__36922\,
            I => \N_1479\
        );

    \I__7204\ : Odrv4
    port map (
            O => \N__36917\,
            I => \N_1479\
        );

    \I__7203\ : Odrv4
    port map (
            O => \N__36914\,
            I => \N_1479\
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__36911\,
            I => \N_1479\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__36908\,
            I => \N_1479\
        );

    \I__7200\ : Odrv4
    port map (
            O => \N__36901\,
            I => \N_1479\
        );

    \I__7199\ : CascadeMux
    port map (
            O => \N__36888\,
            I => \N__36885\
        );

    \I__7198\ : InMux
    port map (
            O => \N__36885\,
            I => \N__36879\
        );

    \I__7197\ : CascadeMux
    port map (
            O => \N__36884\,
            I => \N__36874\
        );

    \I__7196\ : CascadeMux
    port map (
            O => \N__36883\,
            I => \N__36870\
        );

    \I__7195\ : CascadeMux
    port map (
            O => \N__36882\,
            I => \N__36867\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__36879\,
            I => \N__36864\
        );

    \I__7193\ : CascadeMux
    port map (
            O => \N__36878\,
            I => \N__36861\
        );

    \I__7192\ : InMux
    port map (
            O => \N__36877\,
            I => \N__36856\
        );

    \I__7191\ : InMux
    port map (
            O => \N__36874\,
            I => \N__36852\
        );

    \I__7190\ : CascadeMux
    port map (
            O => \N__36873\,
            I => \N__36849\
        );

    \I__7189\ : InMux
    port map (
            O => \N__36870\,
            I => \N__36845\
        );

    \I__7188\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36841\
        );

    \I__7187\ : Span4Mux_v
    port map (
            O => \N__36864\,
            I => \N__36837\
        );

    \I__7186\ : InMux
    port map (
            O => \N__36861\,
            I => \N__36832\
        );

    \I__7185\ : InMux
    port map (
            O => \N__36860\,
            I => \N__36832\
        );

    \I__7184\ : InMux
    port map (
            O => \N__36859\,
            I => \N__36829\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__36856\,
            I => \N__36826\
        );

    \I__7182\ : InMux
    port map (
            O => \N__36855\,
            I => \N__36823\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__36852\,
            I => \N__36820\
        );

    \I__7180\ : InMux
    port map (
            O => \N__36849\,
            I => \N__36814\
        );

    \I__7179\ : InMux
    port map (
            O => \N__36848\,
            I => \N__36814\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__36845\,
            I => \N__36810\
        );

    \I__7177\ : InMux
    port map (
            O => \N__36844\,
            I => \N__36807\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__36841\,
            I => \N__36801\
        );

    \I__7175\ : InMux
    port map (
            O => \N__36840\,
            I => \N__36798\
        );

    \I__7174\ : Span4Mux_h
    port map (
            O => \N__36837\,
            I => \N__36795\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__36832\,
            I => \N__36786\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__36829\,
            I => \N__36786\
        );

    \I__7171\ : Span4Mux_v
    port map (
            O => \N__36826\,
            I => \N__36786\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__36823\,
            I => \N__36786\
        );

    \I__7169\ : Span4Mux_h
    port map (
            O => \N__36820\,
            I => \N__36783\
        );

    \I__7168\ : InMux
    port map (
            O => \N__36819\,
            I => \N__36779\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__36814\,
            I => \N__36776\
        );

    \I__7166\ : InMux
    port map (
            O => \N__36813\,
            I => \N__36773\
        );

    \I__7165\ : Span4Mux_h
    port map (
            O => \N__36810\,
            I => \N__36768\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__36807\,
            I => \N__36768\
        );

    \I__7163\ : InMux
    port map (
            O => \N__36806\,
            I => \N__36763\
        );

    \I__7162\ : InMux
    port map (
            O => \N__36805\,
            I => \N__36763\
        );

    \I__7161\ : InMux
    port map (
            O => \N__36804\,
            I => \N__36760\
        );

    \I__7160\ : Span4Mux_v
    port map (
            O => \N__36801\,
            I => \N__36753\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__36798\,
            I => \N__36753\
        );

    \I__7158\ : Span4Mux_v
    port map (
            O => \N__36795\,
            I => \N__36753\
        );

    \I__7157\ : Span4Mux_v
    port map (
            O => \N__36786\,
            I => \N__36748\
        );

    \I__7156\ : Span4Mux_h
    port map (
            O => \N__36783\,
            I => \N__36748\
        );

    \I__7155\ : InMux
    port map (
            O => \N__36782\,
            I => \N__36745\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__36779\,
            I => \N__36742\
        );

    \I__7153\ : Odrv12
    port map (
            O => \N__36776\,
            I => un7_spon_4
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__36773\,
            I => un7_spon_4
        );

    \I__7151\ : Odrv4
    port map (
            O => \N__36768\,
            I => un7_spon_4
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__36763\,
            I => un7_spon_4
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__36760\,
            I => un7_spon_4
        );

    \I__7148\ : Odrv4
    port map (
            O => \N__36753\,
            I => un7_spon_4
        );

    \I__7147\ : Odrv4
    port map (
            O => \N__36748\,
            I => un7_spon_4
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__36745\,
            I => un7_spon_4
        );

    \I__7145\ : Odrv4
    port map (
            O => \N__36742\,
            I => un7_spon_4
        );

    \I__7144\ : InMux
    port map (
            O => \N__36723\,
            I => \bfn_14_19_0_\
        );

    \I__7143\ : InMux
    port map (
            O => \N__36720\,
            I => \N__36717\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__36717\,
            I => \N__36714\
        );

    \I__7141\ : Span4Mux_v
    port map (
            O => \N__36714\,
            I => \N__36711\
        );

    \I__7140\ : Odrv4
    port map (
            O => \N__36711\,
            I => \sDAC_mem_24Z0Z_3\
        );

    \I__7139\ : InMux
    port map (
            O => \N__36708\,
            I => \N__36705\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__36705\,
            I => \N__36702\
        );

    \I__7137\ : Span4Mux_v
    port map (
            O => \N__36702\,
            I => \N__36699\
        );

    \I__7136\ : Odrv4
    port map (
            O => \N__36699\,
            I => \sDAC_mem_24Z0Z_6\
        );

    \I__7135\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36693\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__36693\,
            I => \N__36690\
        );

    \I__7133\ : Span4Mux_v
    port map (
            O => \N__36690\,
            I => \N__36687\
        );

    \I__7132\ : Span4Mux_v
    port map (
            O => \N__36687\,
            I => \N__36684\
        );

    \I__7131\ : Odrv4
    port map (
            O => \N__36684\,
            I => \sDAC_mem_17Z0Z_2\
        );

    \I__7130\ : CascadeMux
    port map (
            O => \N__36681\,
            I => \N__36678\
        );

    \I__7129\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36675\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__36675\,
            I => \N__36672\
        );

    \I__7127\ : Span4Mux_v
    port map (
            O => \N__36672\,
            I => \N__36669\
        );

    \I__7126\ : Span4Mux_v
    port map (
            O => \N__36669\,
            I => \N__36666\
        );

    \I__7125\ : Span4Mux_v
    port map (
            O => \N__36666\,
            I => \N__36663\
        );

    \I__7124\ : Odrv4
    port map (
            O => \N__36663\,
            I => \sDAC_data_RNO_29Z0Z_5\
        );

    \I__7123\ : InMux
    port map (
            O => \N__36660\,
            I => \N__36656\
        );

    \I__7122\ : InMux
    port map (
            O => \N__36659\,
            I => \N__36650\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__36656\,
            I => \N__36647\
        );

    \I__7120\ : InMux
    port map (
            O => \N__36655\,
            I => \N__36644\
        );

    \I__7119\ : InMux
    port map (
            O => \N__36654\,
            I => \N__36641\
        );

    \I__7118\ : CascadeMux
    port map (
            O => \N__36653\,
            I => \N__36638\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__36650\,
            I => \N__36634\
        );

    \I__7116\ : Span4Mux_h
    port map (
            O => \N__36647\,
            I => \N__36630\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__36644\,
            I => \N__36626\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__36641\,
            I => \N__36623\
        );

    \I__7113\ : InMux
    port map (
            O => \N__36638\,
            I => \N__36620\
        );

    \I__7112\ : InMux
    port map (
            O => \N__36637\,
            I => \N__36617\
        );

    \I__7111\ : Span12Mux_v
    port map (
            O => \N__36634\,
            I => \N__36613\
        );

    \I__7110\ : InMux
    port map (
            O => \N__36633\,
            I => \N__36610\
        );

    \I__7109\ : Span4Mux_h
    port map (
            O => \N__36630\,
            I => \N__36607\
        );

    \I__7108\ : InMux
    port map (
            O => \N__36629\,
            I => \N__36604\
        );

    \I__7107\ : Span4Mux_h
    port map (
            O => \N__36626\,
            I => \N__36599\
        );

    \I__7106\ : Span4Mux_h
    port map (
            O => \N__36623\,
            I => \N__36599\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__36620\,
            I => \N__36596\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__36617\,
            I => \N__36593\
        );

    \I__7103\ : InMux
    port map (
            O => \N__36616\,
            I => \N__36590\
        );

    \I__7102\ : Odrv12
    port map (
            O => \N__36613\,
            I => un7_spon_15
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__36610\,
            I => un7_spon_15
        );

    \I__7100\ : Odrv4
    port map (
            O => \N__36607\,
            I => un7_spon_15
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__36604\,
            I => un7_spon_15
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__36599\,
            I => un7_spon_15
        );

    \I__7097\ : Odrv4
    port map (
            O => \N__36596\,
            I => un7_spon_15
        );

    \I__7096\ : Odrv12
    port map (
            O => \N__36593\,
            I => un7_spon_15
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__36590\,
            I => un7_spon_15
        );

    \I__7094\ : InMux
    port map (
            O => \N__36573\,
            I => \N__36570\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__36570\,
            I => \N__36566\
        );

    \I__7092\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36563\
        );

    \I__7091\ : Span4Mux_v
    port map (
            O => \N__36566\,
            I => \N__36558\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__36563\,
            I => \N__36558\
        );

    \I__7089\ : Odrv4
    port map (
            O => \N__36558\,
            I => \sEEACQZ0Z_15\
        );

    \I__7088\ : CascadeMux
    port map (
            O => \N__36555\,
            I => \N__36552\
        );

    \I__7087\ : InMux
    port map (
            O => \N__36552\,
            I => \N__36549\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__36549\,
            I => \sEEACQ_i_15\
        );

    \I__7085\ : CascadeMux
    port map (
            O => \N__36546\,
            I => \N__36542\
        );

    \I__7084\ : CascadeMux
    port map (
            O => \N__36545\,
            I => \N__36538\
        );

    \I__7083\ : InMux
    port map (
            O => \N__36542\,
            I => \N__36535\
        );

    \I__7082\ : InMux
    port map (
            O => \N__36541\,
            I => \N__36532\
        );

    \I__7081\ : InMux
    port map (
            O => \N__36538\,
            I => \N__36526\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__36535\,
            I => \N__36522\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__36532\,
            I => \N__36518\
        );

    \I__7078\ : InMux
    port map (
            O => \N__36531\,
            I => \N__36514\
        );

    \I__7077\ : InMux
    port map (
            O => \N__36530\,
            I => \N__36511\
        );

    \I__7076\ : InMux
    port map (
            O => \N__36529\,
            I => \N__36508\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__36526\,
            I => \N__36504\
        );

    \I__7074\ : InMux
    port map (
            O => \N__36525\,
            I => \N__36501\
        );

    \I__7073\ : Span4Mux_h
    port map (
            O => \N__36522\,
            I => \N__36498\
        );

    \I__7072\ : InMux
    port map (
            O => \N__36521\,
            I => \N__36495\
        );

    \I__7071\ : Span4Mux_v
    port map (
            O => \N__36518\,
            I => \N__36492\
        );

    \I__7070\ : InMux
    port map (
            O => \N__36517\,
            I => \N__36489\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__36514\,
            I => \N__36486\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__36511\,
            I => \N__36483\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__36508\,
            I => \N__36480\
        );

    \I__7066\ : InMux
    port map (
            O => \N__36507\,
            I => \N__36477\
        );

    \I__7065\ : Span4Mux_h
    port map (
            O => \N__36504\,
            I => \N__36472\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__36501\,
            I => \N__36472\
        );

    \I__7063\ : Span4Mux_v
    port map (
            O => \N__36498\,
            I => \N__36463\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__36495\,
            I => \N__36463\
        );

    \I__7061\ : Span4Mux_h
    port map (
            O => \N__36492\,
            I => \N__36463\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__36489\,
            I => \N__36463\
        );

    \I__7059\ : Span4Mux_v
    port map (
            O => \N__36486\,
            I => \N__36458\
        );

    \I__7058\ : Span4Mux_v
    port map (
            O => \N__36483\,
            I => \N__36458\
        );

    \I__7057\ : Span4Mux_v
    port map (
            O => \N__36480\,
            I => \N__36455\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__36477\,
            I => un7_spon_16
        );

    \I__7055\ : Odrv4
    port map (
            O => \N__36472\,
            I => un7_spon_16
        );

    \I__7054\ : Odrv4
    port map (
            O => \N__36463\,
            I => un7_spon_16
        );

    \I__7053\ : Odrv4
    port map (
            O => \N__36458\,
            I => un7_spon_16
        );

    \I__7052\ : Odrv4
    port map (
            O => \N__36455\,
            I => un7_spon_16
        );

    \I__7051\ : InMux
    port map (
            O => \N__36444\,
            I => \N__36438\
        );

    \I__7050\ : CascadeMux
    port map (
            O => \N__36443\,
            I => \N__36435\
        );

    \I__7049\ : InMux
    port map (
            O => \N__36442\,
            I => \N__36432\
        );

    \I__7048\ : InMux
    port map (
            O => \N__36441\,
            I => \N__36427\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__36438\,
            I => \N__36423\
        );

    \I__7046\ : InMux
    port map (
            O => \N__36435\,
            I => \N__36420\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__36432\,
            I => \N__36417\
        );

    \I__7044\ : InMux
    port map (
            O => \N__36431\,
            I => \N__36413\
        );

    \I__7043\ : InMux
    port map (
            O => \N__36430\,
            I => \N__36410\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__36427\,
            I => \N__36407\
        );

    \I__7041\ : InMux
    port map (
            O => \N__36426\,
            I => \N__36402\
        );

    \I__7040\ : Span4Mux_h
    port map (
            O => \N__36423\,
            I => \N__36397\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__36420\,
            I => \N__36397\
        );

    \I__7038\ : Span4Mux_v
    port map (
            O => \N__36417\,
            I => \N__36394\
        );

    \I__7037\ : InMux
    port map (
            O => \N__36416\,
            I => \N__36391\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__36413\,
            I => \N__36388\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__36410\,
            I => \N__36385\
        );

    \I__7034\ : Span4Mux_v
    port map (
            O => \N__36407\,
            I => \N__36382\
        );

    \I__7033\ : InMux
    port map (
            O => \N__36406\,
            I => \N__36379\
        );

    \I__7032\ : InMux
    port map (
            O => \N__36405\,
            I => \N__36376\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__36402\,
            I => \N__36373\
        );

    \I__7030\ : Span4Mux_v
    port map (
            O => \N__36397\,
            I => \N__36366\
        );

    \I__7029\ : Span4Mux_h
    port map (
            O => \N__36394\,
            I => \N__36366\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__36391\,
            I => \N__36366\
        );

    \I__7027\ : Span4Mux_v
    port map (
            O => \N__36388\,
            I => \N__36361\
        );

    \I__7026\ : Span4Mux_h
    port map (
            O => \N__36385\,
            I => \N__36361\
        );

    \I__7025\ : Odrv4
    port map (
            O => \N__36382\,
            I => un7_spon_17
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__36379\,
            I => un7_spon_17
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__36376\,
            I => un7_spon_17
        );

    \I__7022\ : Odrv12
    port map (
            O => \N__36373\,
            I => un7_spon_17
        );

    \I__7021\ : Odrv4
    port map (
            O => \N__36366\,
            I => un7_spon_17
        );

    \I__7020\ : Odrv4
    port map (
            O => \N__36361\,
            I => un7_spon_17
        );

    \I__7019\ : CascadeMux
    port map (
            O => \N__36348\,
            I => \N__36342\
        );

    \I__7018\ : InMux
    port map (
            O => \N__36347\,
            I => \N__36339\
        );

    \I__7017\ : CascadeMux
    port map (
            O => \N__36346\,
            I => \N__36336\
        );

    \I__7016\ : InMux
    port map (
            O => \N__36345\,
            I => \N__36333\
        );

    \I__7015\ : InMux
    port map (
            O => \N__36342\,
            I => \N__36329\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__36339\,
            I => \N__36324\
        );

    \I__7013\ : InMux
    port map (
            O => \N__36336\,
            I => \N__36320\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__36333\,
            I => \N__36317\
        );

    \I__7011\ : InMux
    port map (
            O => \N__36332\,
            I => \N__36314\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__36329\,
            I => \N__36311\
        );

    \I__7009\ : InMux
    port map (
            O => \N__36328\,
            I => \N__36306\
        );

    \I__7008\ : InMux
    port map (
            O => \N__36327\,
            I => \N__36303\
        );

    \I__7007\ : Span4Mux_v
    port map (
            O => \N__36324\,
            I => \N__36300\
        );

    \I__7006\ : InMux
    port map (
            O => \N__36323\,
            I => \N__36297\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__36320\,
            I => \N__36290\
        );

    \I__7004\ : Span4Mux_v
    port map (
            O => \N__36317\,
            I => \N__36290\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__36314\,
            I => \N__36290\
        );

    \I__7002\ : Span4Mux_h
    port map (
            O => \N__36311\,
            I => \N__36287\
        );

    \I__7001\ : InMux
    port map (
            O => \N__36310\,
            I => \N__36284\
        );

    \I__7000\ : InMux
    port map (
            O => \N__36309\,
            I => \N__36281\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__36306\,
            I => \N__36278\
        );

    \I__6998\ : LocalMux
    port map (
            O => \N__36303\,
            I => \N__36271\
        );

    \I__6997\ : Span4Mux_h
    port map (
            O => \N__36300\,
            I => \N__36271\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__36297\,
            I => \N__36271\
        );

    \I__6995\ : Span4Mux_h
    port map (
            O => \N__36290\,
            I => \N__36268\
        );

    \I__6994\ : Odrv4
    port map (
            O => \N__36287\,
            I => un7_spon_18
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__36284\,
            I => un7_spon_18
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__36281\,
            I => un7_spon_18
        );

    \I__6991\ : Odrv4
    port map (
            O => \N__36278\,
            I => un7_spon_18
        );

    \I__6990\ : Odrv4
    port map (
            O => \N__36271\,
            I => un7_spon_18
        );

    \I__6989\ : Odrv4
    port map (
            O => \N__36268\,
            I => un7_spon_18
        );

    \I__6988\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36248\
        );

    \I__6987\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36244\
        );

    \I__6986\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36241\
        );

    \I__6985\ : InMux
    port map (
            O => \N__36252\,
            I => \N__36238\
        );

    \I__6984\ : InMux
    port map (
            O => \N__36251\,
            I => \N__36235\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__36248\,
            I => \N__36232\
        );

    \I__6982\ : InMux
    port map (
            O => \N__36247\,
            I => \N__36225\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__36244\,
            I => \N__36220\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__36241\,
            I => \N__36220\
        );

    \I__6979\ : LocalMux
    port map (
            O => \N__36238\,
            I => \N__36217\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__36235\,
            I => \N__36214\
        );

    \I__6977\ : Span4Mux_v
    port map (
            O => \N__36232\,
            I => \N__36211\
        );

    \I__6976\ : InMux
    port map (
            O => \N__36231\,
            I => \N__36208\
        );

    \I__6975\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36205\
        );

    \I__6974\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36202\
        );

    \I__6973\ : InMux
    port map (
            O => \N__36228\,
            I => \N__36199\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__36225\,
            I => \N__36196\
        );

    \I__6971\ : Span4Mux_h
    port map (
            O => \N__36220\,
            I => \N__36191\
        );

    \I__6970\ : Span4Mux_h
    port map (
            O => \N__36217\,
            I => \N__36191\
        );

    \I__6969\ : Span4Mux_v
    port map (
            O => \N__36214\,
            I => \N__36184\
        );

    \I__6968\ : Span4Mux_h
    port map (
            O => \N__36211\,
            I => \N__36184\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__36208\,
            I => \N__36184\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__36205\,
            I => un7_spon_19
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__36202\,
            I => un7_spon_19
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__36199\,
            I => un7_spon_19
        );

    \I__6963\ : Odrv4
    port map (
            O => \N__36196\,
            I => un7_spon_19
        );

    \I__6962\ : Odrv4
    port map (
            O => \N__36191\,
            I => un7_spon_19
        );

    \I__6961\ : Odrv4
    port map (
            O => \N__36184\,
            I => un7_spon_19
        );

    \I__6960\ : CascadeMux
    port map (
            O => \N__36171\,
            I => \N__36166\
        );

    \I__6959\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36163\
        );

    \I__6958\ : CascadeMux
    port map (
            O => \N__36169\,
            I => \N__36159\
        );

    \I__6957\ : InMux
    port map (
            O => \N__36166\,
            I => \N__36155\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__36163\,
            I => \N__36152\
        );

    \I__6955\ : InMux
    port map (
            O => \N__36162\,
            I => \N__36149\
        );

    \I__6954\ : InMux
    port map (
            O => \N__36159\,
            I => \N__36141\
        );

    \I__6953\ : InMux
    port map (
            O => \N__36158\,
            I => \N__36141\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__36155\,
            I => \N__36138\
        );

    \I__6951\ : Span4Mux_h
    port map (
            O => \N__36152\,
            I => \N__36133\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__36149\,
            I => \N__36130\
        );

    \I__6949\ : InMux
    port map (
            O => \N__36148\,
            I => \N__36125\
        );

    \I__6948\ : InMux
    port map (
            O => \N__36147\,
            I => \N__36125\
        );

    \I__6947\ : InMux
    port map (
            O => \N__36146\,
            I => \N__36122\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__36141\,
            I => \N__36119\
        );

    \I__6945\ : Span4Mux_v
    port map (
            O => \N__36138\,
            I => \N__36116\
        );

    \I__6944\ : InMux
    port map (
            O => \N__36137\,
            I => \N__36113\
        );

    \I__6943\ : InMux
    port map (
            O => \N__36136\,
            I => \N__36110\
        );

    \I__6942\ : Span4Mux_h
    port map (
            O => \N__36133\,
            I => \N__36107\
        );

    \I__6941\ : Span4Mux_v
    port map (
            O => \N__36130\,
            I => \N__36102\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__36125\,
            I => \N__36102\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__36122\,
            I => \N__36099\
        );

    \I__6938\ : Span4Mux_h
    port map (
            O => \N__36119\,
            I => \N__36096\
        );

    \I__6937\ : Odrv4
    port map (
            O => \N__36116\,
            I => un7_spon_20
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__36113\,
            I => un7_spon_20
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__36110\,
            I => un7_spon_20
        );

    \I__6934\ : Odrv4
    port map (
            O => \N__36107\,
            I => un7_spon_20
        );

    \I__6933\ : Odrv4
    port map (
            O => \N__36102\,
            I => un7_spon_20
        );

    \I__6932\ : Odrv12
    port map (
            O => \N__36099\,
            I => un7_spon_20
        );

    \I__6931\ : Odrv4
    port map (
            O => \N__36096\,
            I => un7_spon_20
        );

    \I__6930\ : InMux
    port map (
            O => \N__36081\,
            I => \N__36076\
        );

    \I__6929\ : CascadeMux
    port map (
            O => \N__36080\,
            I => \N__36073\
        );

    \I__6928\ : InMux
    port map (
            O => \N__36079\,
            I => \N__36069\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__36076\,
            I => \N__36066\
        );

    \I__6926\ : InMux
    port map (
            O => \N__36073\,
            I => \N__36060\
        );

    \I__6925\ : InMux
    port map (
            O => \N__36072\,
            I => \N__36057\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__36069\,
            I => \N__36054\
        );

    \I__6923\ : Span4Mux_h
    port map (
            O => \N__36066\,
            I => \N__36050\
        );

    \I__6922\ : InMux
    port map (
            O => \N__36065\,
            I => \N__36047\
        );

    \I__6921\ : InMux
    port map (
            O => \N__36064\,
            I => \N__36044\
        );

    \I__6920\ : InMux
    port map (
            O => \N__36063\,
            I => \N__36041\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__36060\,
            I => \N__36038\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__36057\,
            I => \N__36035\
        );

    \I__6917\ : Span4Mux_v
    port map (
            O => \N__36054\,
            I => \N__36032\
        );

    \I__6916\ : InMux
    port map (
            O => \N__36053\,
            I => \N__36029\
        );

    \I__6915\ : Span4Mux_h
    port map (
            O => \N__36050\,
            I => \N__36026\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__36047\,
            I => \N__36023\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__36044\,
            I => \N__36018\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__36041\,
            I => \N__36018\
        );

    \I__6911\ : Span4Mux_h
    port map (
            O => \N__36038\,
            I => \N__36013\
        );

    \I__6910\ : Span4Mux_h
    port map (
            O => \N__36035\,
            I => \N__36013\
        );

    \I__6909\ : Odrv4
    port map (
            O => \N__36032\,
            I => un7_spon_21
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__36029\,
            I => un7_spon_21
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__36026\,
            I => un7_spon_21
        );

    \I__6906\ : Odrv4
    port map (
            O => \N__36023\,
            I => un7_spon_21
        );

    \I__6905\ : Odrv12
    port map (
            O => \N__36018\,
            I => un7_spon_21
        );

    \I__6904\ : Odrv4
    port map (
            O => \N__36013\,
            I => un7_spon_21
        );

    \I__6903\ : CascadeMux
    port map (
            O => \N__36000\,
            I => \N__35997\
        );

    \I__6902\ : InMux
    port map (
            O => \N__35997\,
            I => \N__35991\
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__35996\,
            I => \N__35988\
        );

    \I__6900\ : CascadeMux
    port map (
            O => \N__35995\,
            I => \N__35985\
        );

    \I__6899\ : InMux
    port map (
            O => \N__35994\,
            I => \N__35982\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__35991\,
            I => \N__35976\
        );

    \I__6897\ : InMux
    port map (
            O => \N__35988\,
            I => \N__35973\
        );

    \I__6896\ : InMux
    port map (
            O => \N__35985\,
            I => \N__35970\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__35982\,
            I => \N__35967\
        );

    \I__6894\ : InMux
    port map (
            O => \N__35981\,
            I => \N__35964\
        );

    \I__6893\ : CascadeMux
    port map (
            O => \N__35980\,
            I => \N__35961\
        );

    \I__6892\ : CascadeMux
    port map (
            O => \N__35979\,
            I => \N__35957\
        );

    \I__6891\ : Span4Mux_h
    port map (
            O => \N__35976\,
            I => \N__35952\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__35973\,
            I => \N__35952\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__35970\,
            I => \N__35947\
        );

    \I__6888\ : Span4Mux_h
    port map (
            O => \N__35967\,
            I => \N__35944\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__35964\,
            I => \N__35941\
        );

    \I__6886\ : InMux
    port map (
            O => \N__35961\,
            I => \N__35938\
        );

    \I__6885\ : InMux
    port map (
            O => \N__35960\,
            I => \N__35935\
        );

    \I__6884\ : InMux
    port map (
            O => \N__35957\,
            I => \N__35932\
        );

    \I__6883\ : Span4Mux_v
    port map (
            O => \N__35952\,
            I => \N__35929\
        );

    \I__6882\ : InMux
    port map (
            O => \N__35951\,
            I => \N__35926\
        );

    \I__6881\ : InMux
    port map (
            O => \N__35950\,
            I => \N__35923\
        );

    \I__6880\ : Span4Mux_v
    port map (
            O => \N__35947\,
            I => \N__35920\
        );

    \I__6879\ : Span4Mux_h
    port map (
            O => \N__35944\,
            I => \N__35917\
        );

    \I__6878\ : Span4Mux_v
    port map (
            O => \N__35941\,
            I => \N__35912\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__35938\,
            I => \N__35912\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__35935\,
            I => \N__35909\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__35932\,
            I => \N__35906\
        );

    \I__6874\ : Odrv4
    port map (
            O => \N__35929\,
            I => un7_spon_22
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__35926\,
            I => un7_spon_22
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__35923\,
            I => un7_spon_22
        );

    \I__6871\ : Odrv4
    port map (
            O => \N__35920\,
            I => un7_spon_22
        );

    \I__6870\ : Odrv4
    port map (
            O => \N__35917\,
            I => un7_spon_22
        );

    \I__6869\ : Odrv4
    port map (
            O => \N__35912\,
            I => un7_spon_22
        );

    \I__6868\ : Odrv12
    port map (
            O => \N__35909\,
            I => un7_spon_22
        );

    \I__6867\ : Odrv12
    port map (
            O => \N__35906\,
            I => un7_spon_22
        );

    \I__6866\ : CascadeMux
    port map (
            O => \N__35889\,
            I => \N__35885\
        );

    \I__6865\ : CascadeMux
    port map (
            O => \N__35888\,
            I => \N__35882\
        );

    \I__6864\ : InMux
    port map (
            O => \N__35885\,
            I => \N__35878\
        );

    \I__6863\ : InMux
    port map (
            O => \N__35882\,
            I => \N__35874\
        );

    \I__6862\ : CascadeMux
    port map (
            O => \N__35881\,
            I => \N__35871\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__35878\,
            I => \N__35867\
        );

    \I__6860\ : InMux
    port map (
            O => \N__35877\,
            I => \N__35864\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__35874\,
            I => \N__35861\
        );

    \I__6858\ : InMux
    port map (
            O => \N__35871\,
            I => \N__35858\
        );

    \I__6857\ : InMux
    port map (
            O => \N__35870\,
            I => \N__35854\
        );

    \I__6856\ : Span4Mux_h
    port map (
            O => \N__35867\,
            I => \N__35851\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__35864\,
            I => \N__35846\
        );

    \I__6854\ : Span4Mux_h
    port map (
            O => \N__35861\,
            I => \N__35843\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__35858\,
            I => \N__35839\
        );

    \I__6852\ : InMux
    port map (
            O => \N__35857\,
            I => \N__35836\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__35854\,
            I => \N__35833\
        );

    \I__6850\ : Span4Mux_v
    port map (
            O => \N__35851\,
            I => \N__35830\
        );

    \I__6849\ : InMux
    port map (
            O => \N__35850\,
            I => \N__35827\
        );

    \I__6848\ : InMux
    port map (
            O => \N__35849\,
            I => \N__35824\
        );

    \I__6847\ : Span4Mux_v
    port map (
            O => \N__35846\,
            I => \N__35819\
        );

    \I__6846\ : Span4Mux_h
    port map (
            O => \N__35843\,
            I => \N__35819\
        );

    \I__6845\ : InMux
    port map (
            O => \N__35842\,
            I => \N__35816\
        );

    \I__6844\ : Span4Mux_h
    port map (
            O => \N__35839\,
            I => \N__35811\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__35836\,
            I => \N__35811\
        );

    \I__6842\ : Span4Mux_v
    port map (
            O => \N__35833\,
            I => \N__35808\
        );

    \I__6841\ : Odrv4
    port map (
            O => \N__35830\,
            I => un7_spon_8
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__35827\,
            I => un7_spon_8
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__35824\,
            I => un7_spon_8
        );

    \I__6838\ : Odrv4
    port map (
            O => \N__35819\,
            I => un7_spon_8
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__35816\,
            I => un7_spon_8
        );

    \I__6836\ : Odrv4
    port map (
            O => \N__35811\,
            I => un7_spon_8
        );

    \I__6835\ : Odrv4
    port map (
            O => \N__35808\,
            I => un7_spon_8
        );

    \I__6834\ : InMux
    port map (
            O => \N__35793\,
            I => \N__35789\
        );

    \I__6833\ : InMux
    port map (
            O => \N__35792\,
            I => \N__35786\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__35789\,
            I => \N__35783\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__35786\,
            I => \N__35780\
        );

    \I__6830\ : Odrv4
    port map (
            O => \N__35783\,
            I => \sEEACQZ0Z_8\
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__35780\,
            I => \sEEACQZ0Z_8\
        );

    \I__6828\ : InMux
    port map (
            O => \N__35775\,
            I => \N__35772\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__35772\,
            I => \sEEACQ_i_8\
        );

    \I__6826\ : InMux
    port map (
            O => \N__35769\,
            I => \N__35764\
        );

    \I__6825\ : InMux
    port map (
            O => \N__35768\,
            I => \N__35758\
        );

    \I__6824\ : InMux
    port map (
            O => \N__35767\,
            I => \N__35755\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__35764\,
            I => \N__35752\
        );

    \I__6822\ : InMux
    port map (
            O => \N__35763\,
            I => \N__35749\
        );

    \I__6821\ : InMux
    port map (
            O => \N__35762\,
            I => \N__35746\
        );

    \I__6820\ : CascadeMux
    port map (
            O => \N__35761\,
            I => \N__35743\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__35758\,
            I => \N__35740\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__35755\,
            I => \N__35735\
        );

    \I__6817\ : Span4Mux_v
    port map (
            O => \N__35752\,
            I => \N__35732\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__35749\,
            I => \N__35728\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__35746\,
            I => \N__35725\
        );

    \I__6814\ : InMux
    port map (
            O => \N__35743\,
            I => \N__35722\
        );

    \I__6813\ : Span4Mux_v
    port map (
            O => \N__35740\,
            I => \N__35719\
        );

    \I__6812\ : InMux
    port map (
            O => \N__35739\,
            I => \N__35716\
        );

    \I__6811\ : InMux
    port map (
            O => \N__35738\,
            I => \N__35713\
        );

    \I__6810\ : Span4Mux_v
    port map (
            O => \N__35735\,
            I => \N__35708\
        );

    \I__6809\ : Span4Mux_h
    port map (
            O => \N__35732\,
            I => \N__35708\
        );

    \I__6808\ : InMux
    port map (
            O => \N__35731\,
            I => \N__35705\
        );

    \I__6807\ : Span4Mux_h
    port map (
            O => \N__35728\,
            I => \N__35698\
        );

    \I__6806\ : Span4Mux_h
    port map (
            O => \N__35725\,
            I => \N__35698\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__35722\,
            I => \N__35698\
        );

    \I__6804\ : Span4Mux_h
    port map (
            O => \N__35719\,
            I => \N__35695\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__35716\,
            I => un7_spon_9
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__35713\,
            I => un7_spon_9
        );

    \I__6801\ : Odrv4
    port map (
            O => \N__35708\,
            I => un7_spon_9
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__35705\,
            I => un7_spon_9
        );

    \I__6799\ : Odrv4
    port map (
            O => \N__35698\,
            I => un7_spon_9
        );

    \I__6798\ : Odrv4
    port map (
            O => \N__35695\,
            I => un7_spon_9
        );

    \I__6797\ : InMux
    port map (
            O => \N__35682\,
            I => \N__35678\
        );

    \I__6796\ : InMux
    port map (
            O => \N__35681\,
            I => \N__35675\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__35678\,
            I => \N__35672\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__35675\,
            I => \N__35669\
        );

    \I__6793\ : Odrv4
    port map (
            O => \N__35672\,
            I => \sEEACQZ0Z_9\
        );

    \I__6792\ : Odrv4
    port map (
            O => \N__35669\,
            I => \sEEACQZ0Z_9\
        );

    \I__6791\ : CascadeMux
    port map (
            O => \N__35664\,
            I => \N__35661\
        );

    \I__6790\ : InMux
    port map (
            O => \N__35661\,
            I => \N__35658\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__35658\,
            I => \sEEACQ_i_9\
        );

    \I__6788\ : CascadeMux
    port map (
            O => \N__35655\,
            I => \N__35651\
        );

    \I__6787\ : CascadeMux
    port map (
            O => \N__35654\,
            I => \N__35648\
        );

    \I__6786\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35643\
        );

    \I__6785\ : InMux
    port map (
            O => \N__35648\,
            I => \N__35640\
        );

    \I__6784\ : InMux
    port map (
            O => \N__35647\,
            I => \N__35637\
        );

    \I__6783\ : InMux
    port map (
            O => \N__35646\,
            I => \N__35634\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__35643\,
            I => \N__35628\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__35640\,
            I => \N__35624\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__35637\,
            I => \N__35621\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__35634\,
            I => \N__35618\
        );

    \I__6778\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35614\
        );

    \I__6777\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35609\
        );

    \I__6776\ : InMux
    port map (
            O => \N__35631\,
            I => \N__35609\
        );

    \I__6775\ : Span4Mux_h
    port map (
            O => \N__35628\,
            I => \N__35606\
        );

    \I__6774\ : InMux
    port map (
            O => \N__35627\,
            I => \N__35603\
        );

    \I__6773\ : Span4Mux_h
    port map (
            O => \N__35624\,
            I => \N__35598\
        );

    \I__6772\ : Span4Mux_h
    port map (
            O => \N__35621\,
            I => \N__35598\
        );

    \I__6771\ : Span12Mux_s11_v
    port map (
            O => \N__35618\,
            I => \N__35595\
        );

    \I__6770\ : InMux
    port map (
            O => \N__35617\,
            I => \N__35592\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__35614\,
            I => \N__35589\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__35609\,
            I => \N__35586\
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__35606\,
            I => un7_spon_10
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__35603\,
            I => un7_spon_10
        );

    \I__6765\ : Odrv4
    port map (
            O => \N__35598\,
            I => un7_spon_10
        );

    \I__6764\ : Odrv12
    port map (
            O => \N__35595\,
            I => un7_spon_10
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__35592\,
            I => un7_spon_10
        );

    \I__6762\ : Odrv4
    port map (
            O => \N__35589\,
            I => un7_spon_10
        );

    \I__6761\ : Odrv4
    port map (
            O => \N__35586\,
            I => un7_spon_10
        );

    \I__6760\ : InMux
    port map (
            O => \N__35571\,
            I => \N__35568\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__35568\,
            I => \N__35564\
        );

    \I__6758\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35561\
        );

    \I__6757\ : Span4Mux_h
    port map (
            O => \N__35564\,
            I => \N__35558\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__35561\,
            I => \N__35555\
        );

    \I__6755\ : Odrv4
    port map (
            O => \N__35558\,
            I => \sEEACQZ0Z_10\
        );

    \I__6754\ : Odrv12
    port map (
            O => \N__35555\,
            I => \sEEACQZ0Z_10\
        );

    \I__6753\ : CascadeMux
    port map (
            O => \N__35550\,
            I => \N__35547\
        );

    \I__6752\ : InMux
    port map (
            O => \N__35547\,
            I => \N__35544\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__35544\,
            I => \sEEACQ_i_10\
        );

    \I__6750\ : InMux
    port map (
            O => \N__35541\,
            I => \N__35537\
        );

    \I__6749\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35533\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__35537\,
            I => \N__35529\
        );

    \I__6747\ : InMux
    port map (
            O => \N__35536\,
            I => \N__35526\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__35533\,
            I => \N__35523\
        );

    \I__6745\ : InMux
    port map (
            O => \N__35532\,
            I => \N__35517\
        );

    \I__6744\ : Span4Mux_h
    port map (
            O => \N__35529\,
            I => \N__35511\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__35526\,
            I => \N__35511\
        );

    \I__6742\ : Span4Mux_v
    port map (
            O => \N__35523\,
            I => \N__35508\
        );

    \I__6741\ : InMux
    port map (
            O => \N__35522\,
            I => \N__35503\
        );

    \I__6740\ : InMux
    port map (
            O => \N__35521\,
            I => \N__35503\
        );

    \I__6739\ : InMux
    port map (
            O => \N__35520\,
            I => \N__35500\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__35517\,
            I => \N__35497\
        );

    \I__6737\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35493\
        );

    \I__6736\ : Span4Mux_v
    port map (
            O => \N__35511\,
            I => \N__35488\
        );

    \I__6735\ : Span4Mux_h
    port map (
            O => \N__35508\,
            I => \N__35488\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__35503\,
            I => \N__35485\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__35500\,
            I => \N__35482\
        );

    \I__6732\ : Span4Mux_h
    port map (
            O => \N__35497\,
            I => \N__35479\
        );

    \I__6731\ : InMux
    port map (
            O => \N__35496\,
            I => \N__35476\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__35493\,
            I => un7_spon_11
        );

    \I__6729\ : Odrv4
    port map (
            O => \N__35488\,
            I => un7_spon_11
        );

    \I__6728\ : Odrv4
    port map (
            O => \N__35485\,
            I => un7_spon_11
        );

    \I__6727\ : Odrv4
    port map (
            O => \N__35482\,
            I => un7_spon_11
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__35479\,
            I => un7_spon_11
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__35476\,
            I => un7_spon_11
        );

    \I__6724\ : InMux
    port map (
            O => \N__35463\,
            I => \N__35459\
        );

    \I__6723\ : InMux
    port map (
            O => \N__35462\,
            I => \N__35456\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__35459\,
            I => \N__35453\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__35456\,
            I => \N__35450\
        );

    \I__6720\ : Odrv4
    port map (
            O => \N__35453\,
            I => \sEEACQZ0Z_11\
        );

    \I__6719\ : Odrv12
    port map (
            O => \N__35450\,
            I => \sEEACQZ0Z_11\
        );

    \I__6718\ : CascadeMux
    port map (
            O => \N__35445\,
            I => \N__35442\
        );

    \I__6717\ : InMux
    port map (
            O => \N__35442\,
            I => \N__35439\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__35439\,
            I => \sEEACQ_i_11\
        );

    \I__6715\ : InMux
    port map (
            O => \N__35436\,
            I => \N__35432\
        );

    \I__6714\ : InMux
    port map (
            O => \N__35435\,
            I => \N__35429\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__35432\,
            I => \N__35426\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__35429\,
            I => \N__35423\
        );

    \I__6711\ : Odrv4
    port map (
            O => \N__35426\,
            I => \sEEACQZ0Z_12\
        );

    \I__6710\ : Odrv12
    port map (
            O => \N__35423\,
            I => \sEEACQZ0Z_12\
        );

    \I__6709\ : CascadeMux
    port map (
            O => \N__35418\,
            I => \N__35415\
        );

    \I__6708\ : InMux
    port map (
            O => \N__35415\,
            I => \N__35411\
        );

    \I__6707\ : CascadeMux
    port map (
            O => \N__35414\,
            I => \N__35406\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__35411\,
            I => \N__35403\
        );

    \I__6705\ : InMux
    port map (
            O => \N__35410\,
            I => \N__35400\
        );

    \I__6704\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35397\
        );

    \I__6703\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35393\
        );

    \I__6702\ : Span4Mux_h
    port map (
            O => \N__35403\,
            I => \N__35388\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__35400\,
            I => \N__35388\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__35397\,
            I => \N__35385\
        );

    \I__6699\ : CascadeMux
    port map (
            O => \N__35396\,
            I => \N__35381\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__35393\,
            I => \N__35376\
        );

    \I__6697\ : Span4Mux_h
    port map (
            O => \N__35388\,
            I => \N__35373\
        );

    \I__6696\ : Span4Mux_h
    port map (
            O => \N__35385\,
            I => \N__35370\
        );

    \I__6695\ : InMux
    port map (
            O => \N__35384\,
            I => \N__35366\
        );

    \I__6694\ : InMux
    port map (
            O => \N__35381\,
            I => \N__35361\
        );

    \I__6693\ : InMux
    port map (
            O => \N__35380\,
            I => \N__35361\
        );

    \I__6692\ : InMux
    port map (
            O => \N__35379\,
            I => \N__35358\
        );

    \I__6691\ : Span4Mux_v
    port map (
            O => \N__35376\,
            I => \N__35353\
        );

    \I__6690\ : Span4Mux_v
    port map (
            O => \N__35373\,
            I => \N__35353\
        );

    \I__6689\ : Span4Mux_h
    port map (
            O => \N__35370\,
            I => \N__35350\
        );

    \I__6688\ : InMux
    port map (
            O => \N__35369\,
            I => \N__35347\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__35366\,
            I => \N__35344\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__35361\,
            I => \N__35341\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__35358\,
            I => un7_spon_12
        );

    \I__6684\ : Odrv4
    port map (
            O => \N__35353\,
            I => un7_spon_12
        );

    \I__6683\ : Odrv4
    port map (
            O => \N__35350\,
            I => un7_spon_12
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__35347\,
            I => un7_spon_12
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__35344\,
            I => un7_spon_12
        );

    \I__6680\ : Odrv4
    port map (
            O => \N__35341\,
            I => un7_spon_12
        );

    \I__6679\ : CascadeMux
    port map (
            O => \N__35328\,
            I => \N__35325\
        );

    \I__6678\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35322\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__35322\,
            I => \sEEACQ_i_12\
        );

    \I__6676\ : CascadeMux
    port map (
            O => \N__35319\,
            I => \N__35316\
        );

    \I__6675\ : InMux
    port map (
            O => \N__35316\,
            I => \N__35312\
        );

    \I__6674\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35307\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__35312\,
            I => \N__35303\
        );

    \I__6672\ : InMux
    port map (
            O => \N__35311\,
            I => \N__35299\
        );

    \I__6671\ : CascadeMux
    port map (
            O => \N__35310\,
            I => \N__35295\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__35307\,
            I => \N__35292\
        );

    \I__6669\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35288\
        );

    \I__6668\ : Span4Mux_h
    port map (
            O => \N__35303\,
            I => \N__35285\
        );

    \I__6667\ : InMux
    port map (
            O => \N__35302\,
            I => \N__35281\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__35299\,
            I => \N__35278\
        );

    \I__6665\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35273\
        );

    \I__6664\ : InMux
    port map (
            O => \N__35295\,
            I => \N__35273\
        );

    \I__6663\ : Span4Mux_v
    port map (
            O => \N__35292\,
            I => \N__35270\
        );

    \I__6662\ : InMux
    port map (
            O => \N__35291\,
            I => \N__35267\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__35288\,
            I => \N__35264\
        );

    \I__6660\ : Span4Mux_h
    port map (
            O => \N__35285\,
            I => \N__35261\
        );

    \I__6659\ : InMux
    port map (
            O => \N__35284\,
            I => \N__35258\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__35281\,
            I => \N__35255\
        );

    \I__6657\ : Span4Mux_h
    port map (
            O => \N__35278\,
            I => \N__35250\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__35273\,
            I => \N__35250\
        );

    \I__6655\ : Odrv4
    port map (
            O => \N__35270\,
            I => un7_spon_13
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__35267\,
            I => un7_spon_13
        );

    \I__6653\ : Odrv12
    port map (
            O => \N__35264\,
            I => un7_spon_13
        );

    \I__6652\ : Odrv4
    port map (
            O => \N__35261\,
            I => un7_spon_13
        );

    \I__6651\ : LocalMux
    port map (
            O => \N__35258\,
            I => un7_spon_13
        );

    \I__6650\ : Odrv4
    port map (
            O => \N__35255\,
            I => un7_spon_13
        );

    \I__6649\ : Odrv4
    port map (
            O => \N__35250\,
            I => un7_spon_13
        );

    \I__6648\ : InMux
    port map (
            O => \N__35235\,
            I => \N__35232\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__35232\,
            I => \N__35228\
        );

    \I__6646\ : InMux
    port map (
            O => \N__35231\,
            I => \N__35225\
        );

    \I__6645\ : Span4Mux_v
    port map (
            O => \N__35228\,
            I => \N__35222\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__35225\,
            I => \N__35219\
        );

    \I__6643\ : Odrv4
    port map (
            O => \N__35222\,
            I => \sEEACQZ0Z_13\
        );

    \I__6642\ : Odrv12
    port map (
            O => \N__35219\,
            I => \sEEACQZ0Z_13\
        );

    \I__6641\ : InMux
    port map (
            O => \N__35214\,
            I => \N__35211\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__35211\,
            I => \sEEACQ_i_13\
        );

    \I__6639\ : CascadeMux
    port map (
            O => \N__35208\,
            I => \N__35205\
        );

    \I__6638\ : InMux
    port map (
            O => \N__35205\,
            I => \N__35199\
        );

    \I__6637\ : CascadeMux
    port map (
            O => \N__35204\,
            I => \N__35196\
        );

    \I__6636\ : InMux
    port map (
            O => \N__35203\,
            I => \N__35192\
        );

    \I__6635\ : CascadeMux
    port map (
            O => \N__35202\,
            I => \N__35189\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__35199\,
            I => \N__35185\
        );

    \I__6633\ : InMux
    port map (
            O => \N__35196\,
            I => \N__35182\
        );

    \I__6632\ : InMux
    port map (
            O => \N__35195\,
            I => \N__35179\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__35192\,
            I => \N__35176\
        );

    \I__6630\ : InMux
    port map (
            O => \N__35189\,
            I => \N__35173\
        );

    \I__6629\ : InMux
    port map (
            O => \N__35188\,
            I => \N__35170\
        );

    \I__6628\ : Span4Mux_h
    port map (
            O => \N__35185\,
            I => \N__35165\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__35182\,
            I => \N__35165\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__35179\,
            I => \N__35160\
        );

    \I__6625\ : Span4Mux_h
    port map (
            O => \N__35176\,
            I => \N__35157\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__35173\,
            I => \N__35153\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__35170\,
            I => \N__35150\
        );

    \I__6622\ : Span4Mux_v
    port map (
            O => \N__35165\,
            I => \N__35147\
        );

    \I__6621\ : InMux
    port map (
            O => \N__35164\,
            I => \N__35144\
        );

    \I__6620\ : InMux
    port map (
            O => \N__35163\,
            I => \N__35141\
        );

    \I__6619\ : Span4Mux_v
    port map (
            O => \N__35160\,
            I => \N__35136\
        );

    \I__6618\ : Span4Mux_h
    port map (
            O => \N__35157\,
            I => \N__35136\
        );

    \I__6617\ : InMux
    port map (
            O => \N__35156\,
            I => \N__35133\
        );

    \I__6616\ : Span4Mux_v
    port map (
            O => \N__35153\,
            I => \N__35128\
        );

    \I__6615\ : Span4Mux_h
    port map (
            O => \N__35150\,
            I => \N__35128\
        );

    \I__6614\ : Odrv4
    port map (
            O => \N__35147\,
            I => un7_spon_14
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__35144\,
            I => un7_spon_14
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__35141\,
            I => un7_spon_14
        );

    \I__6611\ : Odrv4
    port map (
            O => \N__35136\,
            I => un7_spon_14
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__35133\,
            I => un7_spon_14
        );

    \I__6609\ : Odrv4
    port map (
            O => \N__35128\,
            I => un7_spon_14
        );

    \I__6608\ : InMux
    port map (
            O => \N__35115\,
            I => \N__35112\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__35112\,
            I => \N__35108\
        );

    \I__6606\ : InMux
    port map (
            O => \N__35111\,
            I => \N__35105\
        );

    \I__6605\ : Span4Mux_v
    port map (
            O => \N__35108\,
            I => \N__35100\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__35105\,
            I => \N__35100\
        );

    \I__6603\ : Odrv4
    port map (
            O => \N__35100\,
            I => \sEEACQZ0Z_14\
        );

    \I__6602\ : CascadeMux
    port map (
            O => \N__35097\,
            I => \N__35094\
        );

    \I__6601\ : InMux
    port map (
            O => \N__35094\,
            I => \N__35091\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__35091\,
            I => \sEEACQ_i_14\
        );

    \I__6599\ : InMux
    port map (
            O => \N__35088\,
            I => \N__35085\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__35085\,
            I => \sEEACQ_i_0\
        );

    \I__6597\ : InMux
    port map (
            O => \N__35082\,
            I => \N__35079\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__35079\,
            I => \N__35076\
        );

    \I__6595\ : Span4Mux_v
    port map (
            O => \N__35076\,
            I => \N__35072\
        );

    \I__6594\ : InMux
    port map (
            O => \N__35075\,
            I => \N__35069\
        );

    \I__6593\ : Odrv4
    port map (
            O => \N__35072\,
            I => \sEEACQZ0Z_1\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__35069\,
            I => \sEEACQZ0Z_1\
        );

    \I__6591\ : CascadeMux
    port map (
            O => \N__35064\,
            I => \N__35059\
        );

    \I__6590\ : CascadeMux
    port map (
            O => \N__35063\,
            I => \N__35055\
        );

    \I__6589\ : InMux
    port map (
            O => \N__35062\,
            I => \N__35052\
        );

    \I__6588\ : InMux
    port map (
            O => \N__35059\,
            I => \N__35047\
        );

    \I__6587\ : InMux
    port map (
            O => \N__35058\,
            I => \N__35044\
        );

    \I__6586\ : InMux
    port map (
            O => \N__35055\,
            I => \N__35041\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__35052\,
            I => \N__35038\
        );

    \I__6584\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35035\
        );

    \I__6583\ : InMux
    port map (
            O => \N__35050\,
            I => \N__35031\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__35047\,
            I => \N__35028\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__35044\,
            I => \N__35025\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__35041\,
            I => \N__35020\
        );

    \I__6579\ : Span4Mux_v
    port map (
            O => \N__35038\,
            I => \N__35017\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__35035\,
            I => \N__35014\
        );

    \I__6577\ : InMux
    port map (
            O => \N__35034\,
            I => \N__35011\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__35031\,
            I => \N__35008\
        );

    \I__6575\ : Span4Mux_h
    port map (
            O => \N__35028\,
            I => \N__35003\
        );

    \I__6574\ : Span4Mux_h
    port map (
            O => \N__35025\,
            I => \N__35003\
        );

    \I__6573\ : InMux
    port map (
            O => \N__35024\,
            I => \N__35000\
        );

    \I__6572\ : InMux
    port map (
            O => \N__35023\,
            I => \N__34997\
        );

    \I__6571\ : Span4Mux_v
    port map (
            O => \N__35020\,
            I => \N__34990\
        );

    \I__6570\ : Span4Mux_h
    port map (
            O => \N__35017\,
            I => \N__34990\
        );

    \I__6569\ : Span4Mux_v
    port map (
            O => \N__35014\,
            I => \N__34990\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__35011\,
            I => un7_spon_1
        );

    \I__6567\ : Odrv4
    port map (
            O => \N__35008\,
            I => un7_spon_1
        );

    \I__6566\ : Odrv4
    port map (
            O => \N__35003\,
            I => un7_spon_1
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__35000\,
            I => un7_spon_1
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__34997\,
            I => un7_spon_1
        );

    \I__6563\ : Odrv4
    port map (
            O => \N__34990\,
            I => un7_spon_1
        );

    \I__6562\ : CascadeMux
    port map (
            O => \N__34977\,
            I => \N__34974\
        );

    \I__6561\ : InMux
    port map (
            O => \N__34974\,
            I => \N__34971\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__34971\,
            I => \sEEACQ_i_1\
        );

    \I__6559\ : CascadeMux
    port map (
            O => \N__34968\,
            I => \N__34965\
        );

    \I__6558\ : InMux
    port map (
            O => \N__34965\,
            I => \N__34961\
        );

    \I__6557\ : CascadeMux
    port map (
            O => \N__34964\,
            I => \N__34958\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__34961\,
            I => \N__34953\
        );

    \I__6555\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34950\
        );

    \I__6554\ : InMux
    port map (
            O => \N__34957\,
            I => \N__34946\
        );

    \I__6553\ : InMux
    port map (
            O => \N__34956\,
            I => \N__34943\
        );

    \I__6552\ : Span4Mux_v
    port map (
            O => \N__34953\,
            I => \N__34936\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__34950\,
            I => \N__34936\
        );

    \I__6550\ : InMux
    port map (
            O => \N__34949\,
            I => \N__34933\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__34946\,
            I => \N__34930\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__34943\,
            I => \N__34926\
        );

    \I__6547\ : InMux
    port map (
            O => \N__34942\,
            I => \N__34922\
        );

    \I__6546\ : InMux
    port map (
            O => \N__34941\,
            I => \N__34919\
        );

    \I__6545\ : Span4Mux_h
    port map (
            O => \N__34936\,
            I => \N__34914\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__34933\,
            I => \N__34914\
        );

    \I__6543\ : Span4Mux_h
    port map (
            O => \N__34930\,
            I => \N__34911\
        );

    \I__6542\ : InMux
    port map (
            O => \N__34929\,
            I => \N__34908\
        );

    \I__6541\ : Span12Mux_v
    port map (
            O => \N__34926\,
            I => \N__34905\
        );

    \I__6540\ : InMux
    port map (
            O => \N__34925\,
            I => \N__34902\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__34922\,
            I => \N__34899\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__34919\,
            I => un7_spon_2
        );

    \I__6537\ : Odrv4
    port map (
            O => \N__34914\,
            I => un7_spon_2
        );

    \I__6536\ : Odrv4
    port map (
            O => \N__34911\,
            I => un7_spon_2
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__34908\,
            I => un7_spon_2
        );

    \I__6534\ : Odrv12
    port map (
            O => \N__34905\,
            I => un7_spon_2
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__34902\,
            I => un7_spon_2
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__34899\,
            I => un7_spon_2
        );

    \I__6531\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34881\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__34881\,
            I => \N__34878\
        );

    \I__6529\ : Span4Mux_h
    port map (
            O => \N__34878\,
            I => \N__34874\
        );

    \I__6528\ : InMux
    port map (
            O => \N__34877\,
            I => \N__34871\
        );

    \I__6527\ : Odrv4
    port map (
            O => \N__34874\,
            I => \sEEACQZ0Z_2\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__34871\,
            I => \sEEACQZ0Z_2\
        );

    \I__6525\ : CascadeMux
    port map (
            O => \N__34866\,
            I => \N__34863\
        );

    \I__6524\ : InMux
    port map (
            O => \N__34863\,
            I => \N__34860\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__34860\,
            I => \sEEACQ_i_2\
        );

    \I__6522\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34853\
        );

    \I__6521\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34848\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__34853\,
            I => \N__34845\
        );

    \I__6519\ : InMux
    port map (
            O => \N__34852\,
            I => \N__34842\
        );

    \I__6518\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34839\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__34848\,
            I => \N__34836\
        );

    \I__6516\ : Span4Mux_h
    port map (
            O => \N__34845\,
            I => \N__34828\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__34842\,
            I => \N__34828\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__34839\,
            I => \N__34824\
        );

    \I__6513\ : Span4Mux_v
    port map (
            O => \N__34836\,
            I => \N__34821\
        );

    \I__6512\ : InMux
    port map (
            O => \N__34835\,
            I => \N__34818\
        );

    \I__6511\ : InMux
    port map (
            O => \N__34834\,
            I => \N__34814\
        );

    \I__6510\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34811\
        );

    \I__6509\ : Span4Mux_h
    port map (
            O => \N__34828\,
            I => \N__34808\
        );

    \I__6508\ : InMux
    port map (
            O => \N__34827\,
            I => \N__34805\
        );

    \I__6507\ : Span4Mux_v
    port map (
            O => \N__34824\,
            I => \N__34800\
        );

    \I__6506\ : Span4Mux_h
    port map (
            O => \N__34821\,
            I => \N__34800\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__34818\,
            I => \N__34797\
        );

    \I__6504\ : InMux
    port map (
            O => \N__34817\,
            I => \N__34794\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__34814\,
            I => un7_spon_3
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__34811\,
            I => un7_spon_3
        );

    \I__6501\ : Odrv4
    port map (
            O => \N__34808\,
            I => un7_spon_3
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__34805\,
            I => un7_spon_3
        );

    \I__6499\ : Odrv4
    port map (
            O => \N__34800\,
            I => un7_spon_3
        );

    \I__6498\ : Odrv4
    port map (
            O => \N__34797\,
            I => un7_spon_3
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__34794\,
            I => un7_spon_3
        );

    \I__6496\ : InMux
    port map (
            O => \N__34779\,
            I => \N__34776\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__34776\,
            I => \N__34773\
        );

    \I__6494\ : Span4Mux_h
    port map (
            O => \N__34773\,
            I => \N__34769\
        );

    \I__6493\ : InMux
    port map (
            O => \N__34772\,
            I => \N__34766\
        );

    \I__6492\ : Odrv4
    port map (
            O => \N__34769\,
            I => \sEEACQZ0Z_3\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__34766\,
            I => \sEEACQZ0Z_3\
        );

    \I__6490\ : CascadeMux
    port map (
            O => \N__34761\,
            I => \N__34758\
        );

    \I__6489\ : InMux
    port map (
            O => \N__34758\,
            I => \N__34755\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__34755\,
            I => \sEEACQ_i_3\
        );

    \I__6487\ : InMux
    port map (
            O => \N__34752\,
            I => \N__34749\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__34749\,
            I => \N__34746\
        );

    \I__6485\ : Span4Mux_h
    port map (
            O => \N__34746\,
            I => \N__34742\
        );

    \I__6484\ : InMux
    port map (
            O => \N__34745\,
            I => \N__34739\
        );

    \I__6483\ : Odrv4
    port map (
            O => \N__34742\,
            I => \sEEACQZ0Z_4\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__34739\,
            I => \sEEACQZ0Z_4\
        );

    \I__6481\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34731\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__34731\,
            I => \sEEACQ_i_4\
        );

    \I__6479\ : InMux
    port map (
            O => \N__34728\,
            I => \N__34723\
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__34727\,
            I => \N__34720\
        );

    \I__6477\ : InMux
    port map (
            O => \N__34726\,
            I => \N__34717\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__34723\,
            I => \N__34714\
        );

    \I__6475\ : InMux
    port map (
            O => \N__34720\,
            I => \N__34711\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__34717\,
            I => \N__34707\
        );

    \I__6473\ : Span4Mux_h
    port map (
            O => \N__34714\,
            I => \N__34701\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__34711\,
            I => \N__34701\
        );

    \I__6471\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34696\
        );

    \I__6470\ : Span4Mux_h
    port map (
            O => \N__34707\,
            I => \N__34692\
        );

    \I__6469\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34688\
        );

    \I__6468\ : Span4Mux_v
    port map (
            O => \N__34701\,
            I => \N__34685\
        );

    \I__6467\ : InMux
    port map (
            O => \N__34700\,
            I => \N__34682\
        );

    \I__6466\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34679\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__34696\,
            I => \N__34676\
        );

    \I__6464\ : InMux
    port map (
            O => \N__34695\,
            I => \N__34673\
        );

    \I__6463\ : Span4Mux_h
    port map (
            O => \N__34692\,
            I => \N__34670\
        );

    \I__6462\ : InMux
    port map (
            O => \N__34691\,
            I => \N__34667\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__34688\,
            I => \N__34664\
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__34685\,
            I => un7_spon_5
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__34682\,
            I => un7_spon_5
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__34679\,
            I => un7_spon_5
        );

    \I__6457\ : Odrv12
    port map (
            O => \N__34676\,
            I => un7_spon_5
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__34673\,
            I => un7_spon_5
        );

    \I__6455\ : Odrv4
    port map (
            O => \N__34670\,
            I => un7_spon_5
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__34667\,
            I => un7_spon_5
        );

    \I__6453\ : Odrv4
    port map (
            O => \N__34664\,
            I => un7_spon_5
        );

    \I__6452\ : InMux
    port map (
            O => \N__34647\,
            I => \N__34644\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__34644\,
            I => \N__34641\
        );

    \I__6450\ : Span4Mux_v
    port map (
            O => \N__34641\,
            I => \N__34637\
        );

    \I__6449\ : InMux
    port map (
            O => \N__34640\,
            I => \N__34634\
        );

    \I__6448\ : Odrv4
    port map (
            O => \N__34637\,
            I => \sEEACQZ0Z_5\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__34634\,
            I => \sEEACQZ0Z_5\
        );

    \I__6446\ : CascadeMux
    port map (
            O => \N__34629\,
            I => \N__34626\
        );

    \I__6445\ : InMux
    port map (
            O => \N__34626\,
            I => \N__34623\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__34623\,
            I => \sEEACQ_i_5\
        );

    \I__6443\ : CascadeMux
    port map (
            O => \N__34620\,
            I => \N__34616\
        );

    \I__6442\ : CascadeMux
    port map (
            O => \N__34619\,
            I => \N__34613\
        );

    \I__6441\ : InMux
    port map (
            O => \N__34616\,
            I => \N__34609\
        );

    \I__6440\ : InMux
    port map (
            O => \N__34613\,
            I => \N__34606\
        );

    \I__6439\ : InMux
    port map (
            O => \N__34612\,
            I => \N__34602\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__34609\,
            I => \N__34598\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__34606\,
            I => \N__34595\
        );

    \I__6436\ : InMux
    port map (
            O => \N__34605\,
            I => \N__34591\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__34602\,
            I => \N__34588\
        );

    \I__6434\ : InMux
    port map (
            O => \N__34601\,
            I => \N__34585\
        );

    \I__6433\ : Span4Mux_v
    port map (
            O => \N__34598\,
            I => \N__34582\
        );

    \I__6432\ : Span4Mux_v
    port map (
            O => \N__34595\,
            I => \N__34579\
        );

    \I__6431\ : CascadeMux
    port map (
            O => \N__34594\,
            I => \N__34576\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__34591\,
            I => \N__34571\
        );

    \I__6429\ : Span4Mux_h
    port map (
            O => \N__34588\,
            I => \N__34568\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__34585\,
            I => \N__34564\
        );

    \I__6427\ : Span4Mux_v
    port map (
            O => \N__34582\,
            I => \N__34561\
        );

    \I__6426\ : Span4Mux_v
    port map (
            O => \N__34579\,
            I => \N__34558\
        );

    \I__6425\ : InMux
    port map (
            O => \N__34576\,
            I => \N__34555\
        );

    \I__6424\ : InMux
    port map (
            O => \N__34575\,
            I => \N__34552\
        );

    \I__6423\ : InMux
    port map (
            O => \N__34574\,
            I => \N__34549\
        );

    \I__6422\ : Span4Mux_v
    port map (
            O => \N__34571\,
            I => \N__34544\
        );

    \I__6421\ : Span4Mux_h
    port map (
            O => \N__34568\,
            I => \N__34544\
        );

    \I__6420\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34541\
        );

    \I__6419\ : Span4Mux_h
    port map (
            O => \N__34564\,
            I => \N__34538\
        );

    \I__6418\ : Odrv4
    port map (
            O => \N__34561\,
            I => un7_spon_6
        );

    \I__6417\ : Odrv4
    port map (
            O => \N__34558\,
            I => un7_spon_6
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__34555\,
            I => un7_spon_6
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__34552\,
            I => un7_spon_6
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__34549\,
            I => un7_spon_6
        );

    \I__6413\ : Odrv4
    port map (
            O => \N__34544\,
            I => un7_spon_6
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__34541\,
            I => un7_spon_6
        );

    \I__6411\ : Odrv4
    port map (
            O => \N__34538\,
            I => un7_spon_6
        );

    \I__6410\ : InMux
    port map (
            O => \N__34521\,
            I => \N__34518\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__34518\,
            I => \N__34515\
        );

    \I__6408\ : Span4Mux_v
    port map (
            O => \N__34515\,
            I => \N__34511\
        );

    \I__6407\ : InMux
    port map (
            O => \N__34514\,
            I => \N__34508\
        );

    \I__6406\ : Odrv4
    port map (
            O => \N__34511\,
            I => \sEEACQZ0Z_6\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__34508\,
            I => \sEEACQZ0Z_6\
        );

    \I__6404\ : CascadeMux
    port map (
            O => \N__34503\,
            I => \N__34500\
        );

    \I__6403\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34497\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__34497\,
            I => \sEEACQ_i_6\
        );

    \I__6401\ : CascadeMux
    port map (
            O => \N__34494\,
            I => \N__34490\
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__34493\,
            I => \N__34486\
        );

    \I__6399\ : InMux
    port map (
            O => \N__34490\,
            I => \N__34483\
        );

    \I__6398\ : CascadeMux
    port map (
            O => \N__34489\,
            I => \N__34480\
        );

    \I__6397\ : InMux
    port map (
            O => \N__34486\,
            I => \N__34476\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__34483\,
            I => \N__34472\
        );

    \I__6395\ : InMux
    port map (
            O => \N__34480\,
            I => \N__34469\
        );

    \I__6394\ : InMux
    port map (
            O => \N__34479\,
            I => \N__34466\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__34476\,
            I => \N__34463\
        );

    \I__6392\ : CascadeMux
    port map (
            O => \N__34475\,
            I => \N__34460\
        );

    \I__6391\ : Span4Mux_h
    port map (
            O => \N__34472\,
            I => \N__34455\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__34469\,
            I => \N__34455\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__34466\,
            I => \N__34449\
        );

    \I__6388\ : Span4Mux_h
    port map (
            O => \N__34463\,
            I => \N__34446\
        );

    \I__6387\ : InMux
    port map (
            O => \N__34460\,
            I => \N__34442\
        );

    \I__6386\ : Span4Mux_v
    port map (
            O => \N__34455\,
            I => \N__34439\
        );

    \I__6385\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34436\
        );

    \I__6384\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34433\
        );

    \I__6383\ : InMux
    port map (
            O => \N__34452\,
            I => \N__34430\
        );

    \I__6382\ : Span4Mux_v
    port map (
            O => \N__34449\,
            I => \N__34425\
        );

    \I__6381\ : Span4Mux_h
    port map (
            O => \N__34446\,
            I => \N__34425\
        );

    \I__6380\ : InMux
    port map (
            O => \N__34445\,
            I => \N__34422\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__34442\,
            I => \N__34419\
        );

    \I__6378\ : Odrv4
    port map (
            O => \N__34439\,
            I => un7_spon_7
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__34436\,
            I => un7_spon_7
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__34433\,
            I => un7_spon_7
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__34430\,
            I => un7_spon_7
        );

    \I__6374\ : Odrv4
    port map (
            O => \N__34425\,
            I => un7_spon_7
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__34422\,
            I => un7_spon_7
        );

    \I__6372\ : Odrv4
    port map (
            O => \N__34419\,
            I => un7_spon_7
        );

    \I__6371\ : InMux
    port map (
            O => \N__34404\,
            I => \N__34401\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__34401\,
            I => \N__34398\
        );

    \I__6369\ : Span4Mux_h
    port map (
            O => \N__34398\,
            I => \N__34394\
        );

    \I__6368\ : InMux
    port map (
            O => \N__34397\,
            I => \N__34391\
        );

    \I__6367\ : Odrv4
    port map (
            O => \N__34394\,
            I => \sEEACQZ0Z_7\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__34391\,
            I => \sEEACQZ0Z_7\
        );

    \I__6365\ : InMux
    port map (
            O => \N__34386\,
            I => \N__34383\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__34383\,
            I => \sEEACQ_i_7\
        );

    \I__6363\ : CEMux
    port map (
            O => \N__34380\,
            I => \N__34377\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__34377\,
            I => \N__34374\
        );

    \I__6361\ : Span4Mux_h
    port map (
            O => \N__34374\,
            I => \N__34371\
        );

    \I__6360\ : Span4Mux_h
    port map (
            O => \N__34371\,
            I => \N__34368\
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__34368\,
            I => \sDAC_mem_31_1_sqmuxa\
        );

    \I__6358\ : InMux
    port map (
            O => \N__34365\,
            I => \N__34361\
        );

    \I__6357\ : InMux
    port map (
            O => \N__34364\,
            I => \N__34358\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__34361\,
            I => \N__34355\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__34358\,
            I => \sCounterADCZ0Z_3\
        );

    \I__6354\ : Odrv4
    port map (
            O => \N__34355\,
            I => \sCounterADCZ0Z_3\
        );

    \I__6353\ : InMux
    port map (
            O => \N__34350\,
            I => \N__34346\
        );

    \I__6352\ : InMux
    port map (
            O => \N__34349\,
            I => \N__34343\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__34346\,
            I => \N__34338\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__34343\,
            I => \N__34338\
        );

    \I__6349\ : Odrv4
    port map (
            O => \N__34338\,
            I => \sCounterADCZ0Z_2\
        );

    \I__6348\ : InMux
    port map (
            O => \N__34335\,
            I => \N__34332\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__34332\,
            I => \sEEADC_freqZ0Z_2\
        );

    \I__6346\ : CascadeMux
    port map (
            O => \N__34329\,
            I => \N__34326\
        );

    \I__6345\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34323\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__34323\,
            I => \sEEADC_freqZ0Z_3\
        );

    \I__6343\ : InMux
    port map (
            O => \N__34320\,
            I => \N__34316\
        );

    \I__6342\ : InMux
    port map (
            O => \N__34319\,
            I => \N__34313\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__34316\,
            I => \N__34308\
        );

    \I__6340\ : LocalMux
    port map (
            O => \N__34313\,
            I => \N__34308\
        );

    \I__6339\ : Odrv12
    port map (
            O => \N__34308\,
            I => \sCounterADCZ0Z_5\
        );

    \I__6338\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34301\
        );

    \I__6337\ : InMux
    port map (
            O => \N__34304\,
            I => \N__34298\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__34301\,
            I => \N__34295\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__34298\,
            I => \sCounterADCZ0Z_4\
        );

    \I__6334\ : Odrv4
    port map (
            O => \N__34295\,
            I => \sCounterADCZ0Z_4\
        );

    \I__6333\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34287\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__34287\,
            I => \sEEADC_freqZ0Z_4\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__34284\,
            I => \N__34281\
        );

    \I__6330\ : InMux
    port map (
            O => \N__34281\,
            I => \N__34278\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__34278\,
            I => \sEEADC_freqZ0Z_5\
        );

    \I__6328\ : InMux
    port map (
            O => \N__34275\,
            I => \N__34271\
        );

    \I__6327\ : InMux
    port map (
            O => \N__34274\,
            I => \N__34268\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__34271\,
            I => \N__34265\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__34268\,
            I => \sCounterADCZ0Z_6\
        );

    \I__6324\ : Odrv4
    port map (
            O => \N__34265\,
            I => \sCounterADCZ0Z_6\
        );

    \I__6323\ : InMux
    port map (
            O => \N__34260\,
            I => \N__34256\
        );

    \I__6322\ : InMux
    port map (
            O => \N__34259\,
            I => \N__34253\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__34256\,
            I => \N__34250\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__34253\,
            I => \sCounterADCZ0Z_7\
        );

    \I__6319\ : Odrv12
    port map (
            O => \N__34250\,
            I => \sCounterADCZ0Z_7\
        );

    \I__6318\ : CascadeMux
    port map (
            O => \N__34245\,
            I => \N__34240\
        );

    \I__6317\ : CascadeMux
    port map (
            O => \N__34244\,
            I => \N__34237\
        );

    \I__6316\ : CascadeMux
    port map (
            O => \N__34243\,
            I => \N__34234\
        );

    \I__6315\ : InMux
    port map (
            O => \N__34240\,
            I => \N__34231\
        );

    \I__6314\ : InMux
    port map (
            O => \N__34237\,
            I => \N__34227\
        );

    \I__6313\ : InMux
    port map (
            O => \N__34234\,
            I => \N__34223\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__34231\,
            I => \N__34220\
        );

    \I__6311\ : InMux
    port map (
            O => \N__34230\,
            I => \N__34217\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__34227\,
            I => \N__34214\
        );

    \I__6309\ : InMux
    port map (
            O => \N__34226\,
            I => \N__34211\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__34223\,
            I => \N__34208\
        );

    \I__6307\ : Span4Mux_h
    port map (
            O => \N__34220\,
            I => \N__34202\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__34217\,
            I => \N__34202\
        );

    \I__6305\ : Span4Mux_h
    port map (
            O => \N__34214\,
            I => \N__34197\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__34211\,
            I => \N__34194\
        );

    \I__6303\ : Span4Mux_v
    port map (
            O => \N__34208\,
            I => \N__34191\
        );

    \I__6302\ : InMux
    port map (
            O => \N__34207\,
            I => \N__34188\
        );

    \I__6301\ : Span4Mux_h
    port map (
            O => \N__34202\,
            I => \N__34185\
        );

    \I__6300\ : InMux
    port map (
            O => \N__34201\,
            I => \N__34182\
        );

    \I__6299\ : InMux
    port map (
            O => \N__34200\,
            I => \N__34179\
        );

    \I__6298\ : Span4Mux_h
    port map (
            O => \N__34197\,
            I => \N__34174\
        );

    \I__6297\ : Span4Mux_v
    port map (
            O => \N__34194\,
            I => \N__34174\
        );

    \I__6296\ : Odrv4
    port map (
            O => \N__34191\,
            I => un7_spon_0
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__34188\,
            I => un7_spon_0
        );

    \I__6294\ : Odrv4
    port map (
            O => \N__34185\,
            I => un7_spon_0
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__34182\,
            I => un7_spon_0
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__34179\,
            I => un7_spon_0
        );

    \I__6291\ : Odrv4
    port map (
            O => \N__34174\,
            I => un7_spon_0
        );

    \I__6290\ : InMux
    port map (
            O => \N__34161\,
            I => \N__34158\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__34158\,
            I => \N__34155\
        );

    \I__6288\ : Span4Mux_v
    port map (
            O => \N__34155\,
            I => \N__34151\
        );

    \I__6287\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34148\
        );

    \I__6286\ : Odrv4
    port map (
            O => \N__34151\,
            I => \sEEACQZ0Z_0\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__34148\,
            I => \sEEACQZ0Z_0\
        );

    \I__6284\ : InMux
    port map (
            O => \N__34143\,
            I => \N__34140\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__34140\,
            I => \sDAC_data_RNO_19Z0Z_6\
        );

    \I__6282\ : InMux
    port map (
            O => \N__34137\,
            I => \N__34134\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__34134\,
            I => \sDAC_mem_12Z0Z_2\
        );

    \I__6280\ : InMux
    port map (
            O => \N__34131\,
            I => \N__34128\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__34128\,
            I => \sDAC_mem_12Z0Z_3\
        );

    \I__6278\ : CascadeMux
    port map (
            O => \N__34125\,
            I => \N__34122\
        );

    \I__6277\ : InMux
    port map (
            O => \N__34122\,
            I => \N__34119\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__34119\,
            I => \sDAC_mem_19Z0Z_1\
        );

    \I__6275\ : InMux
    port map (
            O => \N__34116\,
            I => \N__34113\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__34113\,
            I => \sDAC_mem_18Z0Z_1\
        );

    \I__6273\ : InMux
    port map (
            O => \N__34110\,
            I => \N__34107\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__34107\,
            I => \sDAC_mem_19Z0Z_2\
        );

    \I__6271\ : InMux
    port map (
            O => \N__34104\,
            I => \N__34101\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__34101\,
            I => \N__34098\
        );

    \I__6269\ : Odrv12
    port map (
            O => \N__34098\,
            I => \sDAC_data_RNO_30Z0Z_5\
        );

    \I__6268\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34092\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__34092\,
            I => \sDAC_mem_18Z0Z_2\
        );

    \I__6266\ : CEMux
    port map (
            O => \N__34089\,
            I => \N__34085\
        );

    \I__6265\ : CEMux
    port map (
            O => \N__34088\,
            I => \N__34082\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__34085\,
            I => \N__34079\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__34082\,
            I => \sDAC_mem_18_1_sqmuxa\
        );

    \I__6262\ : Odrv12
    port map (
            O => \N__34079\,
            I => \sDAC_mem_18_1_sqmuxa\
        );

    \I__6261\ : CascadeMux
    port map (
            O => \N__34074\,
            I => \sDAC_data_RNO_18Z0Z_5_cascade_\
        );

    \I__6260\ : InMux
    port map (
            O => \N__34071\,
            I => \N__34068\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__34068\,
            I => \sDAC_data_RNO_19Z0Z_5\
        );

    \I__6258\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34062\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__34062\,
            I => \N__34059\
        );

    \I__6256\ : Span4Mux_v
    port map (
            O => \N__34059\,
            I => \N__34056\
        );

    \I__6255\ : Odrv4
    port map (
            O => \N__34056\,
            I => \sDAC_data_2_24_ns_1_5\
        );

    \I__6254\ : CascadeMux
    port map (
            O => \N__34053\,
            I => \sDAC_data_RNO_18Z0Z_6_cascade_\
        );

    \I__6253\ : CascadeMux
    port map (
            O => \N__34050\,
            I => \op_le_op_le_un15_sdacdynlt4_cascade_\
        );

    \I__6252\ : InMux
    port map (
            O => \N__34047\,
            I => \N__34044\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__34044\,
            I => \N__34041\
        );

    \I__6250\ : Odrv12
    port map (
            O => \N__34041\,
            I => un17_sdacdyn_0
        );

    \I__6249\ : InMux
    port map (
            O => \N__34038\,
            I => \N__34035\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__34035\,
            I => \sDAC_mem_10Z0Z_7\
        );

    \I__6247\ : InMux
    port map (
            O => \N__34032\,
            I => \N__34029\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__34029\,
            I => \sDAC_mem_19Z0Z_7\
        );

    \I__6245\ : InMux
    port map (
            O => \N__34026\,
            I => \N__34023\
        );

    \I__6244\ : LocalMux
    port map (
            O => \N__34023\,
            I => \sDAC_mem_18Z0Z_7\
        );

    \I__6243\ : InMux
    port map (
            O => \N__34020\,
            I => \N__34017\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__34017\,
            I => \sDAC_mem_19Z0Z_0\
        );

    \I__6241\ : InMux
    port map (
            O => \N__34014\,
            I => \N__34011\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__34011\,
            I => \sDAC_mem_18Z0Z_0\
        );

    \I__6239\ : CascadeMux
    port map (
            O => \N__34008\,
            I => \N__34005\
        );

    \I__6238\ : InMux
    port map (
            O => \N__34005\,
            I => \N__34002\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__34002\,
            I => \N__33999\
        );

    \I__6236\ : Span4Mux_v
    port map (
            O => \N__33999\,
            I => \N__33996\
        );

    \I__6235\ : Odrv4
    port map (
            O => \N__33996\,
            I => \sDAC_mem_2Z0Z_6\
        );

    \I__6234\ : CascadeMux
    port map (
            O => \N__33993\,
            I => \sDAC_data_2_6_bm_1_9_cascade_\
        );

    \I__6233\ : InMux
    port map (
            O => \N__33990\,
            I => \N__33987\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__33987\,
            I => \sDAC_mem_3Z0Z_6\
        );

    \I__6231\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33981\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__33981\,
            I => \N__33978\
        );

    \I__6229\ : Span4Mux_h
    port map (
            O => \N__33978\,
            I => \N__33975\
        );

    \I__6228\ : Odrv4
    port map (
            O => \N__33975\,
            I => \sDAC_mem_33Z0Z_1\
        );

    \I__6227\ : CascadeMux
    port map (
            O => \N__33972\,
            I => \sDAC_data_RNO_26Z0Z_4_cascade_\
        );

    \I__6226\ : CascadeMux
    port map (
            O => \N__33969\,
            I => \N__33965\
        );

    \I__6225\ : CascadeMux
    port map (
            O => \N__33968\,
            I => \N__33962\
        );

    \I__6224\ : InMux
    port map (
            O => \N__33965\,
            I => \N__33957\
        );

    \I__6223\ : InMux
    port map (
            O => \N__33962\,
            I => \N__33957\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__33957\,
            I => \N__33954\
        );

    \I__6221\ : Span4Mux_v
    port map (
            O => \N__33954\,
            I => \N__33951\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__33951\,
            I => \sDAC_mem_1Z0Z_1\
        );

    \I__6219\ : InMux
    port map (
            O => \N__33948\,
            I => \N__33942\
        );

    \I__6218\ : InMux
    port map (
            O => \N__33947\,
            I => \N__33942\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__33942\,
            I => \sDAC_mem_32Z0Z_1\
        );

    \I__6216\ : InMux
    port map (
            O => \N__33939\,
            I => \N__33936\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__33936\,
            I => \sDAC_data_RNO_27Z0Z_4\
        );

    \I__6214\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33930\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__33930\,
            I => \N__33927\
        );

    \I__6212\ : Span4Mux_v
    port map (
            O => \N__33927\,
            I => \N__33924\
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__33924\,
            I => \sDAC_mem_33Z0Z_2\
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__33921\,
            I => \sDAC_data_RNO_26Z0Z_5_cascade_\
        );

    \I__6209\ : CascadeMux
    port map (
            O => \N__33918\,
            I => \N__33915\
        );

    \I__6208\ : InMux
    port map (
            O => \N__33915\,
            I => \N__33912\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__33912\,
            I => \N__33909\
        );

    \I__6206\ : Odrv12
    port map (
            O => \N__33909\,
            I => \sDAC_data_RNO_14Z0Z_5\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__33906\,
            I => \N__33903\
        );

    \I__6204\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33899\
        );

    \I__6203\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33896\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__33899\,
            I => \sDAC_mem_32Z0Z_2\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__33896\,
            I => \sDAC_mem_32Z0Z_2\
        );

    \I__6200\ : InMux
    port map (
            O => \N__33891\,
            I => \N__33887\
        );

    \I__6199\ : InMux
    port map (
            O => \N__33890\,
            I => \N__33884\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__33887\,
            I => \N__33879\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__33884\,
            I => \N__33879\
        );

    \I__6196\ : Span4Mux_v
    port map (
            O => \N__33879\,
            I => \N__33876\
        );

    \I__6195\ : Odrv4
    port map (
            O => \N__33876\,
            I => \sDAC_mem_1Z0Z_2\
        );

    \I__6194\ : InMux
    port map (
            O => \N__33873\,
            I => \N__33870\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__33870\,
            I => \N__33867\
        );

    \I__6192\ : Odrv4
    port map (
            O => \N__33867\,
            I => \sDAC_data_RNO_27Z0Z_5\
        );

    \I__6191\ : InMux
    port map (
            O => \N__33864\,
            I => \N__33861\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__33861\,
            I => \N__33858\
        );

    \I__6189\ : Span4Mux_v
    port map (
            O => \N__33858\,
            I => \N__33855\
        );

    \I__6188\ : Odrv4
    port map (
            O => \N__33855\,
            I => \sDAC_mem_33Z0Z_5\
        );

    \I__6187\ : CascadeMux
    port map (
            O => \N__33852\,
            I => \sDAC_data_RNO_27Z0Z_8_cascade_\
        );

    \I__6186\ : InMux
    port map (
            O => \N__33849\,
            I => \N__33843\
        );

    \I__6185\ : InMux
    port map (
            O => \N__33848\,
            I => \N__33843\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__33843\,
            I => \sDAC_mem_32Z0Z_5\
        );

    \I__6183\ : InMux
    port map (
            O => \N__33840\,
            I => \N__33837\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__33837\,
            I => \sDAC_data_RNO_26Z0Z_8\
        );

    \I__6181\ : CascadeMux
    port map (
            O => \N__33834\,
            I => \N__33830\
        );

    \I__6180\ : CascadeMux
    port map (
            O => \N__33833\,
            I => \N__33827\
        );

    \I__6179\ : InMux
    port map (
            O => \N__33830\,
            I => \N__33822\
        );

    \I__6178\ : InMux
    port map (
            O => \N__33827\,
            I => \N__33822\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__33822\,
            I => \sDAC_mem_1Z0Z_5\
        );

    \I__6176\ : InMux
    port map (
            O => \N__33819\,
            I => \N__33816\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__33816\,
            I => \N__33813\
        );

    \I__6174\ : Span4Mux_h
    port map (
            O => \N__33813\,
            I => \N__33810\
        );

    \I__6173\ : Odrv4
    port map (
            O => \N__33810\,
            I => \sDAC_mem_33Z0Z_6\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__33807\,
            I => \sDAC_data_RNO_26Z0Z_9_cascade_\
        );

    \I__6171\ : CascadeMux
    port map (
            O => \N__33804\,
            I => \N__33800\
        );

    \I__6170\ : CascadeMux
    port map (
            O => \N__33803\,
            I => \N__33797\
        );

    \I__6169\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33792\
        );

    \I__6168\ : InMux
    port map (
            O => \N__33797\,
            I => \N__33792\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__33792\,
            I => \N__33789\
        );

    \I__6166\ : Odrv4
    port map (
            O => \N__33789\,
            I => \sDAC_mem_32Z0Z_6\
        );

    \I__6165\ : InMux
    port map (
            O => \N__33786\,
            I => \N__33783\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__33783\,
            I => \sDAC_data_RNO_27Z0Z_9\
        );

    \I__6163\ : InMux
    port map (
            O => \N__33780\,
            I => \N__33774\
        );

    \I__6162\ : InMux
    port map (
            O => \N__33779\,
            I => \N__33774\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__33774\,
            I => \sDAC_mem_1Z0Z_6\
        );

    \I__6160\ : CascadeMux
    port map (
            O => \N__33771\,
            I => \sDAC_data_2_5_cascade_\
        );

    \I__6159\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33765\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__33765\,
            I => \N__33762\
        );

    \I__6157\ : Span4Mux_v
    port map (
            O => \N__33762\,
            I => \N__33759\
        );

    \I__6156\ : Odrv4
    port map (
            O => \N__33759\,
            I => \sDAC_dataZ0Z_5\
        );

    \I__6155\ : InMux
    port map (
            O => \N__33756\,
            I => \N__33753\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__33753\,
            I => \N__33750\
        );

    \I__6153\ : Odrv4
    port map (
            O => \N__33750\,
            I => \sDAC_mem_2Z0Z_2\
        );

    \I__6152\ : CascadeMux
    port map (
            O => \N__33747\,
            I => \sDAC_data_2_6_bm_1_5_cascade_\
        );

    \I__6151\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33741\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__33741\,
            I => \sDAC_mem_3Z0Z_2\
        );

    \I__6149\ : InMux
    port map (
            O => \N__33738\,
            I => \N__33735\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__33735\,
            I => \sDAC_data_RNO_15Z0Z_5\
        );

    \I__6147\ : CascadeMux
    port map (
            O => \N__33732\,
            I => \sDAC_data_2_20_am_1_7_cascade_\
        );

    \I__6146\ : CascadeMux
    port map (
            O => \N__33729\,
            I => \sDAC_data_RNO_17Z0Z_7_cascade_\
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__33726\,
            I => \sDAC_data_RNO_8Z0Z_7_cascade_\
        );

    \I__6144\ : InMux
    port map (
            O => \N__33723\,
            I => \N__33720\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__33720\,
            I => \sDAC_data_RNO_7Z0Z_7\
        );

    \I__6142\ : CascadeMux
    port map (
            O => \N__33717\,
            I => \sDAC_data_2_20_am_1_5_cascade_\
        );

    \I__6141\ : CascadeMux
    port map (
            O => \N__33714\,
            I => \sDAC_data_RNO_7Z0Z_5_cascade_\
        );

    \I__6140\ : InMux
    port map (
            O => \N__33711\,
            I => \N__33708\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__33708\,
            I => \sDAC_data_RNO_8Z0Z_5\
        );

    \I__6138\ : InMux
    port map (
            O => \N__33705\,
            I => \N__33702\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__33702\,
            I => \N__33699\
        );

    \I__6136\ : Odrv4
    port map (
            O => \N__33699\,
            I => \sDAC_data_RNO_21Z0Z_5\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__33696\,
            I => \sDAC_data_RNO_10Z0Z_5_cascade_\
        );

    \I__6134\ : InMux
    port map (
            O => \N__33693\,
            I => \N__33690\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__33690\,
            I => \sDAC_data_2_32_ns_1_5\
        );

    \I__6132\ : InMux
    port map (
            O => \N__33687\,
            I => \N__33684\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__33684\,
            I => \N__33681\
        );

    \I__6130\ : Odrv4
    port map (
            O => \N__33681\,
            I => \sDAC_data_RNO_5Z0Z_5\
        );

    \I__6129\ : CascadeMux
    port map (
            O => \N__33678\,
            I => \sDAC_data_2_14_ns_1_5_cascade_\
        );

    \I__6128\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33672\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__33672\,
            I => \N__33669\
        );

    \I__6126\ : Odrv4
    port map (
            O => \N__33669\,
            I => \sDAC_data_RNO_4Z0Z_5\
        );

    \I__6125\ : InMux
    port map (
            O => \N__33666\,
            I => \N__33663\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__33663\,
            I => \sDAC_data_RNO_2Z0Z_5\
        );

    \I__6123\ : CascadeMux
    port map (
            O => \N__33660\,
            I => \sDAC_data_RNO_1Z0Z_5_cascade_\
        );

    \I__6122\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33654\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__33654\,
            I => \sDAC_data_2_41_ns_1_5\
        );

    \I__6120\ : CascadeMux
    port map (
            O => \N__33651\,
            I => \sDAC_data_2_13_am_1_6_cascade_\
        );

    \I__6119\ : InMux
    port map (
            O => \N__33648\,
            I => \N__33645\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__33645\,
            I => \sDAC_mem_4Z0Z_3\
        );

    \I__6117\ : InMux
    port map (
            O => \N__33642\,
            I => \N__33639\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__33639\,
            I => \N__33636\
        );

    \I__6115\ : Span4Mux_v
    port map (
            O => \N__33636\,
            I => \N__33633\
        );

    \I__6114\ : Odrv4
    port map (
            O => \N__33633\,
            I => \sDAC_mem_4Z0Z_4\
        );

    \I__6113\ : CascadeMux
    port map (
            O => \N__33630\,
            I => \sDAC_data_2_13_am_1_7_cascade_\
        );

    \I__6112\ : CascadeMux
    port map (
            O => \N__33627\,
            I => \N__33624\
        );

    \I__6111\ : InMux
    port map (
            O => \N__33624\,
            I => \N__33621\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__33621\,
            I => \sDAC_mem_2Z0Z_0\
        );

    \I__6109\ : CascadeMux
    port map (
            O => \N__33618\,
            I => \sDAC_data_2_6_bm_1_3_cascade_\
        );

    \I__6108\ : InMux
    port map (
            O => \N__33615\,
            I => \N__33612\
        );

    \I__6107\ : LocalMux
    port map (
            O => \N__33612\,
            I => \sDAC_mem_3Z0Z_0\
        );

    \I__6106\ : CascadeMux
    port map (
            O => \N__33609\,
            I => \sDAC_data_RNO_17Z0Z_5_cascade_\
        );

    \I__6105\ : InMux
    port map (
            O => \N__33606\,
            I => \N__33603\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__33603\,
            I => \sDAC_mem_6Z0Z_0\
        );

    \I__6103\ : InMux
    port map (
            O => \N__33600\,
            I => \N__33597\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__33597\,
            I => \sDAC_mem_38Z0Z_1\
        );

    \I__6101\ : CascadeMux
    port map (
            O => \N__33594\,
            I => \sDAC_data_2_13_bm_1_4_cascade_\
        );

    \I__6100\ : InMux
    port map (
            O => \N__33591\,
            I => \N__33588\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__33588\,
            I => \sDAC_mem_6Z0Z_1\
        );

    \I__6098\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33582\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__33582\,
            I => \sDAC_mem_6Z0Z_2\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__33579\,
            I => \sDAC_data_2_13_bm_1_5_cascade_\
        );

    \I__6095\ : CascadeMux
    port map (
            O => \N__33576\,
            I => \sDAC_data_2_13_am_1_5_cascade_\
        );

    \I__6094\ : InMux
    port map (
            O => \N__33573\,
            I => \N__33570\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__33570\,
            I => \sDAC_mem_4Z0Z_2\
        );

    \I__6092\ : InMux
    port map (
            O => \N__33567\,
            I => \N__33532\
        );

    \I__6091\ : InMux
    port map (
            O => \N__33566\,
            I => \N__33532\
        );

    \I__6090\ : InMux
    port map (
            O => \N__33565\,
            I => \N__33532\
        );

    \I__6089\ : InMux
    port map (
            O => \N__33564\,
            I => \N__33532\
        );

    \I__6088\ : InMux
    port map (
            O => \N__33563\,
            I => \N__33523\
        );

    \I__6087\ : InMux
    port map (
            O => \N__33562\,
            I => \N__33523\
        );

    \I__6086\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33523\
        );

    \I__6085\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33523\
        );

    \I__6084\ : InMux
    port map (
            O => \N__33559\,
            I => \N__33514\
        );

    \I__6083\ : InMux
    port map (
            O => \N__33558\,
            I => \N__33514\
        );

    \I__6082\ : InMux
    port map (
            O => \N__33557\,
            I => \N__33514\
        );

    \I__6081\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33514\
        );

    \I__6080\ : InMux
    port map (
            O => \N__33555\,
            I => \N__33505\
        );

    \I__6079\ : InMux
    port map (
            O => \N__33554\,
            I => \N__33505\
        );

    \I__6078\ : InMux
    port map (
            O => \N__33553\,
            I => \N__33505\
        );

    \I__6077\ : InMux
    port map (
            O => \N__33552\,
            I => \N__33505\
        );

    \I__6076\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33494\
        );

    \I__6075\ : InMux
    port map (
            O => \N__33550\,
            I => \N__33494\
        );

    \I__6074\ : InMux
    port map (
            O => \N__33549\,
            I => \N__33494\
        );

    \I__6073\ : InMux
    port map (
            O => \N__33548\,
            I => \N__33494\
        );

    \I__6072\ : InMux
    port map (
            O => \N__33547\,
            I => \N__33485\
        );

    \I__6071\ : InMux
    port map (
            O => \N__33546\,
            I => \N__33485\
        );

    \I__6070\ : InMux
    port map (
            O => \N__33545\,
            I => \N__33485\
        );

    \I__6069\ : InMux
    port map (
            O => \N__33544\,
            I => \N__33485\
        );

    \I__6068\ : InMux
    port map (
            O => \N__33543\,
            I => \N__33479\
        );

    \I__6067\ : InMux
    port map (
            O => \N__33542\,
            I => \N__33479\
        );

    \I__6066\ : InMux
    port map (
            O => \N__33541\,
            I => \N__33476\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__33532\,
            I => \N__33470\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__33523\,
            I => \N__33470\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__33514\,
            I => \N__33465\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__33505\,
            I => \N__33465\
        );

    \I__6061\ : InMux
    port map (
            O => \N__33504\,
            I => \N__33460\
        );

    \I__6060\ : InMux
    port map (
            O => \N__33503\,
            I => \N__33460\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__33494\,
            I => \N__33453\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__33485\,
            I => \N__33450\
        );

    \I__6057\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33447\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__33479\,
            I => \N__33438\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__33476\,
            I => \N__33438\
        );

    \I__6054\ : InMux
    port map (
            O => \N__33475\,
            I => \N__33435\
        );

    \I__6053\ : Span4Mux_h
    port map (
            O => \N__33470\,
            I => \N__33431\
        );

    \I__6052\ : Span4Mux_h
    port map (
            O => \N__33465\,
            I => \N__33428\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__33460\,
            I => \N__33425\
        );

    \I__6050\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33416\
        );

    \I__6049\ : InMux
    port map (
            O => \N__33458\,
            I => \N__33416\
        );

    \I__6048\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33416\
        );

    \I__6047\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33416\
        );

    \I__6046\ : Span4Mux_v
    port map (
            O => \N__33453\,
            I => \N__33409\
        );

    \I__6045\ : Span4Mux_v
    port map (
            O => \N__33450\,
            I => \N__33409\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__33447\,
            I => \N__33409\
        );

    \I__6043\ : InMux
    port map (
            O => \N__33446\,
            I => \N__33400\
        );

    \I__6042\ : InMux
    port map (
            O => \N__33445\,
            I => \N__33400\
        );

    \I__6041\ : InMux
    port map (
            O => \N__33444\,
            I => \N__33400\
        );

    \I__6040\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33400\
        );

    \I__6039\ : Span4Mux_h
    port map (
            O => \N__33438\,
            I => \N__33395\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__33435\,
            I => \N__33395\
        );

    \I__6037\ : InMux
    port map (
            O => \N__33434\,
            I => \N__33392\
        );

    \I__6036\ : Span4Mux_v
    port map (
            O => \N__33431\,
            I => \N__33388\
        );

    \I__6035\ : Span4Mux_h
    port map (
            O => \N__33428\,
            I => \N__33385\
        );

    \I__6034\ : Span4Mux_v
    port map (
            O => \N__33425\,
            I => \N__33380\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__33416\,
            I => \N__33380\
        );

    \I__6032\ : Span4Mux_v
    port map (
            O => \N__33409\,
            I => \N__33375\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__33400\,
            I => \N__33375\
        );

    \I__6030\ : Span4Mux_v
    port map (
            O => \N__33395\,
            I => \N__33370\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__33392\,
            I => \N__33370\
        );

    \I__6028\ : CascadeMux
    port map (
            O => \N__33391\,
            I => \N__33367\
        );

    \I__6027\ : Span4Mux_v
    port map (
            O => \N__33388\,
            I => \N__33364\
        );

    \I__6026\ : Span4Mux_v
    port map (
            O => \N__33385\,
            I => \N__33361\
        );

    \I__6025\ : Span4Mux_v
    port map (
            O => \N__33380\,
            I => \N__33356\
        );

    \I__6024\ : Span4Mux_v
    port map (
            O => \N__33375\,
            I => \N__33356\
        );

    \I__6023\ : Span4Mux_v
    port map (
            O => \N__33370\,
            I => \N__33353\
        );

    \I__6022\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33350\
        );

    \I__6021\ : Span4Mux_h
    port map (
            O => \N__33364\,
            I => \N__33347\
        );

    \I__6020\ : Span4Mux_v
    port map (
            O => \N__33361\,
            I => \N__33344\
        );

    \I__6019\ : Span4Mux_h
    port map (
            O => \N__33356\,
            I => \N__33339\
        );

    \I__6018\ : Span4Mux_v
    port map (
            O => \N__33353\,
            I => \N__33339\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__33350\,
            I => \sEEPointerResetZ0\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__33347\,
            I => \sEEPointerResetZ0\
        );

    \I__6015\ : Odrv4
    port map (
            O => \N__33344\,
            I => \sEEPointerResetZ0\
        );

    \I__6014\ : Odrv4
    port map (
            O => \N__33339\,
            I => \sEEPointerResetZ0\
        );

    \I__6013\ : InMux
    port map (
            O => \N__33330\,
            I => \sRAM_pointer_write_cry_17\
        );

    \I__6012\ : InMux
    port map (
            O => \N__33327\,
            I => \N__33324\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__33324\,
            I => \N__33321\
        );

    \I__6010\ : Span4Mux_h
    port map (
            O => \N__33321\,
            I => \N__33317\
        );

    \I__6009\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33314\
        );

    \I__6008\ : Span4Mux_h
    port map (
            O => \N__33317\,
            I => \N__33311\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__33314\,
            I => \sRAM_pointer_writeZ0Z_18\
        );

    \I__6006\ : Odrv4
    port map (
            O => \N__33311\,
            I => \sRAM_pointer_writeZ0Z_18\
        );

    \I__6005\ : CEMux
    port map (
            O => \N__33306\,
            I => \N__33297\
        );

    \I__6004\ : CEMux
    port map (
            O => \N__33305\,
            I => \N__33297\
        );

    \I__6003\ : CEMux
    port map (
            O => \N__33304\,
            I => \N__33297\
        );

    \I__6002\ : GlobalMux
    port map (
            O => \N__33297\,
            I => \N__33294\
        );

    \I__6001\ : gio2CtrlBuf
    port map (
            O => \N__33294\,
            I => \N_26_g\
        );

    \I__6000\ : CascadeMux
    port map (
            O => \N__33291\,
            I => \N__33288\
        );

    \I__5999\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33278\
        );

    \I__5998\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33278\
        );

    \I__5997\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33278\
        );

    \I__5996\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33274\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__33278\,
            I => \N__33271\
        );

    \I__5994\ : InMux
    port map (
            O => \N__33277\,
            I => \N__33268\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__33274\,
            I => \N__33265\
        );

    \I__5992\ : Span4Mux_v
    port map (
            O => \N__33271\,
            I => \N__33262\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__33268\,
            I => \N__33259\
        );

    \I__5990\ : Span4Mux_h
    port map (
            O => \N__33265\,
            I => \N__33256\
        );

    \I__5989\ : Span4Mux_h
    port map (
            O => \N__33262\,
            I => \N__33251\
        );

    \I__5988\ : Span4Mux_v
    port map (
            O => \N__33259\,
            I => \N__33251\
        );

    \I__5987\ : Sp12to4
    port map (
            O => \N__33256\,
            I => \N__33248\
        );

    \I__5986\ : Span4Mux_v
    port map (
            O => \N__33251\,
            I => \N__33245\
        );

    \I__5985\ : Span12Mux_v
    port map (
            O => \N__33248\,
            I => \N__33240\
        );

    \I__5984\ : Sp12to4
    port map (
            O => \N__33245\,
            I => \N__33240\
        );

    \I__5983\ : Span12Mux_h
    port map (
            O => \N__33240\,
            I => \N__33237\
        );

    \I__5982\ : Odrv12
    port map (
            O => \N__33237\,
            I => spi_cs_ft_c
        );

    \I__5981\ : CascadeMux
    port map (
            O => \N__33234\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_\
        );

    \I__5980\ : InMux
    port map (
            O => \N__33231\,
            I => \N__33225\
        );

    \I__5979\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33225\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__33225\,
            I => \N__33218\
        );

    \I__5977\ : InMux
    port map (
            O => \N__33224\,
            I => \N__33215\
        );

    \I__5976\ : InMux
    port map (
            O => \N__33223\,
            I => \N__33206\
        );

    \I__5975\ : InMux
    port map (
            O => \N__33222\,
            I => \N__33206\
        );

    \I__5974\ : InMux
    port map (
            O => \N__33221\,
            I => \N__33206\
        );

    \I__5973\ : Span4Mux_v
    port map (
            O => \N__33218\,
            I => \N__33201\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__33215\,
            I => \N__33201\
        );

    \I__5971\ : InMux
    port map (
            O => \N__33214\,
            I => \N__33198\
        );

    \I__5970\ : InMux
    port map (
            O => \N__33213\,
            I => \N__33195\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__33206\,
            I => \N__33191\
        );

    \I__5968\ : Span4Mux_v
    port map (
            O => \N__33201\,
            I => \N__33186\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__33198\,
            I => \N__33186\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__33195\,
            I => \N__33183\
        );

    \I__5965\ : InMux
    port map (
            O => \N__33194\,
            I => \N__33180\
        );

    \I__5964\ : Span4Mux_v
    port map (
            O => \N__33191\,
            I => \N__33177\
        );

    \I__5963\ : Span4Mux_v
    port map (
            O => \N__33186\,
            I => \N__33172\
        );

    \I__5962\ : Span4Mux_v
    port map (
            O => \N__33183\,
            I => \N__33172\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__33180\,
            I => \N__33169\
        );

    \I__5960\ : Odrv4
    port map (
            O => \N__33177\,
            I => \spi_slave_inst.spi_csZ0\
        );

    \I__5959\ : Odrv4
    port map (
            O => \N__33172\,
            I => \spi_slave_inst.spi_csZ0\
        );

    \I__5958\ : Odrv4
    port map (
            O => \N__33169\,
            I => \spi_slave_inst.spi_csZ0\
        );

    \I__5957\ : CascadeMux
    port map (
            O => \N__33162\,
            I => \spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_\
        );

    \I__5956\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33156\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__33156\,
            I => \N__33153\
        );

    \I__5954\ : Span4Mux_h
    port map (
            O => \N__33153\,
            I => \N__33150\
        );

    \I__5953\ : Sp12to4
    port map (
            O => \N__33150\,
            I => \N__33146\
        );

    \I__5952\ : InMux
    port map (
            O => \N__33149\,
            I => \N__33143\
        );

    \I__5951\ : Odrv12
    port map (
            O => \N__33146\,
            I => \spi_slave_inst.tx_done_neg_sclk_iZ0\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__33143\,
            I => \spi_slave_inst.tx_done_neg_sclk_iZ0\
        );

    \I__5949\ : CascadeMux
    port map (
            O => \N__33138\,
            I => \N__33135\
        );

    \I__5948\ : InMux
    port map (
            O => \N__33135\,
            I => \N__33132\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__33132\,
            I => \N__33129\
        );

    \I__5946\ : Span12Mux_v
    port map (
            O => \N__33129\,
            I => \N__33126\
        );

    \I__5945\ : Span12Mux_h
    port map (
            O => \N__33126\,
            I => \N__33123\
        );

    \I__5944\ : Odrv12
    port map (
            O => \N__33123\,
            I => spi_miso_flash_c
        );

    \I__5943\ : IoInMux
    port map (
            O => \N__33120\,
            I => \N__33117\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__33117\,
            I => \N__33114\
        );

    \I__5941\ : IoSpan4Mux
    port map (
            O => \N__33114\,
            I => \N__33111\
        );

    \I__5940\ : Span4Mux_s2_h
    port map (
            O => \N__33111\,
            I => \N__33108\
        );

    \I__5939\ : Sp12to4
    port map (
            O => \N__33108\,
            I => \N__33105\
        );

    \I__5938\ : Span12Mux_s8_h
    port map (
            O => \N__33105\,
            I => \N__33102\
        );

    \I__5937\ : Odrv12
    port map (
            O => \N__33102\,
            I => spi_miso_rpi_c
        );

    \I__5936\ : CascadeMux
    port map (
            O => \N__33099\,
            I => \sDAC_data_2_13_bm_1_3_cascade_\
        );

    \I__5935\ : InMux
    port map (
            O => \N__33096\,
            I => \N__33093\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__33093\,
            I => \N__33089\
        );

    \I__5933\ : InMux
    port map (
            O => \N__33092\,
            I => \N__33086\
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__33089\,
            I => \sRAM_pointer_writeZ0Z_10\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__33086\,
            I => \sRAM_pointer_writeZ0Z_10\
        );

    \I__5930\ : InMux
    port map (
            O => \N__33081\,
            I => \sRAM_pointer_write_cry_9\
        );

    \I__5929\ : CascadeMux
    port map (
            O => \N__33078\,
            I => \N__33075\
        );

    \I__5928\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33072\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__33072\,
            I => \N__33068\
        );

    \I__5926\ : InMux
    port map (
            O => \N__33071\,
            I => \N__33065\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__33068\,
            I => \sRAM_pointer_writeZ0Z_11\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__33065\,
            I => \sRAM_pointer_writeZ0Z_11\
        );

    \I__5923\ : InMux
    port map (
            O => \N__33060\,
            I => \sRAM_pointer_write_cry_10\
        );

    \I__5922\ : InMux
    port map (
            O => \N__33057\,
            I => \N__33054\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__33054\,
            I => \N__33051\
        );

    \I__5920\ : Span4Mux_h
    port map (
            O => \N__33051\,
            I => \N__33047\
        );

    \I__5919\ : InMux
    port map (
            O => \N__33050\,
            I => \N__33044\
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__33047\,
            I => \sRAM_pointer_writeZ0Z_12\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__33044\,
            I => \sRAM_pointer_writeZ0Z_12\
        );

    \I__5916\ : InMux
    port map (
            O => \N__33039\,
            I => \sRAM_pointer_write_cry_11\
        );

    \I__5915\ : CascadeMux
    port map (
            O => \N__33036\,
            I => \N__33033\
        );

    \I__5914\ : InMux
    port map (
            O => \N__33033\,
            I => \N__33030\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__33030\,
            I => \N__33026\
        );

    \I__5912\ : InMux
    port map (
            O => \N__33029\,
            I => \N__33023\
        );

    \I__5911\ : Odrv4
    port map (
            O => \N__33026\,
            I => \sRAM_pointer_writeZ0Z_13\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__33023\,
            I => \sRAM_pointer_writeZ0Z_13\
        );

    \I__5909\ : InMux
    port map (
            O => \N__33018\,
            I => \sRAM_pointer_write_cry_12\
        );

    \I__5908\ : InMux
    port map (
            O => \N__33015\,
            I => \N__33012\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__33012\,
            I => \N__33009\
        );

    \I__5906\ : Span4Mux_h
    port map (
            O => \N__33009\,
            I => \N__33005\
        );

    \I__5905\ : InMux
    port map (
            O => \N__33008\,
            I => \N__33002\
        );

    \I__5904\ : Odrv4
    port map (
            O => \N__33005\,
            I => \sRAM_pointer_writeZ0Z_14\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__33002\,
            I => \sRAM_pointer_writeZ0Z_14\
        );

    \I__5902\ : InMux
    port map (
            O => \N__32997\,
            I => \sRAM_pointer_write_cry_13\
        );

    \I__5901\ : InMux
    port map (
            O => \N__32994\,
            I => \N__32991\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__32991\,
            I => \N__32988\
        );

    \I__5899\ : Span4Mux_h
    port map (
            O => \N__32988\,
            I => \N__32984\
        );

    \I__5898\ : InMux
    port map (
            O => \N__32987\,
            I => \N__32981\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__32984\,
            I => \sRAM_pointer_writeZ0Z_15\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__32981\,
            I => \sRAM_pointer_writeZ0Z_15\
        );

    \I__5895\ : InMux
    port map (
            O => \N__32976\,
            I => \sRAM_pointer_write_cry_14\
        );

    \I__5894\ : InMux
    port map (
            O => \N__32973\,
            I => \N__32970\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__32970\,
            I => \N__32966\
        );

    \I__5892\ : InMux
    port map (
            O => \N__32969\,
            I => \N__32963\
        );

    \I__5891\ : Span4Mux_v
    port map (
            O => \N__32966\,
            I => \N__32960\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__32963\,
            I => \sRAM_pointer_writeZ0Z_16\
        );

    \I__5889\ : Odrv4
    port map (
            O => \N__32960\,
            I => \sRAM_pointer_writeZ0Z_16\
        );

    \I__5888\ : InMux
    port map (
            O => \N__32955\,
            I => \bfn_13_20_0_\
        );

    \I__5887\ : InMux
    port map (
            O => \N__32952\,
            I => \N__32949\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__32949\,
            I => \N__32946\
        );

    \I__5885\ : Span4Mux_h
    port map (
            O => \N__32946\,
            I => \N__32943\
        );

    \I__5884\ : Span4Mux_h
    port map (
            O => \N__32943\,
            I => \N__32939\
        );

    \I__5883\ : InMux
    port map (
            O => \N__32942\,
            I => \N__32936\
        );

    \I__5882\ : Odrv4
    port map (
            O => \N__32939\,
            I => \sRAM_pointer_writeZ0Z_17\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__32936\,
            I => \sRAM_pointer_writeZ0Z_17\
        );

    \I__5880\ : InMux
    port map (
            O => \N__32931\,
            I => \sRAM_pointer_write_cry_16\
        );

    \I__5879\ : InMux
    port map (
            O => \N__32928\,
            I => \sRAM_pointer_write_cry_0\
        );

    \I__5878\ : InMux
    port map (
            O => \N__32925\,
            I => \N__32922\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__32922\,
            I => \N__32919\
        );

    \I__5876\ : Span4Mux_h
    port map (
            O => \N__32919\,
            I => \N__32915\
        );

    \I__5875\ : InMux
    port map (
            O => \N__32918\,
            I => \N__32912\
        );

    \I__5874\ : Odrv4
    port map (
            O => \N__32915\,
            I => \sRAM_pointer_writeZ0Z_2\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__32912\,
            I => \sRAM_pointer_writeZ0Z_2\
        );

    \I__5872\ : InMux
    port map (
            O => \N__32907\,
            I => \sRAM_pointer_write_cry_1\
        );

    \I__5871\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32901\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__32901\,
            I => \N__32898\
        );

    \I__5869\ : Span4Mux_h
    port map (
            O => \N__32898\,
            I => \N__32894\
        );

    \I__5868\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32891\
        );

    \I__5867\ : Odrv4
    port map (
            O => \N__32894\,
            I => \sRAM_pointer_writeZ0Z_3\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__32891\,
            I => \sRAM_pointer_writeZ0Z_3\
        );

    \I__5865\ : InMux
    port map (
            O => \N__32886\,
            I => \sRAM_pointer_write_cry_2\
        );

    \I__5864\ : InMux
    port map (
            O => \N__32883\,
            I => \N__32880\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__32880\,
            I => \N__32877\
        );

    \I__5862\ : Span4Mux_h
    port map (
            O => \N__32877\,
            I => \N__32874\
        );

    \I__5861\ : Span4Mux_h
    port map (
            O => \N__32874\,
            I => \N__32870\
        );

    \I__5860\ : InMux
    port map (
            O => \N__32873\,
            I => \N__32867\
        );

    \I__5859\ : Odrv4
    port map (
            O => \N__32870\,
            I => \sRAM_pointer_writeZ0Z_4\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__32867\,
            I => \sRAM_pointer_writeZ0Z_4\
        );

    \I__5857\ : InMux
    port map (
            O => \N__32862\,
            I => \sRAM_pointer_write_cry_3\
        );

    \I__5856\ : CascadeMux
    port map (
            O => \N__32859\,
            I => \N__32856\
        );

    \I__5855\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32853\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__32853\,
            I => \N__32849\
        );

    \I__5853\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32846\
        );

    \I__5852\ : Odrv4
    port map (
            O => \N__32849\,
            I => \sRAM_pointer_writeZ0Z_5\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__32846\,
            I => \sRAM_pointer_writeZ0Z_5\
        );

    \I__5850\ : InMux
    port map (
            O => \N__32841\,
            I => \sRAM_pointer_write_cry_4\
        );

    \I__5849\ : InMux
    port map (
            O => \N__32838\,
            I => \N__32835\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__32835\,
            I => \N__32831\
        );

    \I__5847\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32828\
        );

    \I__5846\ : Odrv4
    port map (
            O => \N__32831\,
            I => \sRAM_pointer_writeZ0Z_6\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__32828\,
            I => \sRAM_pointer_writeZ0Z_6\
        );

    \I__5844\ : InMux
    port map (
            O => \N__32823\,
            I => \sRAM_pointer_write_cry_5\
        );

    \I__5843\ : InMux
    port map (
            O => \N__32820\,
            I => \N__32817\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__32817\,
            I => \N__32813\
        );

    \I__5841\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32810\
        );

    \I__5840\ : Odrv4
    port map (
            O => \N__32813\,
            I => \sRAM_pointer_writeZ0Z_7\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__32810\,
            I => \sRAM_pointer_writeZ0Z_7\
        );

    \I__5838\ : InMux
    port map (
            O => \N__32805\,
            I => \sRAM_pointer_write_cry_6\
        );

    \I__5837\ : InMux
    port map (
            O => \N__32802\,
            I => \N__32799\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__32799\,
            I => \N__32796\
        );

    \I__5835\ : Span4Mux_v
    port map (
            O => \N__32796\,
            I => \N__32792\
        );

    \I__5834\ : InMux
    port map (
            O => \N__32795\,
            I => \N__32789\
        );

    \I__5833\ : Odrv4
    port map (
            O => \N__32792\,
            I => \sRAM_pointer_writeZ0Z_8\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__32789\,
            I => \sRAM_pointer_writeZ0Z_8\
        );

    \I__5831\ : InMux
    port map (
            O => \N__32784\,
            I => \bfn_13_19_0_\
        );

    \I__5830\ : InMux
    port map (
            O => \N__32781\,
            I => \N__32778\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__32778\,
            I => \N__32775\
        );

    \I__5828\ : Span4Mux_v
    port map (
            O => \N__32775\,
            I => \N__32772\
        );

    \I__5827\ : Span4Mux_h
    port map (
            O => \N__32772\,
            I => \N__32768\
        );

    \I__5826\ : InMux
    port map (
            O => \N__32771\,
            I => \N__32765\
        );

    \I__5825\ : Odrv4
    port map (
            O => \N__32768\,
            I => \sRAM_pointer_writeZ0Z_9\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__32765\,
            I => \sRAM_pointer_writeZ0Z_9\
        );

    \I__5823\ : InMux
    port map (
            O => \N__32760\,
            I => \sRAM_pointer_write_cry_8\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__32757\,
            I => \N_107_cascade_\
        );

    \I__5821\ : IoInMux
    port map (
            O => \N__32754\,
            I => \N__32751\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__32751\,
            I => \N__32748\
        );

    \I__5819\ : IoSpan4Mux
    port map (
            O => \N__32748\,
            I => \N__32745\
        );

    \I__5818\ : Span4Mux_s3_h
    port map (
            O => \N__32745\,
            I => \N__32742\
        );

    \I__5817\ : Sp12to4
    port map (
            O => \N__32742\,
            I => \N__32739\
        );

    \I__5816\ : Span12Mux_v
    port map (
            O => \N__32739\,
            I => \N__32736\
        );

    \I__5815\ : Span12Mux_h
    port map (
            O => \N__32736\,
            I => \N__32732\
        );

    \I__5814\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32729\
        );

    \I__5813\ : Odrv12
    port map (
            O => \N__32732\,
            I => \RAM_DATA_cl_5Z0Z_15\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__32729\,
            I => \RAM_DATA_cl_5Z0Z_15\
        );

    \I__5811\ : CascadeMux
    port map (
            O => \N__32724\,
            I => \N_108_cascade_\
        );

    \I__5810\ : IoInMux
    port map (
            O => \N__32721\,
            I => \N__32718\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__32718\,
            I => \N__32715\
        );

    \I__5808\ : IoSpan4Mux
    port map (
            O => \N__32715\,
            I => \N__32712\
        );

    \I__5807\ : IoSpan4Mux
    port map (
            O => \N__32712\,
            I => \N__32709\
        );

    \I__5806\ : Span4Mux_s3_h
    port map (
            O => \N__32709\,
            I => \N__32706\
        );

    \I__5805\ : Span4Mux_h
    port map (
            O => \N__32706\,
            I => \N__32703\
        );

    \I__5804\ : Span4Mux_h
    port map (
            O => \N__32703\,
            I => \N__32699\
        );

    \I__5803\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32696\
        );

    \I__5802\ : Odrv4
    port map (
            O => \N__32699\,
            I => \RAM_DATA_cl_6Z0Z_15\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__32696\,
            I => \RAM_DATA_cl_6Z0Z_15\
        );

    \I__5800\ : InMux
    port map (
            O => \N__32691\,
            I => \N__32672\
        );

    \I__5799\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32665\
        );

    \I__5798\ : InMux
    port map (
            O => \N__32689\,
            I => \N__32665\
        );

    \I__5797\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32665\
        );

    \I__5796\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32658\
        );

    \I__5795\ : InMux
    port map (
            O => \N__32686\,
            I => \N__32658\
        );

    \I__5794\ : InMux
    port map (
            O => \N__32685\,
            I => \N__32658\
        );

    \I__5793\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32649\
        );

    \I__5792\ : InMux
    port map (
            O => \N__32683\,
            I => \N__32649\
        );

    \I__5791\ : InMux
    port map (
            O => \N__32682\,
            I => \N__32649\
        );

    \I__5790\ : InMux
    port map (
            O => \N__32681\,
            I => \N__32649\
        );

    \I__5789\ : InMux
    port map (
            O => \N__32680\,
            I => \N__32640\
        );

    \I__5788\ : InMux
    port map (
            O => \N__32679\,
            I => \N__32640\
        );

    \I__5787\ : InMux
    port map (
            O => \N__32678\,
            I => \N__32640\
        );

    \I__5786\ : InMux
    port map (
            O => \N__32677\,
            I => \N__32640\
        );

    \I__5785\ : CascadeMux
    port map (
            O => \N__32676\,
            I => \N__32637\
        );

    \I__5784\ : CascadeMux
    port map (
            O => \N__32675\,
            I => \N__32628\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__32672\,
            I => \N__32625\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__32665\,
            I => \N__32614\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__32658\,
            I => \N__32614\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__32649\,
            I => \N__32614\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__32640\,
            I => \N__32614\
        );

    \I__5778\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32611\
        );

    \I__5777\ : InMux
    port map (
            O => \N__32636\,
            I => \N__32604\
        );

    \I__5776\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32604\
        );

    \I__5775\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32604\
        );

    \I__5774\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32599\
        );

    \I__5773\ : InMux
    port map (
            O => \N__32632\,
            I => \N__32599\
        );

    \I__5772\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32596\
        );

    \I__5771\ : InMux
    port map (
            O => \N__32628\,
            I => \N__32591\
        );

    \I__5770\ : Span4Mux_v
    port map (
            O => \N__32625\,
            I => \N__32587\
        );

    \I__5769\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32584\
        );

    \I__5768\ : CascadeMux
    port map (
            O => \N__32623\,
            I => \N__32580\
        );

    \I__5767\ : Span4Mux_v
    port map (
            O => \N__32614\,
            I => \N__32569\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__32611\,
            I => \N__32569\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__32604\,
            I => \N__32569\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__32599\,
            I => \N__32569\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__32596\,
            I => \N__32569\
        );

    \I__5762\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32566\
        );

    \I__5761\ : CascadeMux
    port map (
            O => \N__32594\,
            I => \N__32563\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__32591\,
            I => \N__32559\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__32590\,
            I => \N__32555\
        );

    \I__5758\ : Span4Mux_h
    port map (
            O => \N__32587\,
            I => \N__32551\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__32584\,
            I => \N__32548\
        );

    \I__5756\ : IoInMux
    port map (
            O => \N__32583\,
            I => \N__32543\
        );

    \I__5755\ : InMux
    port map (
            O => \N__32580\,
            I => \N__32540\
        );

    \I__5754\ : Span4Mux_v
    port map (
            O => \N__32569\,
            I => \N__32535\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__32566\,
            I => \N__32535\
        );

    \I__5752\ : InMux
    port map (
            O => \N__32563\,
            I => \N__32532\
        );

    \I__5751\ : InMux
    port map (
            O => \N__32562\,
            I => \N__32529\
        );

    \I__5750\ : Span4Mux_v
    port map (
            O => \N__32559\,
            I => \N__32526\
        );

    \I__5749\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32523\
        );

    \I__5748\ : InMux
    port map (
            O => \N__32555\,
            I => \N__32520\
        );

    \I__5747\ : CascadeMux
    port map (
            O => \N__32554\,
            I => \N__32517\
        );

    \I__5746\ : Span4Mux_h
    port map (
            O => \N__32551\,
            I => \N__32510\
        );

    \I__5745\ : Span4Mux_v
    port map (
            O => \N__32548\,
            I => \N__32510\
        );

    \I__5744\ : InMux
    port map (
            O => \N__32547\,
            I => \N__32507\
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__32546\,
            I => \N__32490\
        );

    \I__5742\ : LocalMux
    port map (
            O => \N__32543\,
            I => \N__32487\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__32540\,
            I => \N__32484\
        );

    \I__5740\ : Span4Mux_v
    port map (
            O => \N__32535\,
            I => \N__32479\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__32532\,
            I => \N__32479\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__32529\,
            I => \N__32476\
        );

    \I__5737\ : Span4Mux_v
    port map (
            O => \N__32526\,
            I => \N__32471\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__32523\,
            I => \N__32471\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__32520\,
            I => \N__32463\
        );

    \I__5734\ : InMux
    port map (
            O => \N__32517\,
            I => \N__32456\
        );

    \I__5733\ : InMux
    port map (
            O => \N__32516\,
            I => \N__32456\
        );

    \I__5732\ : CEMux
    port map (
            O => \N__32515\,
            I => \N__32456\
        );

    \I__5731\ : Span4Mux_v
    port map (
            O => \N__32510\,
            I => \N__32451\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__32507\,
            I => \N__32451\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__32506\,
            I => \N__32448\
        );

    \I__5728\ : CascadeMux
    port map (
            O => \N__32505\,
            I => \N__32445\
        );

    \I__5727\ : CascadeMux
    port map (
            O => \N__32504\,
            I => \N__32441\
        );

    \I__5726\ : InMux
    port map (
            O => \N__32503\,
            I => \N__32434\
        );

    \I__5725\ : InMux
    port map (
            O => \N__32502\,
            I => \N__32434\
        );

    \I__5724\ : InMux
    port map (
            O => \N__32501\,
            I => \N__32434\
        );

    \I__5723\ : InMux
    port map (
            O => \N__32500\,
            I => \N__32423\
        );

    \I__5722\ : InMux
    port map (
            O => \N__32499\,
            I => \N__32423\
        );

    \I__5721\ : InMux
    port map (
            O => \N__32498\,
            I => \N__32423\
        );

    \I__5720\ : InMux
    port map (
            O => \N__32497\,
            I => \N__32423\
        );

    \I__5719\ : InMux
    port map (
            O => \N__32496\,
            I => \N__32423\
        );

    \I__5718\ : InMux
    port map (
            O => \N__32495\,
            I => \N__32414\
        );

    \I__5717\ : InMux
    port map (
            O => \N__32494\,
            I => \N__32414\
        );

    \I__5716\ : InMux
    port map (
            O => \N__32493\,
            I => \N__32414\
        );

    \I__5715\ : InMux
    port map (
            O => \N__32490\,
            I => \N__32414\
        );

    \I__5714\ : Span4Mux_s2_h
    port map (
            O => \N__32487\,
            I => \N__32410\
        );

    \I__5713\ : Span4Mux_v
    port map (
            O => \N__32484\,
            I => \N__32407\
        );

    \I__5712\ : Span4Mux_v
    port map (
            O => \N__32479\,
            I => \N__32404\
        );

    \I__5711\ : Span4Mux_h
    port map (
            O => \N__32476\,
            I => \N__32399\
        );

    \I__5710\ : Span4Mux_v
    port map (
            O => \N__32471\,
            I => \N__32399\
        );

    \I__5709\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32391\
        );

    \I__5708\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32391\
        );

    \I__5707\ : InMux
    port map (
            O => \N__32468\,
            I => \N__32391\
        );

    \I__5706\ : InMux
    port map (
            O => \N__32467\,
            I => \N__32386\
        );

    \I__5705\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32386\
        );

    \I__5704\ : Span4Mux_v
    port map (
            O => \N__32463\,
            I => \N__32383\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__32456\,
            I => \N__32380\
        );

    \I__5702\ : Span4Mux_v
    port map (
            O => \N__32451\,
            I => \N__32377\
        );

    \I__5701\ : InMux
    port map (
            O => \N__32448\,
            I => \N__32372\
        );

    \I__5700\ : InMux
    port map (
            O => \N__32445\,
            I => \N__32372\
        );

    \I__5699\ : InMux
    port map (
            O => \N__32444\,
            I => \N__32367\
        );

    \I__5698\ : InMux
    port map (
            O => \N__32441\,
            I => \N__32367\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__32434\,
            I => \N__32364\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__32423\,
            I => \N__32361\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__32414\,
            I => \N__32358\
        );

    \I__5694\ : InMux
    port map (
            O => \N__32413\,
            I => \N__32355\
        );

    \I__5693\ : Sp12to4
    port map (
            O => \N__32410\,
            I => \N__32347\
        );

    \I__5692\ : Span4Mux_h
    port map (
            O => \N__32407\,
            I => \N__32340\
        );

    \I__5691\ : Span4Mux_h
    port map (
            O => \N__32404\,
            I => \N__32340\
        );

    \I__5690\ : Span4Mux_v
    port map (
            O => \N__32399\,
            I => \N__32340\
        );

    \I__5689\ : InMux
    port map (
            O => \N__32398\,
            I => \N__32337\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__32391\,
            I => \N__32332\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__32386\,
            I => \N__32332\
        );

    \I__5686\ : Span4Mux_h
    port map (
            O => \N__32383\,
            I => \N__32327\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__32380\,
            I => \N__32327\
        );

    \I__5684\ : Span4Mux_v
    port map (
            O => \N__32377\,
            I => \N__32323\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__32372\,
            I => \N__32318\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__32367\,
            I => \N__32318\
        );

    \I__5681\ : Span4Mux_v
    port map (
            O => \N__32364\,
            I => \N__32309\
        );

    \I__5680\ : Span4Mux_h
    port map (
            O => \N__32361\,
            I => \N__32309\
        );

    \I__5679\ : Span4Mux_h
    port map (
            O => \N__32358\,
            I => \N__32309\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__32355\,
            I => \N__32309\
        );

    \I__5677\ : InMux
    port map (
            O => \N__32354\,
            I => \N__32302\
        );

    \I__5676\ : InMux
    port map (
            O => \N__32353\,
            I => \N__32302\
        );

    \I__5675\ : InMux
    port map (
            O => \N__32352\,
            I => \N__32302\
        );

    \I__5674\ : InMux
    port map (
            O => \N__32351\,
            I => \N__32299\
        );

    \I__5673\ : InMux
    port map (
            O => \N__32350\,
            I => \N__32296\
        );

    \I__5672\ : Span12Mux_v
    port map (
            O => \N__32347\,
            I => \N__32293\
        );

    \I__5671\ : Span4Mux_v
    port map (
            O => \N__32340\,
            I => \N__32290\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__32337\,
            I => \N__32287\
        );

    \I__5669\ : Span4Mux_v
    port map (
            O => \N__32332\,
            I => \N__32282\
        );

    \I__5668\ : Span4Mux_v
    port map (
            O => \N__32327\,
            I => \N__32282\
        );

    \I__5667\ : IoInMux
    port map (
            O => \N__32326\,
            I => \N__32279\
        );

    \I__5666\ : Sp12to4
    port map (
            O => \N__32323\,
            I => \N__32276\
        );

    \I__5665\ : Span12Mux_s9_v
    port map (
            O => \N__32318\,
            I => \N__32265\
        );

    \I__5664\ : Sp12to4
    port map (
            O => \N__32309\,
            I => \N__32265\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__32302\,
            I => \N__32265\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__32299\,
            I => \N__32265\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__32296\,
            I => \N__32265\
        );

    \I__5660\ : Span12Mux_v
    port map (
            O => \N__32293\,
            I => \N__32262\
        );

    \I__5659\ : Sp12to4
    port map (
            O => \N__32290\,
            I => \N__32259\
        );

    \I__5658\ : Sp12to4
    port map (
            O => \N__32287\,
            I => \N__32254\
        );

    \I__5657\ : Sp12to4
    port map (
            O => \N__32282\,
            I => \N__32254\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__32279\,
            I => \N__32251\
        );

    \I__5655\ : Span12Mux_h
    port map (
            O => \N__32276\,
            I => \N__32246\
        );

    \I__5654\ : Span12Mux_v
    port map (
            O => \N__32265\,
            I => \N__32246\
        );

    \I__5653\ : Span12Mux_h
    port map (
            O => \N__32262\,
            I => \N__32239\
        );

    \I__5652\ : Span12Mux_h
    port map (
            O => \N__32259\,
            I => \N__32239\
        );

    \I__5651\ : Span12Mux_v
    port map (
            O => \N__32254\,
            I => \N__32239\
        );

    \I__5650\ : IoSpan4Mux
    port map (
            O => \N__32251\,
            I => \N__32236\
        );

    \I__5649\ : Odrv12
    port map (
            O => \N__32246\,
            I => \LED3_c\
        );

    \I__5648\ : Odrv12
    port map (
            O => \N__32239\,
            I => \LED3_c\
        );

    \I__5647\ : Odrv4
    port map (
            O => \N__32236\,
            I => \LED3_c\
        );

    \I__5646\ : CascadeMux
    port map (
            O => \N__32229\,
            I => \N__32208\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__32228\,
            I => \N__32205\
        );

    \I__5644\ : CascadeMux
    port map (
            O => \N__32227\,
            I => \N__32202\
        );

    \I__5643\ : CascadeMux
    port map (
            O => \N__32226\,
            I => \N__32199\
        );

    \I__5642\ : InMux
    port map (
            O => \N__32225\,
            I => \N__32187\
        );

    \I__5641\ : InMux
    port map (
            O => \N__32224\,
            I => \N__32187\
        );

    \I__5640\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32187\
        );

    \I__5639\ : InMux
    port map (
            O => \N__32222\,
            I => \N__32187\
        );

    \I__5638\ : CascadeMux
    port map (
            O => \N__32221\,
            I => \N__32172\
        );

    \I__5637\ : CascadeMux
    port map (
            O => \N__32220\,
            I => \N__32169\
        );

    \I__5636\ : CascadeMux
    port map (
            O => \N__32219\,
            I => \N__32166\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__32218\,
            I => \N__32160\
        );

    \I__5634\ : InMux
    port map (
            O => \N__32217\,
            I => \N__32154\
        );

    \I__5633\ : InMux
    port map (
            O => \N__32216\,
            I => \N__32154\
        );

    \I__5632\ : InMux
    port map (
            O => \N__32215\,
            I => \N__32148\
        );

    \I__5631\ : InMux
    port map (
            O => \N__32214\,
            I => \N__32141\
        );

    \I__5630\ : InMux
    port map (
            O => \N__32213\,
            I => \N__32141\
        );

    \I__5629\ : InMux
    port map (
            O => \N__32212\,
            I => \N__32141\
        );

    \I__5628\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32138\
        );

    \I__5627\ : InMux
    port map (
            O => \N__32208\,
            I => \N__32123\
        );

    \I__5626\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32123\
        );

    \I__5625\ : InMux
    port map (
            O => \N__32202\,
            I => \N__32123\
        );

    \I__5624\ : InMux
    port map (
            O => \N__32199\,
            I => \N__32123\
        );

    \I__5623\ : InMux
    port map (
            O => \N__32198\,
            I => \N__32123\
        );

    \I__5622\ : InMux
    port map (
            O => \N__32197\,
            I => \N__32123\
        );

    \I__5621\ : InMux
    port map (
            O => \N__32196\,
            I => \N__32123\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__32187\,
            I => \N__32120\
        );

    \I__5619\ : InMux
    port map (
            O => \N__32186\,
            I => \N__32103\
        );

    \I__5618\ : InMux
    port map (
            O => \N__32185\,
            I => \N__32103\
        );

    \I__5617\ : InMux
    port map (
            O => \N__32184\,
            I => \N__32103\
        );

    \I__5616\ : InMux
    port map (
            O => \N__32183\,
            I => \N__32103\
        );

    \I__5615\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32103\
        );

    \I__5614\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32103\
        );

    \I__5613\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32103\
        );

    \I__5612\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32103\
        );

    \I__5611\ : CascadeMux
    port map (
            O => \N__32178\,
            I => \N__32099\
        );

    \I__5610\ : InMux
    port map (
            O => \N__32177\,
            I => \N__32094\
        );

    \I__5609\ : InMux
    port map (
            O => \N__32176\,
            I => \N__32094\
        );

    \I__5608\ : InMux
    port map (
            O => \N__32175\,
            I => \N__32091\
        );

    \I__5607\ : InMux
    port map (
            O => \N__32172\,
            I => \N__32088\
        );

    \I__5606\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32077\
        );

    \I__5605\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32077\
        );

    \I__5604\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32077\
        );

    \I__5603\ : InMux
    port map (
            O => \N__32164\,
            I => \N__32077\
        );

    \I__5602\ : InMux
    port map (
            O => \N__32163\,
            I => \N__32077\
        );

    \I__5601\ : InMux
    port map (
            O => \N__32160\,
            I => \N__32072\
        );

    \I__5600\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32072\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__32154\,
            I => \N__32069\
        );

    \I__5598\ : InMux
    port map (
            O => \N__32153\,
            I => \N__32063\
        );

    \I__5597\ : InMux
    port map (
            O => \N__32152\,
            I => \N__32058\
        );

    \I__5596\ : InMux
    port map (
            O => \N__32151\,
            I => \N__32058\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__32148\,
            I => \N__32055\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__32141\,
            I => \N__32052\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__32138\,
            I => \N__32049\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__32123\,
            I => \N__32042\
        );

    \I__5591\ : Span4Mux_h
    port map (
            O => \N__32120\,
            I => \N__32042\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32042\
        );

    \I__5589\ : InMux
    port map (
            O => \N__32102\,
            I => \N__32037\
        );

    \I__5588\ : InMux
    port map (
            O => \N__32099\,
            I => \N__32037\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__32094\,
            I => \N__32032\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__32091\,
            I => \N__32032\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__32088\,
            I => \N__32023\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__32077\,
            I => \N__32023\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__32072\,
            I => \N__32023\
        );

    \I__5582\ : Span4Mux_v
    port map (
            O => \N__32069\,
            I => \N__32023\
        );

    \I__5581\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32016\
        );

    \I__5580\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32016\
        );

    \I__5579\ : InMux
    port map (
            O => \N__32066\,
            I => \N__32016\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__32063\,
            I => \N__32009\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__32058\,
            I => \N__32009\
        );

    \I__5576\ : Span12Mux_v
    port map (
            O => \N__32055\,
            I => \N__32009\
        );

    \I__5575\ : Span4Mux_h
    port map (
            O => \N__32052\,
            I => \N__32004\
        );

    \I__5574\ : Span4Mux_h
    port map (
            O => \N__32049\,
            I => \N__32004\
        );

    \I__5573\ : Span4Mux_h
    port map (
            O => \N__32042\,
            I => \N__32001\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__32037\,
            I => \N__31998\
        );

    \I__5571\ : Span4Mux_v
    port map (
            O => \N__32032\,
            I => \N__31993\
        );

    \I__5570\ : Span4Mux_v
    port map (
            O => \N__32023\,
            I => \N__31993\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__32016\,
            I => \un4_sacqtime_cry_23_THRU_CO\
        );

    \I__5568\ : Odrv12
    port map (
            O => \N__32009\,
            I => \un4_sacqtime_cry_23_THRU_CO\
        );

    \I__5567\ : Odrv4
    port map (
            O => \N__32004\,
            I => \un4_sacqtime_cry_23_THRU_CO\
        );

    \I__5566\ : Odrv4
    port map (
            O => \N__32001\,
            I => \un4_sacqtime_cry_23_THRU_CO\
        );

    \I__5565\ : Odrv4
    port map (
            O => \N__31998\,
            I => \un4_sacqtime_cry_23_THRU_CO\
        );

    \I__5564\ : Odrv4
    port map (
            O => \N__31993\,
            I => \un4_sacqtime_cry_23_THRU_CO\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__31980\,
            I => \N_95_cascade_\
        );

    \I__5562\ : InMux
    port map (
            O => \N__31977\,
            I => \N__31974\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__31974\,
            I => \N__31970\
        );

    \I__5560\ : InMux
    port map (
            O => \N__31973\,
            I => \N__31952\
        );

    \I__5559\ : Span4Mux_h
    port map (
            O => \N__31970\,
            I => \N__31949\
        );

    \I__5558\ : InMux
    port map (
            O => \N__31969\,
            I => \N__31927\
        );

    \I__5557\ : InMux
    port map (
            O => \N__31968\,
            I => \N__31927\
        );

    \I__5556\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31927\
        );

    \I__5555\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31922\
        );

    \I__5554\ : InMux
    port map (
            O => \N__31965\,
            I => \N__31922\
        );

    \I__5553\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31917\
        );

    \I__5552\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31917\
        );

    \I__5551\ : InMux
    port map (
            O => \N__31962\,
            I => \N__31897\
        );

    \I__5550\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31897\
        );

    \I__5549\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31897\
        );

    \I__5548\ : InMux
    port map (
            O => \N__31959\,
            I => \N__31897\
        );

    \I__5547\ : InMux
    port map (
            O => \N__31958\,
            I => \N__31897\
        );

    \I__5546\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31897\
        );

    \I__5545\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31892\
        );

    \I__5544\ : InMux
    port map (
            O => \N__31955\,
            I => \N__31892\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__31952\,
            I => \N__31889\
        );

    \I__5542\ : Span4Mux_v
    port map (
            O => \N__31949\,
            I => \N__31886\
        );

    \I__5541\ : InMux
    port map (
            O => \N__31948\,
            I => \N__31873\
        );

    \I__5540\ : InMux
    port map (
            O => \N__31947\,
            I => \N__31873\
        );

    \I__5539\ : InMux
    port map (
            O => \N__31946\,
            I => \N__31873\
        );

    \I__5538\ : InMux
    port map (
            O => \N__31945\,
            I => \N__31873\
        );

    \I__5537\ : InMux
    port map (
            O => \N__31944\,
            I => \N__31866\
        );

    \I__5536\ : InMux
    port map (
            O => \N__31943\,
            I => \N__31866\
        );

    \I__5535\ : InMux
    port map (
            O => \N__31942\,
            I => \N__31866\
        );

    \I__5534\ : InMux
    port map (
            O => \N__31941\,
            I => \N__31849\
        );

    \I__5533\ : InMux
    port map (
            O => \N__31940\,
            I => \N__31849\
        );

    \I__5532\ : InMux
    port map (
            O => \N__31939\,
            I => \N__31849\
        );

    \I__5531\ : InMux
    port map (
            O => \N__31938\,
            I => \N__31849\
        );

    \I__5530\ : InMux
    port map (
            O => \N__31937\,
            I => \N__31849\
        );

    \I__5529\ : InMux
    port map (
            O => \N__31936\,
            I => \N__31849\
        );

    \I__5528\ : InMux
    port map (
            O => \N__31935\,
            I => \N__31849\
        );

    \I__5527\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31849\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__31927\,
            I => \N__31840\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__31922\,
            I => \N__31840\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__31917\,
            I => \N__31840\
        );

    \I__5523\ : InMux
    port map (
            O => \N__31916\,
            I => \N__31835\
        );

    \I__5522\ : InMux
    port map (
            O => \N__31915\,
            I => \N__31835\
        );

    \I__5521\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31824\
        );

    \I__5520\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31824\
        );

    \I__5519\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31824\
        );

    \I__5518\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31824\
        );

    \I__5517\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31824\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__31897\,
            I => \N__31817\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__31892\,
            I => \N__31817\
        );

    \I__5514\ : Span4Mux_v
    port map (
            O => \N__31889\,
            I => \N__31817\
        );

    \I__5513\ : Span4Mux_h
    port map (
            O => \N__31886\,
            I => \N__31814\
        );

    \I__5512\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31805\
        );

    \I__5511\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31805\
        );

    \I__5510\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31805\
        );

    \I__5509\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31805\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__31873\,
            I => \N__31798\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__31866\,
            I => \N__31798\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__31849\,
            I => \N__31798\
        );

    \I__5505\ : InMux
    port map (
            O => \N__31848\,
            I => \N__31793\
        );

    \I__5504\ : InMux
    port map (
            O => \N__31847\,
            I => \N__31793\
        );

    \I__5503\ : Span4Mux_v
    port map (
            O => \N__31840\,
            I => \N__31788\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__31835\,
            I => \N__31788\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__31824\,
            I => \un1_sacqtime_cry_23_THRU_CO\
        );

    \I__5500\ : Odrv4
    port map (
            O => \N__31817\,
            I => \un1_sacqtime_cry_23_THRU_CO\
        );

    \I__5499\ : Odrv4
    port map (
            O => \N__31814\,
            I => \un1_sacqtime_cry_23_THRU_CO\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__31805\,
            I => \un1_sacqtime_cry_23_THRU_CO\
        );

    \I__5497\ : Odrv12
    port map (
            O => \N__31798\,
            I => \un1_sacqtime_cry_23_THRU_CO\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__31793\,
            I => \un1_sacqtime_cry_23_THRU_CO\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__31788\,
            I => \un1_sacqtime_cry_23_THRU_CO\
        );

    \I__5494\ : IoInMux
    port map (
            O => \N__31773\,
            I => \N__31770\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__31770\,
            I => \N__31767\
        );

    \I__5492\ : IoSpan4Mux
    port map (
            O => \N__31767\,
            I => \N__31764\
        );

    \I__5491\ : Span4Mux_s2_h
    port map (
            O => \N__31764\,
            I => \N__31761\
        );

    \I__5490\ : Sp12to4
    port map (
            O => \N__31761\,
            I => \N__31758\
        );

    \I__5489\ : Span12Mux_h
    port map (
            O => \N__31758\,
            I => \N__31754\
        );

    \I__5488\ : InMux
    port map (
            O => \N__31757\,
            I => \N__31751\
        );

    \I__5487\ : Odrv12
    port map (
            O => \N__31754\,
            I => \RAM_DATA_cl_7Z0Z_15\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__31751\,
            I => \RAM_DATA_cl_7Z0Z_15\
        );

    \I__5485\ : IoInMux
    port map (
            O => \N__31746\,
            I => \N__31743\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__31743\,
            I => \N__31740\
        );

    \I__5483\ : IoSpan4Mux
    port map (
            O => \N__31740\,
            I => \N__31737\
        );

    \I__5482\ : IoSpan4Mux
    port map (
            O => \N__31737\,
            I => \N__31734\
        );

    \I__5481\ : Span4Mux_s2_h
    port map (
            O => \N__31734\,
            I => \N__31731\
        );

    \I__5480\ : Sp12to4
    port map (
            O => \N__31731\,
            I => \N__31728\
        );

    \I__5479\ : Span12Mux_h
    port map (
            O => \N__31728\,
            I => \N__31725\
        );

    \I__5478\ : Span12Mux_v
    port map (
            O => \N__31725\,
            I => \N__31721\
        );

    \I__5477\ : InMux
    port map (
            O => \N__31724\,
            I => \N__31718\
        );

    \I__5476\ : Odrv12
    port map (
            O => \N__31721\,
            I => \RAM_DATA_cl_4Z0Z_15\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__31718\,
            I => \RAM_DATA_cl_4Z0Z_15\
        );

    \I__5474\ : InMux
    port map (
            O => \N__31713\,
            I => \N__31698\
        );

    \I__5473\ : InMux
    port map (
            O => \N__31712\,
            I => \N__31698\
        );

    \I__5472\ : InMux
    port map (
            O => \N__31711\,
            I => \N__31698\
        );

    \I__5471\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31698\
        );

    \I__5470\ : InMux
    port map (
            O => \N__31709\,
            I => \N__31686\
        );

    \I__5469\ : InMux
    port map (
            O => \N__31708\,
            I => \N__31686\
        );

    \I__5468\ : InMux
    port map (
            O => \N__31707\,
            I => \N__31686\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__31698\,
            I => \N__31680\
        );

    \I__5466\ : InMux
    port map (
            O => \N__31697\,
            I => \N__31671\
        );

    \I__5465\ : InMux
    port map (
            O => \N__31696\,
            I => \N__31671\
        );

    \I__5464\ : InMux
    port map (
            O => \N__31695\,
            I => \N__31671\
        );

    \I__5463\ : InMux
    port map (
            O => \N__31694\,
            I => \N__31671\
        );

    \I__5462\ : InMux
    port map (
            O => \N__31693\,
            I => \N__31666\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__31686\,
            I => \N__31663\
        );

    \I__5460\ : InMux
    port map (
            O => \N__31685\,
            I => \N__31656\
        );

    \I__5459\ : InMux
    port map (
            O => \N__31684\,
            I => \N__31656\
        );

    \I__5458\ : InMux
    port map (
            O => \N__31683\,
            I => \N__31656\
        );

    \I__5457\ : Span4Mux_h
    port map (
            O => \N__31680\,
            I => \N__31653\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__31671\,
            I => \N__31650\
        );

    \I__5455\ : InMux
    port map (
            O => \N__31670\,
            I => \N__31645\
        );

    \I__5454\ : InMux
    port map (
            O => \N__31669\,
            I => \N__31645\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__31666\,
            I => \N__31642\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__31663\,
            I => \N_71\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__31656\,
            I => \N_71\
        );

    \I__5450\ : Odrv4
    port map (
            O => \N__31653\,
            I => \N_71\
        );

    \I__5449\ : Odrv4
    port map (
            O => \N__31650\,
            I => \N_71\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__31645\,
            I => \N_71\
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__31642\,
            I => \N_71\
        );

    \I__5446\ : InMux
    port map (
            O => \N__31629\,
            I => \N__31626\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__31626\,
            I => \N_105\
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__31623\,
            I => \N__31620\
        );

    \I__5443\ : InMux
    port map (
            O => \N__31620\,
            I => \N__31616\
        );

    \I__5442\ : InMux
    port map (
            O => \N__31619\,
            I => \N__31613\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__31616\,
            I => \sRAM_pointer_writeZ0Z_0\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__31613\,
            I => \sRAM_pointer_writeZ0Z_0\
        );

    \I__5439\ : InMux
    port map (
            O => \N__31608\,
            I => \bfn_13_18_0_\
        );

    \I__5438\ : CascadeMux
    port map (
            O => \N__31605\,
            I => \N__31602\
        );

    \I__5437\ : InMux
    port map (
            O => \N__31602\,
            I => \N__31598\
        );

    \I__5436\ : InMux
    port map (
            O => \N__31601\,
            I => \N__31595\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__31598\,
            I => \sRAM_pointer_writeZ0Z_1\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__31595\,
            I => \sRAM_pointer_writeZ0Z_1\
        );

    \I__5433\ : InMux
    port map (
            O => \N__31590\,
            I => \N__31587\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__31587\,
            I => \N__31584\
        );

    \I__5431\ : Sp12to4
    port map (
            O => \N__31584\,
            I => \N__31581\
        );

    \I__5430\ : Span12Mux_v
    port map (
            O => \N__31581\,
            I => \N__31578\
        );

    \I__5429\ : Span12Mux_h
    port map (
            O => \N__31578\,
            I => \N__31575\
        );

    \I__5428\ : Odrv12
    port map (
            O => \N__31575\,
            I => \ADC4_c\
        );

    \I__5427\ : IoInMux
    port map (
            O => \N__31572\,
            I => \N__31569\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__31569\,
            I => \N__31566\
        );

    \I__5425\ : Span4Mux_s2_v
    port map (
            O => \N__31566\,
            I => \N__31563\
        );

    \I__5424\ : Sp12to4
    port map (
            O => \N__31563\,
            I => \N__31560\
        );

    \I__5423\ : Span12Mux_h
    port map (
            O => \N__31560\,
            I => \N__31557\
        );

    \I__5422\ : Odrv12
    port map (
            O => \N__31557\,
            I => \RAM_DATA_1Z0Z_4\
        );

    \I__5421\ : InMux
    port map (
            O => \N__31554\,
            I => \N__31551\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__31551\,
            I => \N__31548\
        );

    \I__5419\ : Span12Mux_s11_v
    port map (
            O => \N__31548\,
            I => \N__31545\
        );

    \I__5418\ : Span12Mux_h
    port map (
            O => \N__31545\,
            I => \N__31542\
        );

    \I__5417\ : Odrv12
    port map (
            O => \N__31542\,
            I => \ADC6_c\
        );

    \I__5416\ : IoInMux
    port map (
            O => \N__31539\,
            I => \N__31536\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__31536\,
            I => \N__31533\
        );

    \I__5414\ : Span4Mux_s1_v
    port map (
            O => \N__31533\,
            I => \N__31530\
        );

    \I__5413\ : Sp12to4
    port map (
            O => \N__31530\,
            I => \N__31527\
        );

    \I__5412\ : Span12Mux_h
    port map (
            O => \N__31527\,
            I => \N__31524\
        );

    \I__5411\ : Odrv12
    port map (
            O => \N__31524\,
            I => \RAM_DATA_1Z0Z_6\
        );

    \I__5410\ : InMux
    port map (
            O => \N__31521\,
            I => \N__31518\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__31518\,
            I => \N__31515\
        );

    \I__5408\ : Span4Mux_v
    port map (
            O => \N__31515\,
            I => \N__31512\
        );

    \I__5407\ : Sp12to4
    port map (
            O => \N__31512\,
            I => \N__31509\
        );

    \I__5406\ : Span12Mux_h
    port map (
            O => \N__31509\,
            I => \N__31506\
        );

    \I__5405\ : Span12Mux_h
    port map (
            O => \N__31506\,
            I => \N__31503\
        );

    \I__5404\ : Odrv12
    port map (
            O => \N__31503\,
            I => \ADC9_c\
        );

    \I__5403\ : IoInMux
    port map (
            O => \N__31500\,
            I => \N__31497\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__31497\,
            I => \N__31494\
        );

    \I__5401\ : Span4Mux_s3_h
    port map (
            O => \N__31494\,
            I => \N__31491\
        );

    \I__5400\ : Sp12to4
    port map (
            O => \N__31491\,
            I => \N__31488\
        );

    \I__5399\ : Span12Mux_s7_v
    port map (
            O => \N__31488\,
            I => \N__31485\
        );

    \I__5398\ : Span12Mux_h
    port map (
            O => \N__31485\,
            I => \N__31482\
        );

    \I__5397\ : Span12Mux_v
    port map (
            O => \N__31482\,
            I => \N__31479\
        );

    \I__5396\ : Odrv12
    port map (
            O => \N__31479\,
            I => \RAM_DATA_1Z0Z_10\
        );

    \I__5395\ : InMux
    port map (
            O => \N__31476\,
            I => \N__31473\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__31473\,
            I => \N__31470\
        );

    \I__5393\ : Span4Mux_v
    port map (
            O => \N__31470\,
            I => \N__31467\
        );

    \I__5392\ : Sp12to4
    port map (
            O => \N__31467\,
            I => \N__31464\
        );

    \I__5391\ : Span12Mux_h
    port map (
            O => \N__31464\,
            I => \N__31461\
        );

    \I__5390\ : Span12Mux_v
    port map (
            O => \N__31461\,
            I => \N__31458\
        );

    \I__5389\ : Odrv12
    port map (
            O => \N__31458\,
            I => top_tour1_c
        );

    \I__5388\ : IoInMux
    port map (
            O => \N__31455\,
            I => \N__31452\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__31452\,
            I => \N__31449\
        );

    \I__5386\ : IoSpan4Mux
    port map (
            O => \N__31449\,
            I => \N__31446\
        );

    \I__5385\ : Span4Mux_s1_h
    port map (
            O => \N__31446\,
            I => \N__31443\
        );

    \I__5384\ : Sp12to4
    port map (
            O => \N__31443\,
            I => \N__31440\
        );

    \I__5383\ : Span12Mux_h
    port map (
            O => \N__31440\,
            I => \N__31437\
        );

    \I__5382\ : Odrv12
    port map (
            O => \N__31437\,
            I => \RAM_DATA_1Z0Z_11\
        );

    \I__5381\ : InMux
    port map (
            O => \N__31434\,
            I => \N__31431\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__31431\,
            I => \N__31428\
        );

    \I__5379\ : Sp12to4
    port map (
            O => \N__31428\,
            I => \N__31425\
        );

    \I__5378\ : Span12Mux_s9_v
    port map (
            O => \N__31425\,
            I => \N__31422\
        );

    \I__5377\ : Span12Mux_v
    port map (
            O => \N__31422\,
            I => \N__31419\
        );

    \I__5376\ : Span12Mux_h
    port map (
            O => \N__31419\,
            I => \N__31416\
        );

    \I__5375\ : Odrv12
    port map (
            O => \N__31416\,
            I => top_tour2_c
        );

    \I__5374\ : IoInMux
    port map (
            O => \N__31413\,
            I => \N__31410\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__31410\,
            I => \N__31407\
        );

    \I__5372\ : IoSpan4Mux
    port map (
            O => \N__31407\,
            I => \N__31404\
        );

    \I__5371\ : IoSpan4Mux
    port map (
            O => \N__31404\,
            I => \N__31401\
        );

    \I__5370\ : Span4Mux_s2_h
    port map (
            O => \N__31401\,
            I => \N__31398\
        );

    \I__5369\ : Sp12to4
    port map (
            O => \N__31398\,
            I => \N__31395\
        );

    \I__5368\ : Odrv12
    port map (
            O => \N__31395\,
            I => \RAM_DATA_1Z0Z_12\
        );

    \I__5367\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31380\
        );

    \I__5366\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31380\
        );

    \I__5365\ : InMux
    port map (
            O => \N__31390\,
            I => \N__31380\
        );

    \I__5364\ : InMux
    port map (
            O => \N__31389\,
            I => \N__31376\
        );

    \I__5363\ : InMux
    port map (
            O => \N__31388\,
            I => \N__31373\
        );

    \I__5362\ : InMux
    port map (
            O => \N__31387\,
            I => \N__31370\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__31380\,
            I => \N__31367\
        );

    \I__5360\ : InMux
    port map (
            O => \N__31379\,
            I => \N__31364\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__31376\,
            I => \N__31360\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__31373\,
            I => \N__31351\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__31370\,
            I => \N__31351\
        );

    \I__5356\ : Span4Mux_v
    port map (
            O => \N__31367\,
            I => \N__31351\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__31364\,
            I => \N__31351\
        );

    \I__5354\ : InMux
    port map (
            O => \N__31363\,
            I => \N__31346\
        );

    \I__5353\ : Span4Mux_h
    port map (
            O => \N__31360\,
            I => \N__31343\
        );

    \I__5352\ : Span4Mux_h
    port map (
            O => \N__31351\,
            I => \N__31340\
        );

    \I__5351\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31337\
        );

    \I__5350\ : InMux
    port map (
            O => \N__31349\,
            I => \N__31334\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__31346\,
            I => \N__31331\
        );

    \I__5348\ : Span4Mux_h
    port map (
            O => \N__31343\,
            I => \N__31326\
        );

    \I__5347\ : Span4Mux_v
    port map (
            O => \N__31340\,
            I => \N__31326\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__31337\,
            I => \sTrigCounterZ0Z_0\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__31334\,
            I => \sTrigCounterZ0Z_0\
        );

    \I__5344\ : Odrv4
    port map (
            O => \N__31331\,
            I => \sTrigCounterZ0Z_0\
        );

    \I__5343\ : Odrv4
    port map (
            O => \N__31326\,
            I => \sTrigCounterZ0Z_0\
        );

    \I__5342\ : IoInMux
    port map (
            O => \N__31317\,
            I => \N__31314\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__31314\,
            I => \N__31311\
        );

    \I__5340\ : Span12Mux_s3_h
    port map (
            O => \N__31311\,
            I => \N__31308\
        );

    \I__5339\ : Span12Mux_h
    port map (
            O => \N__31308\,
            I => \N__31305\
        );

    \I__5338\ : Odrv12
    port map (
            O => \N__31305\,
            I => \RAM_DATA_1Z0Z_13\
        );

    \I__5337\ : CascadeMux
    port map (
            O => \N__31302\,
            I => \N__31294\
        );

    \I__5336\ : InMux
    port map (
            O => \N__31301\,
            I => \N__31290\
        );

    \I__5335\ : InMux
    port map (
            O => \N__31300\,
            I => \N__31287\
        );

    \I__5334\ : InMux
    port map (
            O => \N__31299\,
            I => \N__31284\
        );

    \I__5333\ : InMux
    port map (
            O => \N__31298\,
            I => \N__31281\
        );

    \I__5332\ : InMux
    port map (
            O => \N__31297\,
            I => \N__31273\
        );

    \I__5331\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31273\
        );

    \I__5330\ : InMux
    port map (
            O => \N__31293\,
            I => \N__31273\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__31290\,
            I => \N__31270\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__31287\,
            I => \N__31263\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__31284\,
            I => \N__31263\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__31281\,
            I => \N__31263\
        );

    \I__5325\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31259\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__31273\,
            I => \N__31256\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__31270\,
            I => \N__31253\
        );

    \I__5322\ : Span4Mux_h
    port map (
            O => \N__31263\,
            I => \N__31250\
        );

    \I__5321\ : InMux
    port map (
            O => \N__31262\,
            I => \N__31247\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__31259\,
            I => \N__31242\
        );

    \I__5319\ : Span4Mux_h
    port map (
            O => \N__31256\,
            I => \N__31242\
        );

    \I__5318\ : Span4Mux_h
    port map (
            O => \N__31253\,
            I => \N__31237\
        );

    \I__5317\ : Span4Mux_v
    port map (
            O => \N__31250\,
            I => \N__31237\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__31247\,
            I => \sTrigCounterZ0Z_1\
        );

    \I__5315\ : Odrv4
    port map (
            O => \N__31242\,
            I => \sTrigCounterZ0Z_1\
        );

    \I__5314\ : Odrv4
    port map (
            O => \N__31237\,
            I => \sTrigCounterZ0Z_1\
        );

    \I__5313\ : IoInMux
    port map (
            O => \N__31230\,
            I => \N__31227\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__31227\,
            I => \N__31224\
        );

    \I__5311\ : Span12Mux_s3_h
    port map (
            O => \N__31224\,
            I => \N__31221\
        );

    \I__5310\ : Span12Mux_h
    port map (
            O => \N__31221\,
            I => \N__31218\
        );

    \I__5309\ : Odrv12
    port map (
            O => \N__31218\,
            I => \RAM_DATA_1Z0Z_14\
        );

    \I__5308\ : InMux
    port map (
            O => \N__31215\,
            I => \N__31212\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__31212\,
            I => \N__31209\
        );

    \I__5306\ : Span4Mux_v
    port map (
            O => \N__31209\,
            I => \N__31206\
        );

    \I__5305\ : Sp12to4
    port map (
            O => \N__31206\,
            I => \N__31203\
        );

    \I__5304\ : Span12Mux_h
    port map (
            O => \N__31203\,
            I => \N__31200\
        );

    \I__5303\ : Odrv12
    port map (
            O => \N__31200\,
            I => \ADC2_c\
        );

    \I__5302\ : IoInMux
    port map (
            O => \N__31197\,
            I => \N__31194\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__31194\,
            I => \N__31191\
        );

    \I__5300\ : Span12Mux_s3_v
    port map (
            O => \N__31191\,
            I => \N__31188\
        );

    \I__5299\ : Span12Mux_h
    port map (
            O => \N__31188\,
            I => \N__31185\
        );

    \I__5298\ : Odrv12
    port map (
            O => \N__31185\,
            I => \RAM_DATA_1Z0Z_2\
        );

    \I__5297\ : CEMux
    port map (
            O => \N__31182\,
            I => \N__31178\
        );

    \I__5296\ : CEMux
    port map (
            O => \N__31181\,
            I => \N__31175\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__31178\,
            I => \N_31_i\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__31175\,
            I => \N_31_i\
        );

    \I__5293\ : CEMux
    port map (
            O => \N__31170\,
            I => \N__31167\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__31167\,
            I => \N__31164\
        );

    \I__5291\ : Span12Mux_v
    port map (
            O => \N__31164\,
            I => \N__31161\
        );

    \I__5290\ : Odrv12
    port map (
            O => \N__31161\,
            I => \sAddress_RNIA6242Z0Z_2\
        );

    \I__5289\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31155\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__31155\,
            I => \sDAC_mem_19Z0Z_4\
        );

    \I__5287\ : InMux
    port map (
            O => \N__31152\,
            I => \N__31149\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__31149\,
            I => \sDAC_mem_18Z0Z_4\
        );

    \I__5285\ : InMux
    port map (
            O => \N__31146\,
            I => \N__31143\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__31143\,
            I => \sDAC_mem_19Z0Z_5\
        );

    \I__5283\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31137\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__31137\,
            I => \sDAC_mem_18Z0Z_5\
        );

    \I__5281\ : InMux
    port map (
            O => \N__31134\,
            I => \N__31131\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__31131\,
            I => \sDAC_mem_19Z0Z_6\
        );

    \I__5279\ : InMux
    port map (
            O => \N__31128\,
            I => \N__31125\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__31125\,
            I => \sDAC_mem_18Z0Z_6\
        );

    \I__5277\ : CEMux
    port map (
            O => \N__31122\,
            I => \N__31119\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__31119\,
            I => \N__31116\
        );

    \I__5275\ : Odrv4
    port map (
            O => \N__31116\,
            I => \sDAC_mem_19_1_sqmuxa\
        );

    \I__5274\ : CEMux
    port map (
            O => \N__31113\,
            I => \N__31110\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__31110\,
            I => \sDAC_mem_32_1_sqmuxa\
        );

    \I__5272\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31101\
        );

    \I__5271\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31098\
        );

    \I__5270\ : InMux
    port map (
            O => \N__31105\,
            I => \N__31095\
        );

    \I__5269\ : InMux
    port map (
            O => \N__31104\,
            I => \N__31091\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__31101\,
            I => \N__31087\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__31098\,
            I => \N__31084\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__31095\,
            I => \N__31081\
        );

    \I__5265\ : InMux
    port map (
            O => \N__31094\,
            I => \N__31078\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__31091\,
            I => \N__31075\
        );

    \I__5263\ : InMux
    port map (
            O => \N__31090\,
            I => \N__31067\
        );

    \I__5262\ : Span4Mux_h
    port map (
            O => \N__31087\,
            I => \N__31064\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__31084\,
            I => \N__31059\
        );

    \I__5260\ : Span4Mux_v
    port map (
            O => \N__31081\,
            I => \N__31059\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__31078\,
            I => \N__31056\
        );

    \I__5258\ : Span4Mux_h
    port map (
            O => \N__31075\,
            I => \N__31053\
        );

    \I__5257\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31048\
        );

    \I__5256\ : InMux
    port map (
            O => \N__31073\,
            I => \N__31048\
        );

    \I__5255\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31045\
        );

    \I__5254\ : InMux
    port map (
            O => \N__31071\,
            I => \N__31040\
        );

    \I__5253\ : InMux
    port map (
            O => \N__31070\,
            I => \N__31040\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__31067\,
            I => \N__31037\
        );

    \I__5251\ : Odrv4
    port map (
            O => \N__31064\,
            I => \N_141\
        );

    \I__5250\ : Odrv4
    port map (
            O => \N__31059\,
            I => \N_141\
        );

    \I__5249\ : Odrv4
    port map (
            O => \N__31056\,
            I => \N_141\
        );

    \I__5248\ : Odrv4
    port map (
            O => \N__31053\,
            I => \N_141\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__31048\,
            I => \N_141\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__31045\,
            I => \N_141\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__31040\,
            I => \N_141\
        );

    \I__5244\ : Odrv4
    port map (
            O => \N__31037\,
            I => \N_141\
        );

    \I__5243\ : CEMux
    port map (
            O => \N__31020\,
            I => \N__31017\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__31017\,
            I => \N__31013\
        );

    \I__5241\ : CEMux
    port map (
            O => \N__31016\,
            I => \N__31010\
        );

    \I__5240\ : Span4Mux_h
    port map (
            O => \N__31013\,
            I => \N__31005\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__31010\,
            I => \N__31005\
        );

    \I__5238\ : Span4Mux_h
    port map (
            O => \N__31005\,
            I => \N__31002\
        );

    \I__5237\ : Odrv4
    port map (
            O => \N__31002\,
            I => \sEETrigCounter_1_sqmuxa\
        );

    \I__5236\ : CascadeMux
    port map (
            O => \N__30999\,
            I => \N_1480_cascade_\
        );

    \I__5235\ : InMux
    port map (
            O => \N__30996\,
            I => \N__30993\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__30993\,
            I => \N__30988\
        );

    \I__5233\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30985\
        );

    \I__5232\ : InMux
    port map (
            O => \N__30991\,
            I => \N__30982\
        );

    \I__5231\ : Odrv4
    port map (
            O => \N__30988\,
            I => un1_spointer11_5_0_2
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__30985\,
            I => un1_spointer11_5_0_2
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__30982\,
            I => un1_spointer11_5_0_2
        );

    \I__5228\ : CEMux
    port map (
            O => \N__30975\,
            I => \N__30972\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__30972\,
            I => \N__30969\
        );

    \I__5226\ : Span4Mux_v
    port map (
            O => \N__30969\,
            I => \N__30966\
        );

    \I__5225\ : Odrv4
    port map (
            O => \N__30966\,
            I => \sAddress_RNIA6242_2Z0Z_2\
        );

    \I__5224\ : CascadeMux
    port map (
            O => \N__30963\,
            I => \N_280_cascade_\
        );

    \I__5223\ : CEMux
    port map (
            O => \N__30960\,
            I => \N__30957\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__30957\,
            I => \sDAC_mem_17_1_sqmuxa\
        );

    \I__5221\ : InMux
    port map (
            O => \N__30954\,
            I => \N__30951\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__30951\,
            I => \N__30948\
        );

    \I__5219\ : Span4Mux_v
    port map (
            O => \N__30948\,
            I => \N__30943\
        );

    \I__5218\ : InMux
    port map (
            O => \N__30947\,
            I => \N__30938\
        );

    \I__5217\ : InMux
    port map (
            O => \N__30946\,
            I => \N__30938\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__30943\,
            I => \sAddressZ0Z_6\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__30938\,
            I => \sAddressZ0Z_6\
        );

    \I__5214\ : CascadeMux
    port map (
            O => \N__30933\,
            I => \N__30930\
        );

    \I__5213\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30927\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__30927\,
            I => \N__30923\
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__30926\,
            I => \N__30919\
        );

    \I__5210\ : Span4Mux_h
    port map (
            O => \N__30923\,
            I => \N__30916\
        );

    \I__5209\ : InMux
    port map (
            O => \N__30922\,
            I => \N__30911\
        );

    \I__5208\ : InMux
    port map (
            O => \N__30919\,
            I => \N__30911\
        );

    \I__5207\ : Odrv4
    port map (
            O => \N__30916\,
            I => \sAddressZ0Z_7\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__30911\,
            I => \sAddressZ0Z_7\
        );

    \I__5205\ : InMux
    port map (
            O => \N__30906\,
            I => \N__30903\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__30903\,
            I => \sEEPonPoff_1_sqmuxa_0_a2_1\
        );

    \I__5203\ : CEMux
    port map (
            O => \N__30900\,
            I => \N__30897\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__30897\,
            I => \N__30893\
        );

    \I__5201\ : CEMux
    port map (
            O => \N__30896\,
            I => \N__30890\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__30893\,
            I => \N__30887\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__30890\,
            I => \N__30884\
        );

    \I__5198\ : Span4Mux_h
    port map (
            O => \N__30887\,
            I => \N__30881\
        );

    \I__5197\ : Sp12to4
    port map (
            O => \N__30884\,
            I => \N__30878\
        );

    \I__5196\ : Odrv4
    port map (
            O => \N__30881\,
            I => \sEEPon_1_sqmuxa\
        );

    \I__5195\ : Odrv12
    port map (
            O => \N__30878\,
            I => \sEEPon_1_sqmuxa\
        );

    \I__5194\ : InMux
    port map (
            O => \N__30873\,
            I => \N__30861\
        );

    \I__5193\ : InMux
    port map (
            O => \N__30872\,
            I => \N__30861\
        );

    \I__5192\ : InMux
    port map (
            O => \N__30871\,
            I => \N__30861\
        );

    \I__5191\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30861\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__30861\,
            I => \N_291\
        );

    \I__5189\ : CEMux
    port map (
            O => \N__30858\,
            I => \N__30855\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__30855\,
            I => \N__30852\
        );

    \I__5187\ : Odrv4
    port map (
            O => \N__30852\,
            I => \sDAC_mem_33_1_sqmuxa\
        );

    \I__5186\ : InMux
    port map (
            O => \N__30849\,
            I => \N__30846\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__30846\,
            I => \sDAC_mem_23Z0Z_2\
        );

    \I__5184\ : InMux
    port map (
            O => \N__30843\,
            I => \N__30840\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__30840\,
            I => \sDAC_mem_22Z0Z_2\
        );

    \I__5182\ : InMux
    port map (
            O => \N__30837\,
            I => \N__30834\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__30834\,
            I => \sDAC_mem_23Z0Z_3\
        );

    \I__5180\ : InMux
    port map (
            O => \N__30831\,
            I => \N__30828\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__30828\,
            I => \sDAC_mem_22Z0Z_3\
        );

    \I__5178\ : InMux
    port map (
            O => \N__30825\,
            I => \N__30822\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__30822\,
            I => \sDAC_mem_23Z0Z_4\
        );

    \I__5176\ : InMux
    port map (
            O => \N__30819\,
            I => \N__30816\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__30816\,
            I => \sDAC_mem_22Z0Z_4\
        );

    \I__5174\ : CascadeMux
    port map (
            O => \N__30813\,
            I => \N_291_cascade_\
        );

    \I__5173\ : CEMux
    port map (
            O => \N__30810\,
            I => \N__30807\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__30807\,
            I => \N__30804\
        );

    \I__5171\ : Span4Mux_h
    port map (
            O => \N__30804\,
            I => \N__30801\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__30801\,
            I => \N__30798\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__30798\,
            I => \sEEPonPoff_1_sqmuxa\
        );

    \I__5168\ : InMux
    port map (
            O => \N__30795\,
            I => \N__30791\
        );

    \I__5167\ : InMux
    port map (
            O => \N__30794\,
            I => \N__30788\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__30791\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__30788\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0\
        );

    \I__5164\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30779\
        );

    \I__5163\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30776\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__30779\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__30776\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1\
        );

    \I__5160\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30767\
        );

    \I__5159\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30764\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__30767\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__30764\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2\
        );

    \I__5156\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30755\
        );

    \I__5155\ : InMux
    port map (
            O => \N__30758\,
            I => \N__30752\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__30755\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__30752\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3\
        );

    \I__5152\ : InMux
    port map (
            O => \N__30747\,
            I => \N__30743\
        );

    \I__5151\ : InMux
    port map (
            O => \N__30746\,
            I => \N__30740\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__30743\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__30740\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4\
        );

    \I__5148\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30731\
        );

    \I__5147\ : InMux
    port map (
            O => \N__30734\,
            I => \N__30728\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__30731\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__30728\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5\
        );

    \I__5144\ : InMux
    port map (
            O => \N__30723\,
            I => \N__30719\
        );

    \I__5143\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30716\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__30719\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__30716\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6\
        );

    \I__5140\ : InMux
    port map (
            O => \N__30711\,
            I => \N__30708\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__30708\,
            I => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7\
        );

    \I__5138\ : ClkMux
    port map (
            O => \N__30705\,
            I => \N__30678\
        );

    \I__5137\ : ClkMux
    port map (
            O => \N__30704\,
            I => \N__30678\
        );

    \I__5136\ : ClkMux
    port map (
            O => \N__30703\,
            I => \N__30678\
        );

    \I__5135\ : ClkMux
    port map (
            O => \N__30702\,
            I => \N__30678\
        );

    \I__5134\ : ClkMux
    port map (
            O => \N__30701\,
            I => \N__30678\
        );

    \I__5133\ : ClkMux
    port map (
            O => \N__30700\,
            I => \N__30678\
        );

    \I__5132\ : ClkMux
    port map (
            O => \N__30699\,
            I => \N__30678\
        );

    \I__5131\ : ClkMux
    port map (
            O => \N__30698\,
            I => \N__30678\
        );

    \I__5130\ : ClkMux
    port map (
            O => \N__30697\,
            I => \N__30678\
        );

    \I__5129\ : GlobalMux
    port map (
            O => \N__30678\,
            I => \N__30675\
        );

    \I__5128\ : gio2CtrlBuf
    port map (
            O => \N__30675\,
            I => spi_sclk_g
        );

    \I__5127\ : CEMux
    port map (
            O => \N__30672\,
            I => \N__30668\
        );

    \I__5126\ : CEMux
    port map (
            O => \N__30671\,
            I => \N__30665\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__30668\,
            I => \N__30661\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__30665\,
            I => \N__30658\
        );

    \I__5123\ : CEMux
    port map (
            O => \N__30664\,
            I => \N__30655\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__30661\,
            I => \N__30652\
        );

    \I__5121\ : Span4Mux_h
    port map (
            O => \N__30658\,
            I => \N__30649\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__30655\,
            I => \N__30646\
        );

    \I__5119\ : Odrv4
    port map (
            O => \N__30652\,
            I => \spi_slave_inst.spi_cs_iZ0\
        );

    \I__5118\ : Odrv4
    port map (
            O => \N__30649\,
            I => \spi_slave_inst.spi_cs_iZ0\
        );

    \I__5117\ : Odrv4
    port map (
            O => \N__30646\,
            I => \spi_slave_inst.spi_cs_iZ0\
        );

    \I__5116\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30636\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__30636\,
            I => \N__30633\
        );

    \I__5114\ : Span12Mux_s11_v
    port map (
            O => \N__30633\,
            I => \N__30630\
        );

    \I__5113\ : Span12Mux_h
    port map (
            O => \N__30630\,
            I => \N__30627\
        );

    \I__5112\ : Odrv12
    port map (
            O => \N__30627\,
            I => \ADC8_c\
        );

    \I__5111\ : IoInMux
    port map (
            O => \N__30624\,
            I => \N__30621\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__30621\,
            I => \N__30618\
        );

    \I__5109\ : IoSpan4Mux
    port map (
            O => \N__30618\,
            I => \N__30615\
        );

    \I__5108\ : Span4Mux_s3_h
    port map (
            O => \N__30615\,
            I => \N__30612\
        );

    \I__5107\ : Sp12to4
    port map (
            O => \N__30612\,
            I => \N__30609\
        );

    \I__5106\ : Span12Mux_h
    port map (
            O => \N__30609\,
            I => \N__30606\
        );

    \I__5105\ : Span12Mux_v
    port map (
            O => \N__30606\,
            I => \N__30603\
        );

    \I__5104\ : Odrv12
    port map (
            O => \N__30603\,
            I => \RAM_DATA_1Z0Z_9\
        );

    \I__5103\ : IoInMux
    port map (
            O => \N__30600\,
            I => \N__30597\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__30597\,
            I => \N__30594\
        );

    \I__5101\ : Span4Mux_s2_h
    port map (
            O => \N__30594\,
            I => \N__30591\
        );

    \I__5100\ : Sp12to4
    port map (
            O => \N__30591\,
            I => \N__30588\
        );

    \I__5099\ : Span12Mux_v
    port map (
            O => \N__30588\,
            I => \N__30585\
        );

    \I__5098\ : Span12Mux_h
    port map (
            O => \N__30585\,
            I => \N__30582\
        );

    \I__5097\ : Odrv12
    port map (
            O => \N__30582\,
            I => \RAM_DATA_1Z0Z_15\
        );

    \I__5096\ : IoInMux
    port map (
            O => \N__30579\,
            I => \N__30576\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__30576\,
            I => \N__30573\
        );

    \I__5094\ : IoSpan4Mux
    port map (
            O => \N__30573\,
            I => \N__30570\
        );

    \I__5093\ : Span4Mux_s1_v
    port map (
            O => \N__30570\,
            I => \N__30567\
        );

    \I__5092\ : Sp12to4
    port map (
            O => \N__30567\,
            I => \N__30564\
        );

    \I__5091\ : Span12Mux_h
    port map (
            O => \N__30564\,
            I => \N__30561\
        );

    \I__5090\ : Odrv12
    port map (
            O => \N__30561\,
            I => \RAM_DATA_1Z0Z_7\
        );

    \I__5089\ : IoInMux
    port map (
            O => \N__30558\,
            I => \N__30555\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__30555\,
            I => \N__30552\
        );

    \I__5087\ : Span4Mux_s2_v
    port map (
            O => \N__30552\,
            I => \N__30549\
        );

    \I__5086\ : Span4Mux_h
    port map (
            O => \N__30549\,
            I => \N__30546\
        );

    \I__5085\ : Span4Mux_h
    port map (
            O => \N__30546\,
            I => \N__30543\
        );

    \I__5084\ : Span4Mux_h
    port map (
            O => \N__30543\,
            I => \N__30540\
        );

    \I__5083\ : Span4Mux_v
    port map (
            O => \N__30540\,
            I => \N__30536\
        );

    \I__5082\ : InMux
    port map (
            O => \N__30539\,
            I => \N__30533\
        );

    \I__5081\ : Odrv4
    port map (
            O => \N__30536\,
            I => \RAM_DATA_cl_1Z0Z_15\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__30533\,
            I => \RAM_DATA_cl_1Z0Z_15\
        );

    \I__5079\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30525\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__30525\,
            I => \N_100\
        );

    \I__5077\ : IoInMux
    port map (
            O => \N__30522\,
            I => \N__30519\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__30519\,
            I => \N__30516\
        );

    \I__5075\ : IoSpan4Mux
    port map (
            O => \N__30516\,
            I => \N__30513\
        );

    \I__5074\ : IoSpan4Mux
    port map (
            O => \N__30513\,
            I => \N__30510\
        );

    \I__5073\ : Span4Mux_s3_h
    port map (
            O => \N__30510\,
            I => \N__30507\
        );

    \I__5072\ : Sp12to4
    port map (
            O => \N__30507\,
            I => \N__30504\
        );

    \I__5071\ : Span12Mux_h
    port map (
            O => \N__30504\,
            I => \N__30500\
        );

    \I__5070\ : InMux
    port map (
            O => \N__30503\,
            I => \N__30497\
        );

    \I__5069\ : Odrv12
    port map (
            O => \N__30500\,
            I => \RAM_DATA_cl_13Z0Z_15\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__30497\,
            I => \RAM_DATA_cl_13Z0Z_15\
        );

    \I__5067\ : InMux
    port map (
            O => \N__30492\,
            I => \N__30489\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__30489\,
            I => \N_97\
        );

    \I__5065\ : IoInMux
    port map (
            O => \N__30486\,
            I => \N__30483\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__30483\,
            I => \N__30480\
        );

    \I__5063\ : IoSpan4Mux
    port map (
            O => \N__30480\,
            I => \N__30477\
        );

    \I__5062\ : IoSpan4Mux
    port map (
            O => \N__30477\,
            I => \N__30474\
        );

    \I__5061\ : Sp12to4
    port map (
            O => \N__30474\,
            I => \N__30471\
        );

    \I__5060\ : Span12Mux_s7_h
    port map (
            O => \N__30471\,
            I => \N__30467\
        );

    \I__5059\ : InMux
    port map (
            O => \N__30470\,
            I => \N__30464\
        );

    \I__5058\ : Odrv12
    port map (
            O => \N__30467\,
            I => \RAM_DATA_cl_2Z0Z_15\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__30464\,
            I => \RAM_DATA_cl_2Z0Z_15\
        );

    \I__5056\ : InMux
    port map (
            O => \N__30459\,
            I => \N__30456\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__30456\,
            I => \N_101\
        );

    \I__5054\ : InMux
    port map (
            O => \N__30453\,
            I => \N__30450\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__30450\,
            I => \N_103\
        );

    \I__5052\ : IoInMux
    port map (
            O => \N__30447\,
            I => \N__30444\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__30444\,
            I => \N__30441\
        );

    \I__5050\ : Span4Mux_s3_v
    port map (
            O => \N__30441\,
            I => \N__30438\
        );

    \I__5049\ : Span4Mux_h
    port map (
            O => \N__30438\,
            I => \N__30435\
        );

    \I__5048\ : Span4Mux_h
    port map (
            O => \N__30435\,
            I => \N__30432\
        );

    \I__5047\ : Span4Mux_h
    port map (
            O => \N__30432\,
            I => \N__30428\
        );

    \I__5046\ : InMux
    port map (
            O => \N__30431\,
            I => \N__30425\
        );

    \I__5045\ : Odrv4
    port map (
            O => \N__30428\,
            I => \RAM_DATA_cl_3Z0Z_15\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__30425\,
            I => \RAM_DATA_cl_3Z0Z_15\
        );

    \I__5043\ : InMux
    port map (
            O => \N__30420\,
            I => \N__30417\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__30417\,
            I => \N__30414\
        );

    \I__5041\ : Span12Mux_v
    port map (
            O => \N__30414\,
            I => \N__30411\
        );

    \I__5040\ : Span12Mux_h
    port map (
            O => \N__30411\,
            I => \N__30408\
        );

    \I__5039\ : Odrv12
    port map (
            O => \N__30408\,
            I => spi_mosi_ft_c
        );

    \I__5038\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30402\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__30402\,
            I => \N__30399\
        );

    \I__5036\ : Span4Mux_v
    port map (
            O => \N__30399\,
            I => \N__30396\
        );

    \I__5035\ : Sp12to4
    port map (
            O => \N__30396\,
            I => \N__30393\
        );

    \I__5034\ : Span12Mux_h
    port map (
            O => \N__30393\,
            I => \N__30389\
        );

    \I__5033\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30386\
        );

    \I__5032\ : Odrv12
    port map (
            O => \N__30389\,
            I => \sRAM_pointer_readZ0Z_11\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__30386\,
            I => \sRAM_pointer_readZ0Z_11\
        );

    \I__5030\ : IoInMux
    port map (
            O => \N__30381\,
            I => \N__30378\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__30378\,
            I => \N__30375\
        );

    \I__5028\ : IoSpan4Mux
    port map (
            O => \N__30375\,
            I => \N__30372\
        );

    \I__5027\ : Span4Mux_s1_h
    port map (
            O => \N__30372\,
            I => \N__30369\
        );

    \I__5026\ : Span4Mux_v
    port map (
            O => \N__30369\,
            I => \N__30366\
        );

    \I__5025\ : Sp12to4
    port map (
            O => \N__30366\,
            I => \N__30363\
        );

    \I__5024\ : Span12Mux_v
    port map (
            O => \N__30363\,
            I => \N__30360\
        );

    \I__5023\ : Span12Mux_h
    port map (
            O => \N__30360\,
            I => \N__30357\
        );

    \I__5022\ : Odrv12
    port map (
            O => \N__30357\,
            I => \RAM_ADD_c_11\
        );

    \I__5021\ : CascadeMux
    port map (
            O => \N__30354\,
            I => \N__30351\
        );

    \I__5020\ : InMux
    port map (
            O => \N__30351\,
            I => \N__30348\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__30348\,
            I => \N__30345\
        );

    \I__5018\ : Span4Mux_v
    port map (
            O => \N__30345\,
            I => \N__30342\
        );

    \I__5017\ : Span4Mux_v
    port map (
            O => \N__30342\,
            I => \N__30339\
        );

    \I__5016\ : Sp12to4
    port map (
            O => \N__30339\,
            I => \N__30335\
        );

    \I__5015\ : InMux
    port map (
            O => \N__30338\,
            I => \N__30332\
        );

    \I__5014\ : Odrv12
    port map (
            O => \N__30335\,
            I => \sRAM_pointer_readZ0Z_12\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__30332\,
            I => \sRAM_pointer_readZ0Z_12\
        );

    \I__5012\ : IoInMux
    port map (
            O => \N__30327\,
            I => \N__30324\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__30324\,
            I => \N__30321\
        );

    \I__5010\ : Span12Mux_s4_h
    port map (
            O => \N__30321\,
            I => \N__30318\
        );

    \I__5009\ : Span12Mux_v
    port map (
            O => \N__30318\,
            I => \N__30315\
        );

    \I__5008\ : Span12Mux_h
    port map (
            O => \N__30315\,
            I => \N__30312\
        );

    \I__5007\ : Odrv12
    port map (
            O => \N__30312\,
            I => \RAM_ADD_c_12\
        );

    \I__5006\ : InMux
    port map (
            O => \N__30309\,
            I => \N__30306\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__30306\,
            I => \N__30303\
        );

    \I__5004\ : Span12Mux_h
    port map (
            O => \N__30303\,
            I => \N__30299\
        );

    \I__5003\ : InMux
    port map (
            O => \N__30302\,
            I => \N__30296\
        );

    \I__5002\ : Odrv12
    port map (
            O => \N__30299\,
            I => \sRAM_pointer_readZ0Z_13\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__30296\,
            I => \sRAM_pointer_readZ0Z_13\
        );

    \I__5000\ : IoInMux
    port map (
            O => \N__30291\,
            I => \N__30288\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__30288\,
            I => \N__30285\
        );

    \I__4998\ : Span4Mux_s3_h
    port map (
            O => \N__30285\,
            I => \N__30282\
        );

    \I__4997\ : Sp12to4
    port map (
            O => \N__30282\,
            I => \N__30279\
        );

    \I__4996\ : Span12Mux_s10_v
    port map (
            O => \N__30279\,
            I => \N__30276\
        );

    \I__4995\ : Span12Mux_h
    port map (
            O => \N__30276\,
            I => \N__30273\
        );

    \I__4994\ : Span12Mux_v
    port map (
            O => \N__30273\,
            I => \N__30270\
        );

    \I__4993\ : Odrv12
    port map (
            O => \N__30270\,
            I => \RAM_ADD_c_13\
        );

    \I__4992\ : CEMux
    port map (
            O => \N__30267\,
            I => \N__30264\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__30264\,
            I => \N__30259\
        );

    \I__4990\ : CEMux
    port map (
            O => \N__30263\,
            I => \N__30256\
        );

    \I__4989\ : CEMux
    port map (
            O => \N__30262\,
            I => \N__30253\
        );

    \I__4988\ : Span4Mux_v
    port map (
            O => \N__30259\,
            I => \N__30248\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__30256\,
            I => \N__30248\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__30253\,
            I => \N__30243\
        );

    \I__4985\ : Span4Mux_v
    port map (
            O => \N__30248\,
            I => \N__30243\
        );

    \I__4984\ : Odrv4
    port map (
            O => \N__30243\,
            I => \N_67_i\
        );

    \I__4983\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30237\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__30237\,
            I => \N__30234\
        );

    \I__4981\ : Span4Mux_v
    port map (
            O => \N__30234\,
            I => \N__30231\
        );

    \I__4980\ : Sp12to4
    port map (
            O => \N__30231\,
            I => \N__30228\
        );

    \I__4979\ : Span12Mux_h
    port map (
            O => \N__30228\,
            I => \N__30225\
        );

    \I__4978\ : Odrv12
    port map (
            O => \N__30225\,
            I => \ADC3_c\
        );

    \I__4977\ : IoInMux
    port map (
            O => \N__30222\,
            I => \N__30219\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__30219\,
            I => \N__30216\
        );

    \I__4975\ : Span4Mux_s0_v
    port map (
            O => \N__30216\,
            I => \N__30213\
        );

    \I__4974\ : Sp12to4
    port map (
            O => \N__30213\,
            I => \N__30210\
        );

    \I__4973\ : Span12Mux_h
    port map (
            O => \N__30210\,
            I => \N__30207\
        );

    \I__4972\ : Odrv12
    port map (
            O => \N__30207\,
            I => \RAM_DATA_1Z0Z_3\
        );

    \I__4971\ : InMux
    port map (
            O => \N__30204\,
            I => \N__30201\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__30201\,
            I => \N__30198\
        );

    \I__4969\ : Span4Mux_v
    port map (
            O => \N__30198\,
            I => \N__30195\
        );

    \I__4968\ : Sp12to4
    port map (
            O => \N__30195\,
            I => \N__30192\
        );

    \I__4967\ : Span12Mux_h
    port map (
            O => \N__30192\,
            I => \N__30189\
        );

    \I__4966\ : Odrv12
    port map (
            O => \N__30189\,
            I => \ADC0_c\
        );

    \I__4965\ : IoInMux
    port map (
            O => \N__30186\,
            I => \N__30183\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__30183\,
            I => \N__30180\
        );

    \I__4963\ : Span4Mux_s3_v
    port map (
            O => \N__30180\,
            I => \N__30177\
        );

    \I__4962\ : Span4Mux_h
    port map (
            O => \N__30177\,
            I => \N__30174\
        );

    \I__4961\ : Sp12to4
    port map (
            O => \N__30174\,
            I => \N__30171\
        );

    \I__4960\ : Span12Mux_s8_v
    port map (
            O => \N__30171\,
            I => \N__30168\
        );

    \I__4959\ : Odrv12
    port map (
            O => \N__30168\,
            I => \RAM_DATA_1Z0Z_0\
        );

    \I__4958\ : InMux
    port map (
            O => \N__30165\,
            I => \N__30162\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__30162\,
            I => \N__30159\
        );

    \I__4956\ : Span4Mux_v
    port map (
            O => \N__30159\,
            I => \N__30156\
        );

    \I__4955\ : Sp12to4
    port map (
            O => \N__30156\,
            I => \N__30153\
        );

    \I__4954\ : Span12Mux_h
    port map (
            O => \N__30153\,
            I => \N__30150\
        );

    \I__4953\ : Odrv12
    port map (
            O => \N__30150\,
            I => \ADC5_c\
        );

    \I__4952\ : IoInMux
    port map (
            O => \N__30147\,
            I => \N__30144\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__30144\,
            I => \N__30141\
        );

    \I__4950\ : IoSpan4Mux
    port map (
            O => \N__30141\,
            I => \N__30138\
        );

    \I__4949\ : Span4Mux_s2_v
    port map (
            O => \N__30138\,
            I => \N__30135\
        );

    \I__4948\ : Sp12to4
    port map (
            O => \N__30135\,
            I => \N__30132\
        );

    \I__4947\ : Span12Mux_s10_v
    port map (
            O => \N__30132\,
            I => \N__30129\
        );

    \I__4946\ : Span12Mux_h
    port map (
            O => \N__30129\,
            I => \N__30126\
        );

    \I__4945\ : Odrv12
    port map (
            O => \N__30126\,
            I => \RAM_DATA_1Z0Z_5\
        );

    \I__4944\ : InMux
    port map (
            O => \N__30123\,
            I => \N__30120\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__30120\,
            I => \N__30117\
        );

    \I__4942\ : Span4Mux_v
    port map (
            O => \N__30117\,
            I => \N__30114\
        );

    \I__4941\ : Sp12to4
    port map (
            O => \N__30114\,
            I => \N__30111\
        );

    \I__4940\ : Span12Mux_h
    port map (
            O => \N__30111\,
            I => \N__30108\
        );

    \I__4939\ : Odrv12
    port map (
            O => \N__30108\,
            I => \ADC1_c\
        );

    \I__4938\ : IoInMux
    port map (
            O => \N__30105\,
            I => \N__30102\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__30102\,
            I => \N__30099\
        );

    \I__4936\ : Span12Mux_s9_v
    port map (
            O => \N__30099\,
            I => \N__30096\
        );

    \I__4935\ : Span12Mux_h
    port map (
            O => \N__30096\,
            I => \N__30093\
        );

    \I__4934\ : Odrv12
    port map (
            O => \N__30093\,
            I => \RAM_DATA_1Z0Z_1\
        );

    \I__4933\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30087\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__30087\,
            I => \N__30084\
        );

    \I__4931\ : Span12Mux_s9_v
    port map (
            O => \N__30084\,
            I => \N__30081\
        );

    \I__4930\ : Span12Mux_h
    port map (
            O => \N__30081\,
            I => \N__30078\
        );

    \I__4929\ : Odrv12
    port map (
            O => \N__30078\,
            I => \ADC7_c\
        );

    \I__4928\ : IoInMux
    port map (
            O => \N__30075\,
            I => \N__30072\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__30072\,
            I => \N__30069\
        );

    \I__4926\ : Span4Mux_s0_h
    port map (
            O => \N__30069\,
            I => \N__30066\
        );

    \I__4925\ : Span4Mux_v
    port map (
            O => \N__30066\,
            I => \N__30063\
        );

    \I__4924\ : Sp12to4
    port map (
            O => \N__30063\,
            I => \N__30060\
        );

    \I__4923\ : Span12Mux_v
    port map (
            O => \N__30060\,
            I => \N__30057\
        );

    \I__4922\ : Span12Mux_h
    port map (
            O => \N__30057\,
            I => \N__30054\
        );

    \I__4921\ : Odrv12
    port map (
            O => \N__30054\,
            I => \RAM_DATA_1Z0Z_8\
        );

    \I__4920\ : InMux
    port map (
            O => \N__30051\,
            I => \N__30048\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__30048\,
            I => \N__30045\
        );

    \I__4918\ : Span4Mux_h
    port map (
            O => \N__30045\,
            I => \N__30042\
        );

    \I__4917\ : Sp12to4
    port map (
            O => \N__30042\,
            I => \N__30039\
        );

    \I__4916\ : Span12Mux_v
    port map (
            O => \N__30039\,
            I => \N__30036\
        );

    \I__4915\ : Span12Mux_h
    port map (
            O => \N__30036\,
            I => \N__30033\
        );

    \I__4914\ : Odrv12
    port map (
            O => \N__30033\,
            I => \RAM_DATA_in_11\
        );

    \I__4913\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30027\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__30027\,
            I => \N__30024\
        );

    \I__4911\ : Span4Mux_v
    port map (
            O => \N__30024\,
            I => \N__30021\
        );

    \I__4910\ : Span4Mux_v
    port map (
            O => \N__30021\,
            I => \N__30018\
        );

    \I__4909\ : Sp12to4
    port map (
            O => \N__30018\,
            I => \N__30015\
        );

    \I__4908\ : Span12Mux_h
    port map (
            O => \N__30015\,
            I => \N__30012\
        );

    \I__4907\ : Odrv12
    port map (
            O => \N__30012\,
            I => \RAM_DATA_in_3\
        );

    \I__4906\ : InMux
    port map (
            O => \N__30009\,
            I => \N__30006\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__30006\,
            I => \N__30003\
        );

    \I__4904\ : Span4Mux_h
    port map (
            O => \N__30003\,
            I => \N__30000\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__30000\,
            I => \spi_data_misoZ0Z_3\
        );

    \I__4902\ : InMux
    port map (
            O => \N__29997\,
            I => \N__29994\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__29994\,
            I => \N__29991\
        );

    \I__4900\ : Span4Mux_v
    port map (
            O => \N__29991\,
            I => \N__29988\
        );

    \I__4899\ : Sp12to4
    port map (
            O => \N__29988\,
            I => \N__29985\
        );

    \I__4898\ : Span12Mux_v
    port map (
            O => \N__29985\,
            I => \N__29982\
        );

    \I__4897\ : Span12Mux_h
    port map (
            O => \N__29982\,
            I => \N__29979\
        );

    \I__4896\ : Odrv12
    port map (
            O => \N__29979\,
            I => \RAM_DATA_in_12\
        );

    \I__4895\ : CascadeMux
    port map (
            O => \N__29976\,
            I => \N__29973\
        );

    \I__4894\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29970\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__29970\,
            I => \N__29967\
        );

    \I__4892\ : Span4Mux_v
    port map (
            O => \N__29967\,
            I => \N__29964\
        );

    \I__4891\ : Span4Mux_v
    port map (
            O => \N__29964\,
            I => \N__29961\
        );

    \I__4890\ : Sp12to4
    port map (
            O => \N__29961\,
            I => \N__29958\
        );

    \I__4889\ : Span12Mux_h
    port map (
            O => \N__29958\,
            I => \N__29955\
        );

    \I__4888\ : Odrv12
    port map (
            O => \N__29955\,
            I => \RAM_DATA_in_4\
        );

    \I__4887\ : InMux
    port map (
            O => \N__29952\,
            I => \N__29949\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__29949\,
            I => \N__29946\
        );

    \I__4885\ : Span4Mux_v
    port map (
            O => \N__29946\,
            I => \N__29943\
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__29943\,
            I => \spi_data_misoZ0Z_4\
        );

    \I__4883\ : CEMux
    port map (
            O => \N__29940\,
            I => \N__29934\
        );

    \I__4882\ : InMux
    port map (
            O => \N__29939\,
            I => \N__29926\
        );

    \I__4881\ : InMux
    port map (
            O => \N__29938\,
            I => \N__29926\
        );

    \I__4880\ : InMux
    port map (
            O => \N__29937\,
            I => \N__29926\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__29934\,
            I => \N__29917\
        );

    \I__4878\ : InMux
    port map (
            O => \N__29933\,
            I => \N__29914\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__29926\,
            I => \N__29911\
        );

    \I__4876\ : InMux
    port map (
            O => \N__29925\,
            I => \N__29898\
        );

    \I__4875\ : InMux
    port map (
            O => \N__29924\,
            I => \N__29898\
        );

    \I__4874\ : InMux
    port map (
            O => \N__29923\,
            I => \N__29898\
        );

    \I__4873\ : InMux
    port map (
            O => \N__29922\,
            I => \N__29898\
        );

    \I__4872\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29898\
        );

    \I__4871\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29898\
        );

    \I__4870\ : Odrv4
    port map (
            O => \N__29917\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__29914\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__4868\ : Odrv4
    port map (
            O => \N__29911\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__29898\,
            I => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\
        );

    \I__4866\ : InMux
    port map (
            O => \N__29889\,
            I => \N__29886\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__29886\,
            I => \N__29883\
        );

    \I__4864\ : Span4Mux_v
    port map (
            O => \N__29883\,
            I => \N__29880\
        );

    \I__4863\ : Sp12to4
    port map (
            O => \N__29880\,
            I => \N__29877\
        );

    \I__4862\ : Span12Mux_h
    port map (
            O => \N__29877\,
            I => \N__29874\
        );

    \I__4861\ : Odrv12
    port map (
            O => \N__29874\,
            I => \RAM_DATA_in_5\
        );

    \I__4860\ : CascadeMux
    port map (
            O => \N__29871\,
            I => \N__29865\
        );

    \I__4859\ : CascadeMux
    port map (
            O => \N__29870\,
            I => \N__29861\
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__29869\,
            I => \N__29857\
        );

    \I__4857\ : CascadeMux
    port map (
            O => \N__29868\,
            I => \N__29853\
        );

    \I__4856\ : InMux
    port map (
            O => \N__29865\,
            I => \N__29838\
        );

    \I__4855\ : InMux
    port map (
            O => \N__29864\,
            I => \N__29838\
        );

    \I__4854\ : InMux
    port map (
            O => \N__29861\,
            I => \N__29838\
        );

    \I__4853\ : InMux
    port map (
            O => \N__29860\,
            I => \N__29838\
        );

    \I__4852\ : InMux
    port map (
            O => \N__29857\,
            I => \N__29838\
        );

    \I__4851\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29838\
        );

    \I__4850\ : InMux
    port map (
            O => \N__29853\,
            I => \N__29833\
        );

    \I__4849\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29833\
        );

    \I__4848\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29830\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__29838\,
            I => \N_75\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__29833\,
            I => \N_75\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__29830\,
            I => \N_75\
        );

    \I__4844\ : InMux
    port map (
            O => \N__29823\,
            I => \N__29820\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__29820\,
            I => \N__29817\
        );

    \I__4842\ : Span4Mux_v
    port map (
            O => \N__29817\,
            I => \N__29814\
        );

    \I__4841\ : Span4Mux_h
    port map (
            O => \N__29814\,
            I => \N__29811\
        );

    \I__4840\ : Span4Mux_h
    port map (
            O => \N__29811\,
            I => \N__29808\
        );

    \I__4839\ : Span4Mux_h
    port map (
            O => \N__29808\,
            I => \N__29805\
        );

    \I__4838\ : IoSpan4Mux
    port map (
            O => \N__29805\,
            I => \N__29802\
        );

    \I__4837\ : Odrv4
    port map (
            O => \N__29802\,
            I => \RAM_DATA_in_13\
        );

    \I__4836\ : InMux
    port map (
            O => \N__29799\,
            I => \N__29796\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__29796\,
            I => \N__29793\
        );

    \I__4834\ : Span4Mux_v
    port map (
            O => \N__29793\,
            I => \N__29790\
        );

    \I__4833\ : Odrv4
    port map (
            O => \N__29790\,
            I => \spi_data_misoZ0Z_5\
        );

    \I__4832\ : CEMux
    port map (
            O => \N__29787\,
            I => \N__29784\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__29784\,
            I => \N__29781\
        );

    \I__4830\ : Span4Mux_v
    port map (
            O => \N__29781\,
            I => \N__29777\
        );

    \I__4829\ : CEMux
    port map (
            O => \N__29780\,
            I => \N__29774\
        );

    \I__4828\ : Span4Mux_h
    port map (
            O => \N__29777\,
            I => \N__29771\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__29774\,
            I => \N__29768\
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__29771\,
            I => \N_6\
        );

    \I__4825\ : Odrv12
    port map (
            O => \N__29768\,
            I => \N_6\
        );

    \I__4824\ : InMux
    port map (
            O => \N__29763\,
            I => \N__29760\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__29760\,
            I => \N__29757\
        );

    \I__4822\ : Span4Mux_h
    port map (
            O => \N__29757\,
            I => \N__29754\
        );

    \I__4821\ : Sp12to4
    port map (
            O => \N__29754\,
            I => \N__29751\
        );

    \I__4820\ : Span12Mux_v
    port map (
            O => \N__29751\,
            I => \N__29747\
        );

    \I__4819\ : InMux
    port map (
            O => \N__29750\,
            I => \N__29744\
        );

    \I__4818\ : Odrv12
    port map (
            O => \N__29747\,
            I => \sRAM_pointer_readZ0Z_0\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__29744\,
            I => \sRAM_pointer_readZ0Z_0\
        );

    \I__4816\ : IoInMux
    port map (
            O => \N__29739\,
            I => \N__29736\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__29736\,
            I => \N__29733\
        );

    \I__4814\ : Span4Mux_s1_v
    port map (
            O => \N__29733\,
            I => \N__29730\
        );

    \I__4813\ : Span4Mux_v
    port map (
            O => \N__29730\,
            I => \N__29727\
        );

    \I__4812\ : Span4Mux_h
    port map (
            O => \N__29727\,
            I => \N__29724\
        );

    \I__4811\ : Span4Mux_v
    port map (
            O => \N__29724\,
            I => \N__29721\
        );

    \I__4810\ : Odrv4
    port map (
            O => \N__29721\,
            I => \RAM_ADD_c_0\
        );

    \I__4809\ : InMux
    port map (
            O => \N__29718\,
            I => \N__29715\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__29715\,
            I => \N__29712\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__29712\,
            I => \N__29709\
        );

    \I__4806\ : Span4Mux_v
    port map (
            O => \N__29709\,
            I => \N__29706\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__29706\,
            I => \reset_rpi_ibuf_RNI7JCVZ0\
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__29703\,
            I => \N__29700\
        );

    \I__4803\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29694\
        );

    \I__4802\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29694\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__29694\,
            I => \N__29691\
        );

    \I__4800\ : Odrv4
    port map (
            O => \N__29691\,
            I => \sRAM_ADD_0_sqmuxa_i_0\
        );

    \I__4799\ : InMux
    port map (
            O => \N__29688\,
            I => \N__29685\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__29685\,
            I => \N__29682\
        );

    \I__4797\ : Span4Mux_v
    port map (
            O => \N__29682\,
            I => \N__29679\
        );

    \I__4796\ : Sp12to4
    port map (
            O => \N__29679\,
            I => \N__29676\
        );

    \I__4795\ : Span12Mux_h
    port map (
            O => \N__29676\,
            I => \N__29672\
        );

    \I__4794\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29669\
        );

    \I__4793\ : Odrv12
    port map (
            O => \N__29672\,
            I => \sRAM_pointer_readZ0Z_1\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__29669\,
            I => \sRAM_pointer_readZ0Z_1\
        );

    \I__4791\ : IoInMux
    port map (
            O => \N__29664\,
            I => \N__29661\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__29661\,
            I => \N__29658\
        );

    \I__4789\ : Span4Mux_s3_v
    port map (
            O => \N__29658\,
            I => \N__29655\
        );

    \I__4788\ : Span4Mux_h
    port map (
            O => \N__29655\,
            I => \N__29652\
        );

    \I__4787\ : Sp12to4
    port map (
            O => \N__29652\,
            I => \N__29649\
        );

    \I__4786\ : Odrv12
    port map (
            O => \N__29649\,
            I => \RAM_ADD_c_1\
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__29646\,
            I => \N__29643\
        );

    \I__4784\ : InMux
    port map (
            O => \N__29643\,
            I => \N__29640\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__29640\,
            I => \N__29637\
        );

    \I__4782\ : Span4Mux_h
    port map (
            O => \N__29637\,
            I => \N__29634\
        );

    \I__4781\ : Span4Mux_h
    port map (
            O => \N__29634\,
            I => \N__29631\
        );

    \I__4780\ : Span4Mux_h
    port map (
            O => \N__29631\,
            I => \N__29627\
        );

    \I__4779\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29624\
        );

    \I__4778\ : Span4Mux_v
    port map (
            O => \N__29627\,
            I => \N__29621\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__29624\,
            I => \sRAM_pointer_readZ0Z_10\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__29621\,
            I => \sRAM_pointer_readZ0Z_10\
        );

    \I__4775\ : IoInMux
    port map (
            O => \N__29616\,
            I => \N__29613\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__29613\,
            I => \N__29610\
        );

    \I__4773\ : IoSpan4Mux
    port map (
            O => \N__29610\,
            I => \N__29607\
        );

    \I__4772\ : Span4Mux_s0_h
    port map (
            O => \N__29607\,
            I => \N__29604\
        );

    \I__4771\ : Span4Mux_v
    port map (
            O => \N__29604\,
            I => \N__29601\
        );

    \I__4770\ : Sp12to4
    port map (
            O => \N__29601\,
            I => \N__29598\
        );

    \I__4769\ : Span12Mux_v
    port map (
            O => \N__29598\,
            I => \N__29595\
        );

    \I__4768\ : Span12Mux_h
    port map (
            O => \N__29595\,
            I => \N__29592\
        );

    \I__4767\ : Odrv12
    port map (
            O => \N__29592\,
            I => \RAM_ADD_c_10\
        );

    \I__4766\ : InMux
    port map (
            O => \N__29589\,
            I => \sCounterADC_cry_1\
        );

    \I__4765\ : InMux
    port map (
            O => \N__29586\,
            I => \sCounterADC_cry_2\
        );

    \I__4764\ : InMux
    port map (
            O => \N__29583\,
            I => \sCounterADC_cry_3\
        );

    \I__4763\ : InMux
    port map (
            O => \N__29580\,
            I => \sCounterADC_cry_4\
        );

    \I__4762\ : InMux
    port map (
            O => \N__29577\,
            I => \sCounterADC_cry_5\
        );

    \I__4761\ : InMux
    port map (
            O => \N__29574\,
            I => \sCounterADC_cry_6\
        );

    \I__4760\ : InMux
    port map (
            O => \N__29571\,
            I => \N__29568\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__29568\,
            I => \N__29565\
        );

    \I__4758\ : Span4Mux_h
    port map (
            O => \N__29565\,
            I => \N__29562\
        );

    \I__4757\ : Span4Mux_v
    port map (
            O => \N__29562\,
            I => \N__29559\
        );

    \I__4756\ : Sp12to4
    port map (
            O => \N__29559\,
            I => \N__29556\
        );

    \I__4755\ : Span12Mux_v
    port map (
            O => \N__29556\,
            I => \N__29553\
        );

    \I__4754\ : Span12Mux_h
    port map (
            O => \N__29553\,
            I => \N__29550\
        );

    \I__4753\ : Odrv12
    port map (
            O => \N__29550\,
            I => \RAM_DATA_in_8\
        );

    \I__4752\ : CascadeMux
    port map (
            O => \N__29547\,
            I => \N__29544\
        );

    \I__4751\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29541\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29538\
        );

    \I__4749\ : Span4Mux_v
    port map (
            O => \N__29538\,
            I => \N__29535\
        );

    \I__4748\ : Sp12to4
    port map (
            O => \N__29535\,
            I => \N__29532\
        );

    \I__4747\ : Span12Mux_h
    port map (
            O => \N__29532\,
            I => \N__29529\
        );

    \I__4746\ : Odrv12
    port map (
            O => \N__29529\,
            I => \RAM_DATA_in_0\
        );

    \I__4745\ : InMux
    port map (
            O => \N__29526\,
            I => \N__29523\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__29523\,
            I => \N__29520\
        );

    \I__4743\ : Sp12to4
    port map (
            O => \N__29520\,
            I => \N__29517\
        );

    \I__4742\ : Odrv12
    port map (
            O => \N__29517\,
            I => \spi_data_misoZ0Z_0\
        );

    \I__4741\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29511\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__29511\,
            I => \N__29508\
        );

    \I__4739\ : Span12Mux_h
    port map (
            O => \N__29508\,
            I => \N__29505\
        );

    \I__4738\ : Span12Mux_v
    port map (
            O => \N__29505\,
            I => \N__29502\
        );

    \I__4737\ : Odrv12
    port map (
            O => \N__29502\,
            I => \RAM_DATA_in_9\
        );

    \I__4736\ : InMux
    port map (
            O => \N__29499\,
            I => \N__29496\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__29496\,
            I => \N__29493\
        );

    \I__4734\ : Sp12to4
    port map (
            O => \N__29493\,
            I => \N__29490\
        );

    \I__4733\ : Span12Mux_v
    port map (
            O => \N__29490\,
            I => \N__29487\
        );

    \I__4732\ : Span12Mux_h
    port map (
            O => \N__29487\,
            I => \N__29484\
        );

    \I__4731\ : Odrv12
    port map (
            O => \N__29484\,
            I => \RAM_DATA_in_1\
        );

    \I__4730\ : InMux
    port map (
            O => \N__29481\,
            I => \N__29478\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__29478\,
            I => \N__29475\
        );

    \I__4728\ : Span4Mux_h
    port map (
            O => \N__29475\,
            I => \N__29472\
        );

    \I__4727\ : Odrv4
    port map (
            O => \N__29472\,
            I => \spi_data_misoZ0Z_1\
        );

    \I__4726\ : InMux
    port map (
            O => \N__29469\,
            I => \N__29466\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__29466\,
            I => \N__29463\
        );

    \I__4724\ : Span4Mux_h
    port map (
            O => \N__29463\,
            I => \N__29460\
        );

    \I__4723\ : Span4Mux_h
    port map (
            O => \N__29460\,
            I => \N__29457\
        );

    \I__4722\ : Sp12to4
    port map (
            O => \N__29457\,
            I => \N__29454\
        );

    \I__4721\ : Span12Mux_v
    port map (
            O => \N__29454\,
            I => \N__29451\
        );

    \I__4720\ : Span12Mux_v
    port map (
            O => \N__29451\,
            I => \N__29448\
        );

    \I__4719\ : Odrv12
    port map (
            O => \N__29448\,
            I => \RAM_DATA_in_10\
        );

    \I__4718\ : CascadeMux
    port map (
            O => \N__29445\,
            I => \N__29442\
        );

    \I__4717\ : InMux
    port map (
            O => \N__29442\,
            I => \N__29439\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__29439\,
            I => \N__29436\
        );

    \I__4715\ : Span4Mux_v
    port map (
            O => \N__29436\,
            I => \N__29433\
        );

    \I__4714\ : Span4Mux_v
    port map (
            O => \N__29433\,
            I => \N__29430\
        );

    \I__4713\ : Sp12to4
    port map (
            O => \N__29430\,
            I => \N__29427\
        );

    \I__4712\ : Span12Mux_h
    port map (
            O => \N__29427\,
            I => \N__29424\
        );

    \I__4711\ : Odrv12
    port map (
            O => \N__29424\,
            I => \RAM_DATA_in_2\
        );

    \I__4710\ : InMux
    port map (
            O => \N__29421\,
            I => \N__29418\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__29418\,
            I => \N__29415\
        );

    \I__4708\ : Span4Mux_h
    port map (
            O => \N__29415\,
            I => \N__29412\
        );

    \I__4707\ : Odrv4
    port map (
            O => \N__29412\,
            I => \spi_data_misoZ0Z_2\
        );

    \I__4706\ : InMux
    port map (
            O => \N__29409\,
            I => \N__29406\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__29406\,
            I => \N__29403\
        );

    \I__4704\ : Span4Mux_h
    port map (
            O => \N__29403\,
            I => \N__29400\
        );

    \I__4703\ : Odrv4
    port map (
            O => \N__29400\,
            I => \sEEPoffZ0Z_11\
        );

    \I__4702\ : InMux
    port map (
            O => \N__29397\,
            I => \N__29394\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__29394\,
            I => \N__29391\
        );

    \I__4700\ : Span4Mux_v
    port map (
            O => \N__29391\,
            I => \N__29388\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__29388\,
            I => \sEEPoffZ0Z_12\
        );

    \I__4698\ : InMux
    port map (
            O => \N__29385\,
            I => \N__29382\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__29382\,
            I => \N__29379\
        );

    \I__4696\ : Odrv4
    port map (
            O => \N__29379\,
            I => \sEEPoffZ0Z_13\
        );

    \I__4695\ : InMux
    port map (
            O => \N__29376\,
            I => \N__29373\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__29373\,
            I => \N__29370\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__29370\,
            I => \sEEPoffZ0Z_14\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__29367\,
            I => \N__29364\
        );

    \I__4691\ : InMux
    port map (
            O => \N__29364\,
            I => \N__29361\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__29361\,
            I => \N__29358\
        );

    \I__4689\ : Odrv4
    port map (
            O => \N__29358\,
            I => \sEEPoffZ0Z_15\
        );

    \I__4688\ : InMux
    port map (
            O => \N__29355\,
            I => \N__29352\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__29352\,
            I => \N__29349\
        );

    \I__4686\ : Odrv4
    port map (
            O => \N__29349\,
            I => \sEEPoffZ0Z_8\
        );

    \I__4685\ : InMux
    port map (
            O => \N__29346\,
            I => \N__29343\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__29343\,
            I => \N__29340\
        );

    \I__4683\ : Odrv12
    port map (
            O => \N__29340\,
            I => \sEEPoffZ0Z_9\
        );

    \I__4682\ : CEMux
    port map (
            O => \N__29337\,
            I => \N__29334\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__29334\,
            I => \N__29331\
        );

    \I__4680\ : Span4Mux_v
    port map (
            O => \N__29331\,
            I => \N__29328\
        );

    \I__4679\ : Span4Mux_h
    port map (
            O => \N__29328\,
            I => \N__29325\
        );

    \I__4678\ : Odrv4
    port map (
            O => \N__29325\,
            I => \sAddress_RNIA6242_1Z0Z_2\
        );

    \I__4677\ : InMux
    port map (
            O => \N__29322\,
            I => \bfn_12_15_0_\
        );

    \I__4676\ : InMux
    port map (
            O => \N__29319\,
            I => \sCounterADC_cry_0\
        );

    \I__4675\ : InMux
    port map (
            O => \N__29316\,
            I => \N__29313\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__29313\,
            I => \N__29310\
        );

    \I__4673\ : Odrv12
    port map (
            O => \N__29310\,
            I => \sEEPoffZ0Z_0\
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__29307\,
            I => \N__29304\
        );

    \I__4671\ : InMux
    port map (
            O => \N__29304\,
            I => \N__29301\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__29301\,
            I => \N__29298\
        );

    \I__4669\ : Span4Mux_h
    port map (
            O => \N__29298\,
            I => \N__29295\
        );

    \I__4668\ : Odrv4
    port map (
            O => \N__29295\,
            I => \sEEPoffZ0Z_1\
        );

    \I__4667\ : InMux
    port map (
            O => \N__29292\,
            I => \N__29289\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__29289\,
            I => \N__29286\
        );

    \I__4665\ : Odrv4
    port map (
            O => \N__29286\,
            I => \sEEPoffZ0Z_2\
        );

    \I__4664\ : InMux
    port map (
            O => \N__29283\,
            I => \N__29280\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__29280\,
            I => \N__29277\
        );

    \I__4662\ : Odrv4
    port map (
            O => \N__29277\,
            I => \sEEPoffZ0Z_3\
        );

    \I__4661\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29271\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__29271\,
            I => \N__29268\
        );

    \I__4659\ : Odrv4
    port map (
            O => \N__29268\,
            I => \sEEPoffZ0Z_4\
        );

    \I__4658\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29262\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__29262\,
            I => \N__29259\
        );

    \I__4656\ : Odrv12
    port map (
            O => \N__29259\,
            I => \sEEPoffZ0Z_5\
        );

    \I__4655\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29253\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__29253\,
            I => \N__29250\
        );

    \I__4653\ : Odrv12
    port map (
            O => \N__29250\,
            I => \sEEPoffZ0Z_6\
        );

    \I__4652\ : InMux
    port map (
            O => \N__29247\,
            I => \N__29244\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__29244\,
            I => \N__29241\
        );

    \I__4650\ : Odrv12
    port map (
            O => \N__29241\,
            I => \sEEPoffZ0Z_7\
        );

    \I__4649\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29235\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__29235\,
            I => \N__29232\
        );

    \I__4647\ : Odrv12
    port map (
            O => \N__29232\,
            I => \sEEPoffZ0Z_10\
        );

    \I__4646\ : InMux
    port map (
            O => \N__29229\,
            I => \N__29226\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__29226\,
            I => \N__29223\
        );

    \I__4644\ : Odrv12
    port map (
            O => \N__29223\,
            I => \spi_slave_inst.un1_spointer11_2_0_a2_0_6_4\
        );

    \I__4643\ : CascadeMux
    port map (
            O => \N__29220\,
            I => \spi_slave_inst.un1_spointer11_2_0_a2_0_6_5_cascade_\
        );

    \I__4642\ : InMux
    port map (
            O => \N__29217\,
            I => \N__29214\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__29214\,
            I => \N__29210\
        );

    \I__4640\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29207\
        );

    \I__4639\ : Span4Mux_h
    port map (
            O => \N__29210\,
            I => \N__29202\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__29207\,
            I => \N__29202\
        );

    \I__4637\ : Odrv4
    port map (
            O => \N__29202\,
            I => un1_spointer11_2_0
        );

    \I__4636\ : CascadeMux
    port map (
            O => \N__29199\,
            I => \N_285_cascade_\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__29196\,
            I => \N__29193\
        );

    \I__4634\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29185\
        );

    \I__4633\ : InMux
    port map (
            O => \N__29192\,
            I => \N__29180\
        );

    \I__4632\ : InMux
    port map (
            O => \N__29191\,
            I => \N__29180\
        );

    \I__4631\ : InMux
    port map (
            O => \N__29190\,
            I => \N__29177\
        );

    \I__4630\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29173\
        );

    \I__4629\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29170\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__29185\,
            I => \N__29167\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__29180\,
            I => \N__29162\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__29177\,
            I => \N__29162\
        );

    \I__4625\ : InMux
    port map (
            O => \N__29176\,
            I => \N__29159\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__29173\,
            I => \sPointerZ0Z_0\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__29170\,
            I => \sPointerZ0Z_0\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__29167\,
            I => \sPointerZ0Z_0\
        );

    \I__4621\ : Odrv4
    port map (
            O => \N__29162\,
            I => \sPointerZ0Z_0\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__29159\,
            I => \sPointerZ0Z_0\
        );

    \I__4619\ : CascadeMux
    port map (
            O => \N__29148\,
            I => \N_116_cascade_\
        );

    \I__4618\ : InMux
    port map (
            O => \N__29145\,
            I => \N__29141\
        );

    \I__4617\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29138\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__29141\,
            I => \N_159\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__29138\,
            I => \N_159\
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__29133\,
            I => \N_117_cascade_\
        );

    \I__4613\ : InMux
    port map (
            O => \N__29130\,
            I => \N__29124\
        );

    \I__4612\ : InMux
    port map (
            O => \N__29129\,
            I => \N__29121\
        );

    \I__4611\ : InMux
    port map (
            O => \N__29128\,
            I => \N__29118\
        );

    \I__4610\ : InMux
    port map (
            O => \N__29127\,
            I => \N__29115\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__29124\,
            I => \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__29121\,
            I => \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__29118\,
            I => \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__29115\,
            I => \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1\
        );

    \I__4605\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29090\
        );

    \I__4604\ : InMux
    port map (
            O => \N__29105\,
            I => \N__29085\
        );

    \I__4603\ : InMux
    port map (
            O => \N__29104\,
            I => \N__29085\
        );

    \I__4602\ : InMux
    port map (
            O => \N__29103\,
            I => \N__29073\
        );

    \I__4601\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29073\
        );

    \I__4600\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29073\
        );

    \I__4599\ : InMux
    port map (
            O => \N__29100\,
            I => \N__29073\
        );

    \I__4598\ : InMux
    port map (
            O => \N__29099\,
            I => \N__29073\
        );

    \I__4597\ : InMux
    port map (
            O => \N__29098\,
            I => \N__29064\
        );

    \I__4596\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29064\
        );

    \I__4595\ : InMux
    port map (
            O => \N__29096\,
            I => \N__29064\
        );

    \I__4594\ : InMux
    port map (
            O => \N__29095\,
            I => \N__29064\
        );

    \I__4593\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29061\
        );

    \I__4592\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29057\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__29090\,
            I => \N__29054\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__29085\,
            I => \N__29051\
        );

    \I__4589\ : InMux
    port map (
            O => \N__29084\,
            I => \N__29048\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__29073\,
            I => \N__29045\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__29064\,
            I => \N__29042\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__29061\,
            I => \N__29037\
        );

    \I__4585\ : InMux
    port map (
            O => \N__29060\,
            I => \N__29034\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__29057\,
            I => \N__29031\
        );

    \I__4583\ : Span4Mux_v
    port map (
            O => \N__29054\,
            I => \N__29024\
        );

    \I__4582\ : Span4Mux_v
    port map (
            O => \N__29051\,
            I => \N__29024\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__29048\,
            I => \N__29024\
        );

    \I__4580\ : Span4Mux_v
    port map (
            O => \N__29045\,
            I => \N__29019\
        );

    \I__4579\ : Span4Mux_h
    port map (
            O => \N__29042\,
            I => \N__29019\
        );

    \I__4578\ : InMux
    port map (
            O => \N__29041\,
            I => \N__29014\
        );

    \I__4577\ : InMux
    port map (
            O => \N__29040\,
            I => \N__29014\
        );

    \I__4576\ : Span12Mux_h
    port map (
            O => \N__29037\,
            I => \N__29011\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__29034\,
            I => \N__29006\
        );

    \I__4574\ : Span12Mux_v
    port map (
            O => \N__29031\,
            I => \N__29006\
        );

    \I__4573\ : Span4Mux_h
    port map (
            O => \N__29024\,
            I => \N__29003\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__29019\,
            I => \N__29000\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__29014\,
            I => \sEETrigInternalZ0\
        );

    \I__4570\ : Odrv12
    port map (
            O => \N__29011\,
            I => \sEETrigInternalZ0\
        );

    \I__4569\ : Odrv12
    port map (
            O => \N__29006\,
            I => \sEETrigInternalZ0\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__29003\,
            I => \sEETrigInternalZ0\
        );

    \I__4567\ : Odrv4
    port map (
            O => \N__29000\,
            I => \sEETrigInternalZ0\
        );

    \I__4566\ : CEMux
    port map (
            O => \N__28989\,
            I => \N__28985\
        );

    \I__4565\ : CEMux
    port map (
            O => \N__28988\,
            I => \N__28982\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__28985\,
            I => \N__28977\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__28982\,
            I => \N__28977\
        );

    \I__4562\ : Sp12to4
    port map (
            O => \N__28977\,
            I => \N__28974\
        );

    \I__4561\ : Odrv12
    port map (
            O => \N__28974\,
            I => \sDAC_mem_23_1_sqmuxa\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__28971\,
            I => \N_275_cascade_\
        );

    \I__4559\ : CascadeMux
    port map (
            O => \N__28968\,
            I => \N_360_cascade_\
        );

    \I__4558\ : InMux
    port map (
            O => \N__28965\,
            I => \N__28962\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__28962\,
            I => \N_269\
        );

    \I__4556\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28956\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__28956\,
            I => \N__28953\
        );

    \I__4554\ : Span4Mux_h
    port map (
            O => \N__28953\,
            I => \N__28950\
        );

    \I__4553\ : Span4Mux_h
    port map (
            O => \N__28950\,
            I => \N__28947\
        );

    \I__4552\ : Odrv4
    port map (
            O => \N__28947\,
            I => \N_132\
        );

    \I__4551\ : CEMux
    port map (
            O => \N__28944\,
            I => \N__28941\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__28941\,
            I => \N__28938\
        );

    \I__4549\ : Odrv12
    port map (
            O => \N__28938\,
            I => \sAddress_RNIA6242_0Z0Z_0\
        );

    \I__4548\ : CascadeMux
    port map (
            O => \N__28935\,
            I => \N__28932\
        );

    \I__4547\ : InMux
    port map (
            O => \N__28932\,
            I => \N__28929\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__28929\,
            I => un1_spointer11_7_0_tz
        );

    \I__4545\ : CascadeMux
    port map (
            O => \N__28926\,
            I => \un1_spointer11_7_0_tz_cascade_\
        );

    \I__4544\ : CEMux
    port map (
            O => \N__28923\,
            I => \N__28920\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__28920\,
            I => \N__28917\
        );

    \I__4542\ : Odrv12
    port map (
            O => \N__28917\,
            I => \sAddress_RNID9242Z0Z_3\
        );

    \I__4541\ : CascadeMux
    port map (
            O => \N__28914\,
            I => \un1_spointer11_5_0_2_cascade_\
        );

    \I__4540\ : CEMux
    port map (
            O => \N__28911\,
            I => \N__28908\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__28908\,
            I => \N__28905\
        );

    \I__4538\ : Span4Mux_v
    port map (
            O => \N__28905\,
            I => \N__28902\
        );

    \I__4537\ : Odrv4
    port map (
            O => \N__28902\,
            I => \sAddress_RNIA6242_0Z0Z_2\
        );

    \I__4536\ : InMux
    port map (
            O => \N__28899\,
            I => \N__28896\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__28896\,
            I => \N__28893\
        );

    \I__4534\ : Odrv4
    port map (
            O => \N__28893\,
            I => \sDAC_dataZ0Z_0\
        );

    \I__4533\ : InMux
    port map (
            O => \N__28890\,
            I => \N__28887\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__28887\,
            I => \N__28884\
        );

    \I__4531\ : Span4Mux_h
    port map (
            O => \N__28884\,
            I => \N__28881\
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__28881\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_0\
        );

    \I__4529\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28875\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__28875\,
            I => \N__28872\
        );

    \I__4527\ : Span4Mux_h
    port map (
            O => \N__28872\,
            I => \N__28869\
        );

    \I__4526\ : Odrv4
    port map (
            O => \N__28869\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_7\
        );

    \I__4525\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28863\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__28863\,
            I => \N__28860\
        );

    \I__4523\ : Span4Mux_h
    port map (
            O => \N__28860\,
            I => \N__28857\
        );

    \I__4522\ : Odrv4
    port map (
            O => \N__28857\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_8\
        );

    \I__4521\ : InMux
    port map (
            O => \N__28854\,
            I => \N__28851\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__28851\,
            I => \N__28848\
        );

    \I__4519\ : Span4Mux_v
    port map (
            O => \N__28848\,
            I => \N__28845\
        );

    \I__4518\ : Odrv4
    port map (
            O => \N__28845\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_9\
        );

    \I__4517\ : CEMux
    port map (
            O => \N__28842\,
            I => \N__28838\
        );

    \I__4516\ : CEMux
    port map (
            O => \N__28841\,
            I => \N__28834\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__28838\,
            I => \N__28831\
        );

    \I__4514\ : CascadeMux
    port map (
            O => \N__28837\,
            I => \N__28828\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__28834\,
            I => \N__28825\
        );

    \I__4512\ : Span4Mux_v
    port map (
            O => \N__28831\,
            I => \N__28822\
        );

    \I__4511\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28819\
        );

    \I__4510\ : Odrv12
    port map (
            O => \N__28825\,
            I => \spi_master_inst.spi_data_path_u1.tx_ready_iZ0\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__28822\,
            I => \spi_master_inst.spi_data_path_u1.tx_ready_iZ0\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__28819\,
            I => \spi_master_inst.spi_data_path_u1.tx_ready_iZ0\
        );

    \I__4507\ : InMux
    port map (
            O => \N__28812\,
            I => \N__28809\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__28809\,
            I => \N__28806\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__28806\,
            I => \N__28802\
        );

    \I__4504\ : InMux
    port map (
            O => \N__28805\,
            I => \N__28799\
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__28802\,
            I => \spi_slave_inst.rx_done_reg1_iZ0\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__28799\,
            I => \spi_slave_inst.rx_done_reg1_iZ0\
        );

    \I__4501\ : InMux
    port map (
            O => \N__28794\,
            I => \N__28789\
        );

    \I__4500\ : InMux
    port map (
            O => \N__28793\,
            I => \N__28784\
        );

    \I__4499\ : InMux
    port map (
            O => \N__28792\,
            I => \N__28784\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__28789\,
            I => \N__28781\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__28784\,
            I => \N__28778\
        );

    \I__4496\ : Span4Mux_h
    port map (
            O => \N__28781\,
            I => \N__28775\
        );

    \I__4495\ : Span12Mux_v
    port map (
            O => \N__28778\,
            I => \N__28772\
        );

    \I__4494\ : Odrv4
    port map (
            O => \N__28775\,
            I => \spi_slave_inst.rx_done_reg2_iZ0\
        );

    \I__4493\ : Odrv12
    port map (
            O => \N__28772\,
            I => \spi_slave_inst.rx_done_reg2_iZ0\
        );

    \I__4492\ : CEMux
    port map (
            O => \N__28767\,
            I => \N__28764\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__28764\,
            I => \spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541\
        );

    \I__4490\ : InMux
    port map (
            O => \N__28761\,
            I => \N__28758\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__28758\,
            I => \N__28755\
        );

    \I__4488\ : Odrv12
    port map (
            O => \N__28755\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_10\
        );

    \I__4487\ : InMux
    port map (
            O => \N__28752\,
            I => \N__28749\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__28749\,
            I => \N__28746\
        );

    \I__4485\ : Span4Mux_v
    port map (
            O => \N__28746\,
            I => \N__28743\
        );

    \I__4484\ : Span4Mux_h
    port map (
            O => \N__28743\,
            I => \N__28740\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__28740\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_13\
        );

    \I__4482\ : InMux
    port map (
            O => \N__28737\,
            I => \N__28734\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__28734\,
            I => \N__28731\
        );

    \I__4480\ : Odrv4
    port map (
            O => \N__28731\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_4\
        );

    \I__4479\ : InMux
    port map (
            O => \N__28728\,
            I => \N__28725\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__28725\,
            I => \N__28722\
        );

    \I__4477\ : Odrv12
    port map (
            O => \N__28722\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_5\
        );

    \I__4476\ : InMux
    port map (
            O => \N__28719\,
            I => \N__28716\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__28716\,
            I => \N__28713\
        );

    \I__4474\ : Sp12to4
    port map (
            O => \N__28713\,
            I => \N__28710\
        );

    \I__4473\ : Span12Mux_v
    port map (
            O => \N__28710\,
            I => \N__28707\
        );

    \I__4472\ : Span12Mux_h
    port map (
            O => \N__28707\,
            I => \N__28704\
        );

    \I__4471\ : Odrv12
    port map (
            O => \N__28704\,
            I => spi_sclk_ft_c
        );

    \I__4470\ : IoInMux
    port map (
            O => \N__28701\,
            I => \N__28698\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__28698\,
            I => \N__28695\
        );

    \I__4468\ : Span4Mux_s3_v
    port map (
            O => \N__28695\,
            I => \N__28692\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__28692\,
            I => spi_sclk
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__28689\,
            I => \N__28686\
        );

    \I__4465\ : InMux
    port map (
            O => \N__28686\,
            I => \N__28683\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__28683\,
            I => \N__28680\
        );

    \I__4463\ : Span4Mux_v
    port map (
            O => \N__28680\,
            I => \N__28677\
        );

    \I__4462\ : Span4Mux_h
    port map (
            O => \N__28677\,
            I => \N__28674\
        );

    \I__4461\ : Span4Mux_h
    port map (
            O => \N__28674\,
            I => \N__28670\
        );

    \I__4460\ : InMux
    port map (
            O => \N__28673\,
            I => \N__28667\
        );

    \I__4459\ : Odrv4
    port map (
            O => \N__28670\,
            I => \sRAM_pointer_readZ0Z_3\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__28667\,
            I => \sRAM_pointer_readZ0Z_3\
        );

    \I__4457\ : IoInMux
    port map (
            O => \N__28662\,
            I => \N__28659\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__28659\,
            I => \N__28656\
        );

    \I__4455\ : Span12Mux_s9_v
    port map (
            O => \N__28656\,
            I => \N__28653\
        );

    \I__4454\ : Odrv12
    port map (
            O => \N__28653\,
            I => \RAM_ADD_c_3\
        );

    \I__4453\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28647\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__28647\,
            I => \N__28644\
        );

    \I__4451\ : Span4Mux_v
    port map (
            O => \N__28644\,
            I => \N__28641\
        );

    \I__4450\ : Span4Mux_h
    port map (
            O => \N__28641\,
            I => \N__28638\
        );

    \I__4449\ : Span4Mux_h
    port map (
            O => \N__28638\,
            I => \N__28634\
        );

    \I__4448\ : InMux
    port map (
            O => \N__28637\,
            I => \N__28631\
        );

    \I__4447\ : Odrv4
    port map (
            O => \N__28634\,
            I => \sRAM_pointer_readZ0Z_4\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__28631\,
            I => \sRAM_pointer_readZ0Z_4\
        );

    \I__4445\ : IoInMux
    port map (
            O => \N__28626\,
            I => \N__28623\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__28623\,
            I => \N__28620\
        );

    \I__4443\ : Span4Mux_s1_v
    port map (
            O => \N__28620\,
            I => \N__28617\
        );

    \I__4442\ : Span4Mux_v
    port map (
            O => \N__28617\,
            I => \N__28614\
        );

    \I__4441\ : Span4Mux_v
    port map (
            O => \N__28614\,
            I => \N__28611\
        );

    \I__4440\ : Sp12to4
    port map (
            O => \N__28611\,
            I => \N__28608\
        );

    \I__4439\ : Odrv12
    port map (
            O => \N__28608\,
            I => \RAM_ADD_c_4\
        );

    \I__4438\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28602\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__28602\,
            I => \N__28599\
        );

    \I__4436\ : Span4Mux_v
    port map (
            O => \N__28599\,
            I => \N__28596\
        );

    \I__4435\ : Span4Mux_h
    port map (
            O => \N__28596\,
            I => \N__28593\
        );

    \I__4434\ : Span4Mux_h
    port map (
            O => \N__28593\,
            I => \N__28589\
        );

    \I__4433\ : InMux
    port map (
            O => \N__28592\,
            I => \N__28586\
        );

    \I__4432\ : Odrv4
    port map (
            O => \N__28589\,
            I => \sRAM_pointer_readZ0Z_5\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__28586\,
            I => \sRAM_pointer_readZ0Z_5\
        );

    \I__4430\ : IoInMux
    port map (
            O => \N__28581\,
            I => \N__28578\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__28578\,
            I => \N__28575\
        );

    \I__4428\ : Span4Mux_s2_h
    port map (
            O => \N__28575\,
            I => \N__28572\
        );

    \I__4427\ : Span4Mux_v
    port map (
            O => \N__28572\,
            I => \N__28569\
        );

    \I__4426\ : Sp12to4
    port map (
            O => \N__28569\,
            I => \N__28566\
        );

    \I__4425\ : Span12Mux_s9_h
    port map (
            O => \N__28566\,
            I => \N__28563\
        );

    \I__4424\ : Odrv12
    port map (
            O => \N__28563\,
            I => \RAM_ADD_c_5\
        );

    \I__4423\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28557\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__28557\,
            I => \N__28554\
        );

    \I__4421\ : Span4Mux_v
    port map (
            O => \N__28554\,
            I => \N__28551\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__28551\,
            I => \N__28548\
        );

    \I__4419\ : Span4Mux_h
    port map (
            O => \N__28548\,
            I => \N__28544\
        );

    \I__4418\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28541\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__28544\,
            I => \sRAM_pointer_readZ0Z_6\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__28541\,
            I => \sRAM_pointer_readZ0Z_6\
        );

    \I__4415\ : IoInMux
    port map (
            O => \N__28536\,
            I => \N__28533\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__28533\,
            I => \N__28530\
        );

    \I__4413\ : Span4Mux_s2_h
    port map (
            O => \N__28530\,
            I => \N__28527\
        );

    \I__4412\ : Span4Mux_h
    port map (
            O => \N__28527\,
            I => \N__28524\
        );

    \I__4411\ : Span4Mux_h
    port map (
            O => \N__28524\,
            I => \N__28521\
        );

    \I__4410\ : Sp12to4
    port map (
            O => \N__28521\,
            I => \N__28518\
        );

    \I__4409\ : Span12Mux_s8_v
    port map (
            O => \N__28518\,
            I => \N__28515\
        );

    \I__4408\ : Odrv12
    port map (
            O => \N__28515\,
            I => \RAM_ADD_c_6\
        );

    \I__4407\ : CascadeMux
    port map (
            O => \N__28512\,
            I => \N__28509\
        );

    \I__4406\ : InMux
    port map (
            O => \N__28509\,
            I => \N__28506\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__28506\,
            I => \N__28503\
        );

    \I__4404\ : Sp12to4
    port map (
            O => \N__28503\,
            I => \N__28500\
        );

    \I__4403\ : Span12Mux_v
    port map (
            O => \N__28500\,
            I => \N__28496\
        );

    \I__4402\ : InMux
    port map (
            O => \N__28499\,
            I => \N__28493\
        );

    \I__4401\ : Odrv12
    port map (
            O => \N__28496\,
            I => \sRAM_pointer_readZ0Z_7\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__28493\,
            I => \sRAM_pointer_readZ0Z_7\
        );

    \I__4399\ : IoInMux
    port map (
            O => \N__28488\,
            I => \N__28485\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__28485\,
            I => \N__28482\
        );

    \I__4397\ : Span4Mux_s3_h
    port map (
            O => \N__28482\,
            I => \N__28479\
        );

    \I__4396\ : Span4Mux_h
    port map (
            O => \N__28479\,
            I => \N__28476\
        );

    \I__4395\ : Span4Mux_h
    port map (
            O => \N__28476\,
            I => \N__28473\
        );

    \I__4394\ : Sp12to4
    port map (
            O => \N__28473\,
            I => \N__28470\
        );

    \I__4393\ : Span12Mux_s8_v
    port map (
            O => \N__28470\,
            I => \N__28467\
        );

    \I__4392\ : Odrv12
    port map (
            O => \N__28467\,
            I => \RAM_ADD_c_7\
        );

    \I__4391\ : InMux
    port map (
            O => \N__28464\,
            I => \N__28461\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__28461\,
            I => \N__28458\
        );

    \I__4389\ : Span4Mux_v
    port map (
            O => \N__28458\,
            I => \N__28455\
        );

    \I__4388\ : Span4Mux_h
    port map (
            O => \N__28455\,
            I => \N__28452\
        );

    \I__4387\ : Span4Mux_h
    port map (
            O => \N__28452\,
            I => \N__28448\
        );

    \I__4386\ : InMux
    port map (
            O => \N__28451\,
            I => \N__28445\
        );

    \I__4385\ : Odrv4
    port map (
            O => \N__28448\,
            I => \sRAM_pointer_readZ0Z_8\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__28445\,
            I => \sRAM_pointer_readZ0Z_8\
        );

    \I__4383\ : IoInMux
    port map (
            O => \N__28440\,
            I => \N__28437\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__28437\,
            I => \N__28434\
        );

    \I__4381\ : IoSpan4Mux
    port map (
            O => \N__28434\,
            I => \N__28431\
        );

    \I__4380\ : Span4Mux_s3_h
    port map (
            O => \N__28431\,
            I => \N__28428\
        );

    \I__4379\ : Sp12to4
    port map (
            O => \N__28428\,
            I => \N__28425\
        );

    \I__4378\ : Span12Mux_h
    port map (
            O => \N__28425\,
            I => \N__28422\
        );

    \I__4377\ : Odrv12
    port map (
            O => \N__28422\,
            I => \RAM_ADD_c_8\
        );

    \I__4376\ : CascadeMux
    port map (
            O => \N__28419\,
            I => \N__28416\
        );

    \I__4375\ : InMux
    port map (
            O => \N__28416\,
            I => \N__28413\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__28413\,
            I => \N__28410\
        );

    \I__4373\ : Span4Mux_v
    port map (
            O => \N__28410\,
            I => \N__28407\
        );

    \I__4372\ : Sp12to4
    port map (
            O => \N__28407\,
            I => \N__28404\
        );

    \I__4371\ : Span12Mux_h
    port map (
            O => \N__28404\,
            I => \N__28400\
        );

    \I__4370\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28397\
        );

    \I__4369\ : Odrv12
    port map (
            O => \N__28400\,
            I => \sRAM_pointer_readZ0Z_9\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__28397\,
            I => \sRAM_pointer_readZ0Z_9\
        );

    \I__4367\ : IoInMux
    port map (
            O => \N__28392\,
            I => \N__28389\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__28389\,
            I => \N__28386\
        );

    \I__4365\ : IoSpan4Mux
    port map (
            O => \N__28386\,
            I => \N__28383\
        );

    \I__4364\ : IoSpan4Mux
    port map (
            O => \N__28383\,
            I => \N__28380\
        );

    \I__4363\ : Sp12to4
    port map (
            O => \N__28380\,
            I => \N__28377\
        );

    \I__4362\ : Span12Mux_s7_h
    port map (
            O => \N__28377\,
            I => \N__28374\
        );

    \I__4361\ : Odrv12
    port map (
            O => \N__28374\,
            I => \RAM_ADD_c_9\
        );

    \I__4360\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28368\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__28368\,
            I => \N__28365\
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__28365\,
            I => \N_102\
        );

    \I__4357\ : IoInMux
    port map (
            O => \N__28362\,
            I => \N__28359\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__28359\,
            I => \N__28356\
        );

    \I__4355\ : IoSpan4Mux
    port map (
            O => \N__28356\,
            I => \N__28353\
        );

    \I__4354\ : Sp12to4
    port map (
            O => \N__28353\,
            I => \N__28349\
        );

    \I__4353\ : InMux
    port map (
            O => \N__28352\,
            I => \N__28346\
        );

    \I__4352\ : Span12Mux_s7_h
    port map (
            O => \N__28349\,
            I => \N__28343\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__28346\,
            I => \N__28340\
        );

    \I__4350\ : Span12Mux_v
    port map (
            O => \N__28343\,
            I => \N__28337\
        );

    \I__4349\ : Span4Mux_h
    port map (
            O => \N__28340\,
            I => \N__28334\
        );

    \I__4348\ : Odrv12
    port map (
            O => \N__28337\,
            I => \RAM_DATA_cl_15Z0Z_15\
        );

    \I__4347\ : Odrv4
    port map (
            O => \N__28334\,
            I => \RAM_DATA_cl_15Z0Z_15\
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__28329\,
            I => \N_96_cascade_\
        );

    \I__4345\ : IoInMux
    port map (
            O => \N__28326\,
            I => \N__28323\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__28323\,
            I => \N__28320\
        );

    \I__4343\ : IoSpan4Mux
    port map (
            O => \N__28320\,
            I => \N__28317\
        );

    \I__4342\ : Span4Mux_s2_v
    port map (
            O => \N__28317\,
            I => \N__28314\
        );

    \I__4341\ : Sp12to4
    port map (
            O => \N__28314\,
            I => \N__28311\
        );

    \I__4340\ : Span12Mux_s10_v
    port map (
            O => \N__28311\,
            I => \N__28307\
        );

    \I__4339\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28304\
        );

    \I__4338\ : Odrv12
    port map (
            O => \N__28307\,
            I => \RAM_DATA_cl_8Z0Z_15\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__28304\,
            I => \RAM_DATA_cl_8Z0Z_15\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__28299\,
            I => \N__28296\
        );

    \I__4335\ : InMux
    port map (
            O => \N__28296\,
            I => \N__28293\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__28293\,
            I => \N__28290\
        );

    \I__4333\ : Sp12to4
    port map (
            O => \N__28290\,
            I => \N__28286\
        );

    \I__4332\ : InMux
    port map (
            O => \N__28289\,
            I => \N__28283\
        );

    \I__4331\ : Span12Mux_v
    port map (
            O => \N__28286\,
            I => \N__28280\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__28283\,
            I => \sRAM_pointer_readZ0Z_14\
        );

    \I__4329\ : Odrv12
    port map (
            O => \N__28280\,
            I => \sRAM_pointer_readZ0Z_14\
        );

    \I__4328\ : IoInMux
    port map (
            O => \N__28275\,
            I => \N__28272\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__28272\,
            I => \N__28269\
        );

    \I__4326\ : IoSpan4Mux
    port map (
            O => \N__28269\,
            I => \N__28266\
        );

    \I__4325\ : Span4Mux_s1_h
    port map (
            O => \N__28266\,
            I => \N__28263\
        );

    \I__4324\ : Span4Mux_h
    port map (
            O => \N__28263\,
            I => \N__28260\
        );

    \I__4323\ : Sp12to4
    port map (
            O => \N__28260\,
            I => \N__28257\
        );

    \I__4322\ : Span12Mux_v
    port map (
            O => \N__28257\,
            I => \N__28254\
        );

    \I__4321\ : Span12Mux_h
    port map (
            O => \N__28254\,
            I => \N__28251\
        );

    \I__4320\ : Odrv12
    port map (
            O => \N__28251\,
            I => \RAM_ADD_c_14\
        );

    \I__4319\ : InMux
    port map (
            O => \N__28248\,
            I => \N__28245\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__28245\,
            I => \N__28242\
        );

    \I__4317\ : Span12Mux_v
    port map (
            O => \N__28242\,
            I => \N__28238\
        );

    \I__4316\ : InMux
    port map (
            O => \N__28241\,
            I => \N__28235\
        );

    \I__4315\ : Odrv12
    port map (
            O => \N__28238\,
            I => \sRAM_pointer_readZ0Z_15\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__28235\,
            I => \sRAM_pointer_readZ0Z_15\
        );

    \I__4313\ : IoInMux
    port map (
            O => \N__28230\,
            I => \N__28227\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__28227\,
            I => \N__28224\
        );

    \I__4311\ : IoSpan4Mux
    port map (
            O => \N__28224\,
            I => \N__28221\
        );

    \I__4310\ : Span4Mux_s2_h
    port map (
            O => \N__28221\,
            I => \N__28218\
        );

    \I__4309\ : Sp12to4
    port map (
            O => \N__28218\,
            I => \N__28215\
        );

    \I__4308\ : Span12Mux_s10_h
    port map (
            O => \N__28215\,
            I => \N__28212\
        );

    \I__4307\ : Odrv12
    port map (
            O => \N__28212\,
            I => \RAM_ADD_c_15\
        );

    \I__4306\ : InMux
    port map (
            O => \N__28209\,
            I => \N__28206\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__28206\,
            I => \N__28203\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__28203\,
            I => \N__28200\
        );

    \I__4303\ : Span4Mux_h
    port map (
            O => \N__28200\,
            I => \N__28196\
        );

    \I__4302\ : InMux
    port map (
            O => \N__28199\,
            I => \N__28193\
        );

    \I__4301\ : Span4Mux_v
    port map (
            O => \N__28196\,
            I => \N__28190\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__28193\,
            I => \sRAM_pointer_readZ0Z_16\
        );

    \I__4299\ : Odrv4
    port map (
            O => \N__28190\,
            I => \sRAM_pointer_readZ0Z_16\
        );

    \I__4298\ : IoInMux
    port map (
            O => \N__28185\,
            I => \N__28182\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__28182\,
            I => \N__28179\
        );

    \I__4296\ : Span12Mux_s5_h
    port map (
            O => \N__28179\,
            I => \N__28176\
        );

    \I__4295\ : Span12Mux_v
    port map (
            O => \N__28176\,
            I => \N__28173\
        );

    \I__4294\ : Span12Mux_h
    port map (
            O => \N__28173\,
            I => \N__28170\
        );

    \I__4293\ : Span12Mux_v
    port map (
            O => \N__28170\,
            I => \N__28167\
        );

    \I__4292\ : Odrv12
    port map (
            O => \N__28167\,
            I => \RAM_ADD_c_16\
        );

    \I__4291\ : InMux
    port map (
            O => \N__28164\,
            I => \N__28161\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__28161\,
            I => \N__28158\
        );

    \I__4289\ : Span4Mux_h
    port map (
            O => \N__28158\,
            I => \N__28155\
        );

    \I__4288\ : Span4Mux_h
    port map (
            O => \N__28155\,
            I => \N__28152\
        );

    \I__4287\ : Span4Mux_v
    port map (
            O => \N__28152\,
            I => \N__28148\
        );

    \I__4286\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28145\
        );

    \I__4285\ : Odrv4
    port map (
            O => \N__28148\,
            I => \sRAM_pointer_readZ0Z_17\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__28145\,
            I => \sRAM_pointer_readZ0Z_17\
        );

    \I__4283\ : IoInMux
    port map (
            O => \N__28140\,
            I => \N__28137\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__28137\,
            I => \N__28134\
        );

    \I__4281\ : Sp12to4
    port map (
            O => \N__28134\,
            I => \N__28131\
        );

    \I__4280\ : Span12Mux_h
    port map (
            O => \N__28131\,
            I => \N__28128\
        );

    \I__4279\ : Odrv12
    port map (
            O => \N__28128\,
            I => \RAM_ADD_c_17\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__28125\,
            I => \N__28122\
        );

    \I__4277\ : InMux
    port map (
            O => \N__28122\,
            I => \N__28119\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__28119\,
            I => \N__28116\
        );

    \I__4275\ : Span4Mux_v
    port map (
            O => \N__28116\,
            I => \N__28113\
        );

    \I__4274\ : Span4Mux_h
    port map (
            O => \N__28113\,
            I => \N__28110\
        );

    \I__4273\ : Span4Mux_h
    port map (
            O => \N__28110\,
            I => \N__28106\
        );

    \I__4272\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28103\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__28106\,
            I => \sRAM_pointer_readZ0Z_18\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__28103\,
            I => \sRAM_pointer_readZ0Z_18\
        );

    \I__4269\ : IoInMux
    port map (
            O => \N__28098\,
            I => \N__28095\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__28095\,
            I => \N__28092\
        );

    \I__4267\ : Span12Mux_s5_h
    port map (
            O => \N__28092\,
            I => \N__28089\
        );

    \I__4266\ : Span12Mux_h
    port map (
            O => \N__28089\,
            I => \N__28086\
        );

    \I__4265\ : Span12Mux_v
    port map (
            O => \N__28086\,
            I => \N__28083\
        );

    \I__4264\ : Odrv12
    port map (
            O => \N__28083\,
            I => \RAM_ADD_c_18\
        );

    \I__4263\ : InMux
    port map (
            O => \N__28080\,
            I => \N__28077\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__28077\,
            I => \N__28074\
        );

    \I__4261\ : Span4Mux_v
    port map (
            O => \N__28074\,
            I => \N__28071\
        );

    \I__4260\ : Span4Mux_h
    port map (
            O => \N__28071\,
            I => \N__28068\
        );

    \I__4259\ : Span4Mux_h
    port map (
            O => \N__28068\,
            I => \N__28064\
        );

    \I__4258\ : InMux
    port map (
            O => \N__28067\,
            I => \N__28061\
        );

    \I__4257\ : Odrv4
    port map (
            O => \N__28064\,
            I => \sRAM_pointer_readZ0Z_2\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__28061\,
            I => \sRAM_pointer_readZ0Z_2\
        );

    \I__4255\ : IoInMux
    port map (
            O => \N__28056\,
            I => \N__28053\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28050\
        );

    \I__4253\ : Span4Mux_s2_v
    port map (
            O => \N__28050\,
            I => \N__28047\
        );

    \I__4252\ : Span4Mux_h
    port map (
            O => \N__28047\,
            I => \N__28044\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__28044\,
            I => \N__28041\
        );

    \I__4250\ : Odrv4
    port map (
            O => \N__28041\,
            I => \RAM_ADD_c_2\
        );

    \I__4249\ : InMux
    port map (
            O => \N__28038\,
            I => \N__28035\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__28035\,
            I => \N__28031\
        );

    \I__4247\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28028\
        );

    \I__4246\ : Span4Mux_h
    port map (
            O => \N__28031\,
            I => \N__28025\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__28028\,
            I => \sCounterRAMZ0Z_2\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__28025\,
            I => \sCounterRAMZ0Z_2\
        );

    \I__4243\ : InMux
    port map (
            O => \N__28020\,
            I => \N__28017\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__28017\,
            I => \N__28014\
        );

    \I__4241\ : Span4Mux_v
    port map (
            O => \N__28014\,
            I => \N__28010\
        );

    \I__4240\ : InMux
    port map (
            O => \N__28013\,
            I => \N__28007\
        );

    \I__4239\ : Span4Mux_h
    port map (
            O => \N__28010\,
            I => \N__28004\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__28007\,
            I => \sCounterRAMZ0Z_1\
        );

    \I__4237\ : Odrv4
    port map (
            O => \N__28004\,
            I => \sCounterRAMZ0Z_1\
        );

    \I__4236\ : CascadeMux
    port map (
            O => \N__27999\,
            I => \spi_data_miso_0_sqmuxa_2_i_o2_5_cascade_\
        );

    \I__4235\ : InMux
    port map (
            O => \N__27996\,
            I => \N__27993\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__27993\,
            I => \N__27990\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__27990\,
            I => \N__27987\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__27987\,
            I => spi_data_miso_0_sqmuxa_2_i_o2_4
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__27984\,
            I => \N_75_cascade_\
        );

    \I__4230\ : InMux
    port map (
            O => \N__27981\,
            I => \N__27975\
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__27980\,
            I => \N__27972\
        );

    \I__4228\ : InMux
    port map (
            O => \N__27979\,
            I => \N__27969\
        );

    \I__4227\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27966\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__27975\,
            I => \N__27963\
        );

    \I__4225\ : InMux
    port map (
            O => \N__27972\,
            I => \N__27960\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__27969\,
            I => \N__27957\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__27966\,
            I => \N__27953\
        );

    \I__4222\ : Span4Mux_h
    port map (
            O => \N__27963\,
            I => \N__27948\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__27960\,
            I => \N__27948\
        );

    \I__4220\ : Span4Mux_h
    port map (
            O => \N__27957\,
            I => \N__27945\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__27956\,
            I => \N__27942\
        );

    \I__4218\ : Span4Mux_h
    port map (
            O => \N__27953\,
            I => \N__27939\
        );

    \I__4217\ : Span4Mux_v
    port map (
            O => \N__27948\,
            I => \N__27936\
        );

    \I__4216\ : Span4Mux_h
    port map (
            O => \N__27945\,
            I => \N__27933\
        );

    \I__4215\ : InMux
    port map (
            O => \N__27942\,
            I => \N__27930\
        );

    \I__4214\ : Span4Mux_h
    port map (
            O => \N__27939\,
            I => \N__27927\
        );

    \I__4213\ : Span4Mux_v
    port map (
            O => \N__27936\,
            I => \N__27924\
        );

    \I__4212\ : Span4Mux_v
    port map (
            O => \N__27933\,
            I => \N__27921\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__27930\,
            I => \sSPI_MSB0LSBZ0Z1\
        );

    \I__4210\ : Odrv4
    port map (
            O => \N__27927\,
            I => \sSPI_MSB0LSBZ0Z1\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__27924\,
            I => \sSPI_MSB0LSBZ0Z1\
        );

    \I__4208\ : Odrv4
    port map (
            O => \N__27921\,
            I => \sSPI_MSB0LSBZ0Z1\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__27912\,
            I => \N__27908\
        );

    \I__4206\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27904\
        );

    \I__4205\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27901\
        );

    \I__4204\ : InMux
    port map (
            O => \N__27907\,
            I => \N__27898\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__27904\,
            I => \N__27894\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__27901\,
            I => \N__27889\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__27898\,
            I => \N__27889\
        );

    \I__4200\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27886\
        );

    \I__4199\ : Span4Mux_h
    port map (
            O => \N__27894\,
            I => \N__27883\
        );

    \I__4198\ : Span4Mux_v
    port map (
            O => \N__27889\,
            I => \N__27879\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__27886\,
            I => \N__27876\
        );

    \I__4196\ : Span4Mux_h
    port map (
            O => \N__27883\,
            I => \N__27873\
        );

    \I__4195\ : InMux
    port map (
            O => \N__27882\,
            I => \N__27870\
        );

    \I__4194\ : Span4Mux_h
    port map (
            O => \N__27879\,
            I => \N__27865\
        );

    \I__4193\ : Span4Mux_v
    port map (
            O => \N__27876\,
            I => \N__27865\
        );

    \I__4192\ : Odrv4
    port map (
            O => \N__27873\,
            I => \spi_mosi_ready_prev3_RNILKERZ0\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__27870\,
            I => \spi_mosi_ready_prev3_RNILKERZ0\
        );

    \I__4190\ : Odrv4
    port map (
            O => \N__27865\,
            I => \spi_mosi_ready_prev3_RNILKERZ0\
        );

    \I__4189\ : InMux
    port map (
            O => \N__27858\,
            I => \N__27855\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__27855\,
            I => \N_88\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__27852\,
            I => \N_88_cascade_\
        );

    \I__4186\ : IoInMux
    port map (
            O => \N__27849\,
            I => \N__27846\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__27846\,
            I => \N__27843\
        );

    \I__4184\ : Span4Mux_s1_h
    port map (
            O => \N__27843\,
            I => \N__27840\
        );

    \I__4183\ : Span4Mux_h
    port map (
            O => \N__27840\,
            I => \N__27837\
        );

    \I__4182\ : Span4Mux_h
    port map (
            O => \N__27837\,
            I => \N__27834\
        );

    \I__4181\ : Span4Mux_h
    port map (
            O => \N__27834\,
            I => \N__27831\
        );

    \I__4180\ : Span4Mux_v
    port map (
            O => \N__27831\,
            I => \N__27828\
        );

    \I__4179\ : Odrv4
    port map (
            O => \N__27828\,
            I => \N_28\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__27825\,
            I => \N_93_cascade_\
        );

    \I__4177\ : IoInMux
    port map (
            O => \N__27822\,
            I => \N__27819\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__27819\,
            I => \N__27816\
        );

    \I__4175\ : Span4Mux_s0_v
    port map (
            O => \N__27816\,
            I => \N__27813\
        );

    \I__4174\ : Span4Mux_h
    port map (
            O => \N__27813\,
            I => \N__27810\
        );

    \I__4173\ : Sp12to4
    port map (
            O => \N__27810\,
            I => \N__27807\
        );

    \I__4172\ : Span12Mux_h
    port map (
            O => \N__27807\,
            I => \N__27803\
        );

    \I__4171\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27800\
        );

    \I__4170\ : Odrv12
    port map (
            O => \N__27803\,
            I => \RAM_DATA_cl_9Z0Z_15\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__27800\,
            I => \RAM_DATA_cl_9Z0Z_15\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__27795\,
            I => \N_98_cascade_\
        );

    \I__4167\ : IoInMux
    port map (
            O => \N__27792\,
            I => \N__27789\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__27789\,
            I => \N__27786\
        );

    \I__4165\ : IoSpan4Mux
    port map (
            O => \N__27786\,
            I => \N__27783\
        );

    \I__4164\ : Span4Mux_s2_v
    port map (
            O => \N__27783\,
            I => \N__27780\
        );

    \I__4163\ : Sp12to4
    port map (
            O => \N__27780\,
            I => \N__27777\
        );

    \I__4162\ : Span12Mux_s10_v
    port map (
            O => \N__27777\,
            I => \N__27773\
        );

    \I__4161\ : InMux
    port map (
            O => \N__27776\,
            I => \N__27770\
        );

    \I__4160\ : Odrv12
    port map (
            O => \N__27773\,
            I => \RAM_DATA_clZ0Z_15\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__27770\,
            I => \RAM_DATA_clZ0Z_15\
        );

    \I__4158\ : InMux
    port map (
            O => \N__27765\,
            I => \N__27762\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__27762\,
            I => \N__27759\
        );

    \I__4156\ : Span4Mux_v
    port map (
            O => \N__27759\,
            I => \N__27756\
        );

    \I__4155\ : Span4Mux_h
    port map (
            O => \N__27756\,
            I => \N__27753\
        );

    \I__4154\ : Sp12to4
    port map (
            O => \N__27753\,
            I => \N__27750\
        );

    \I__4153\ : Span12Mux_v
    port map (
            O => \N__27750\,
            I => \N__27747\
        );

    \I__4152\ : Span12Mux_h
    port map (
            O => \N__27747\,
            I => \N__27744\
        );

    \I__4151\ : Odrv12
    port map (
            O => \N__27744\,
            I => \RAM_DATA_in_6\
        );

    \I__4150\ : CascadeMux
    port map (
            O => \N__27741\,
            I => \N__27738\
        );

    \I__4149\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27735\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27732\
        );

    \I__4147\ : Span4Mux_v
    port map (
            O => \N__27732\,
            I => \N__27729\
        );

    \I__4146\ : Sp12to4
    port map (
            O => \N__27729\,
            I => \N__27726\
        );

    \I__4145\ : Span12Mux_h
    port map (
            O => \N__27726\,
            I => \N__27723\
        );

    \I__4144\ : Odrv12
    port map (
            O => \N__27723\,
            I => \RAM_DATA_in_14\
        );

    \I__4143\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27717\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__27717\,
            I => \N__27714\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__27714\,
            I => \spi_data_misoZ0Z_6\
        );

    \I__4140\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27708\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__27708\,
            I => \N__27705\
        );

    \I__4138\ : Span4Mux_v
    port map (
            O => \N__27705\,
            I => \N__27702\
        );

    \I__4137\ : Span4Mux_h
    port map (
            O => \N__27702\,
            I => \N__27699\
        );

    \I__4136\ : Sp12to4
    port map (
            O => \N__27699\,
            I => \N__27696\
        );

    \I__4135\ : Span12Mux_v
    port map (
            O => \N__27696\,
            I => \N__27693\
        );

    \I__4134\ : Span12Mux_h
    port map (
            O => \N__27693\,
            I => \N__27690\
        );

    \I__4133\ : Odrv12
    port map (
            O => \N__27690\,
            I => \RAM_DATA_in_7\
        );

    \I__4132\ : InMux
    port map (
            O => \N__27687\,
            I => \N__27684\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__27684\,
            I => \N__27681\
        );

    \I__4130\ : Span4Mux_v
    port map (
            O => \N__27681\,
            I => \N__27678\
        );

    \I__4129\ : Sp12to4
    port map (
            O => \N__27678\,
            I => \N__27675\
        );

    \I__4128\ : Span12Mux_h
    port map (
            O => \N__27675\,
            I => \N__27672\
        );

    \I__4127\ : Odrv12
    port map (
            O => \N__27672\,
            I => \RAM_DATA_in_15\
        );

    \I__4126\ : InMux
    port map (
            O => \N__27669\,
            I => \N__27666\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__27666\,
            I => \N__27663\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__27663\,
            I => \spi_data_misoZ0Z_7\
        );

    \I__4123\ : IoInMux
    port map (
            O => \N__27660\,
            I => \N__27657\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__27657\,
            I => \N__27654\
        );

    \I__4121\ : IoSpan4Mux
    port map (
            O => \N__27654\,
            I => \N__27651\
        );

    \I__4120\ : Span4Mux_s2_h
    port map (
            O => \N__27651\,
            I => \N__27648\
        );

    \I__4119\ : Span4Mux_h
    port map (
            O => \N__27648\,
            I => \N__27645\
        );

    \I__4118\ : Sp12to4
    port map (
            O => \N__27645\,
            I => \N__27642\
        );

    \I__4117\ : Span12Mux_h
    port map (
            O => \N__27642\,
            I => \N__27639\
        );

    \I__4116\ : Odrv12
    port map (
            O => \N__27639\,
            I => \RAM_nWE_0_i\
        );

    \I__4115\ : InMux
    port map (
            O => \N__27636\,
            I => \N__27632\
        );

    \I__4114\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27629\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__27632\,
            I => \N__27626\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__27629\,
            I => \sADC_clk_prevZ0\
        );

    \I__4111\ : Odrv12
    port map (
            O => \N__27626\,
            I => \sADC_clk_prevZ0\
        );

    \I__4110\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27618\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__27618\,
            I => \N__27612\
        );

    \I__4108\ : InMux
    port map (
            O => \N__27617\,
            I => \N__27607\
        );

    \I__4107\ : InMux
    port map (
            O => \N__27616\,
            I => \N__27607\
        );

    \I__4106\ : IoInMux
    port map (
            O => \N__27615\,
            I => \N__27603\
        );

    \I__4105\ : Span4Mux_h
    port map (
            O => \N__27612\,
            I => \N__27597\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__27607\,
            I => \N__27597\
        );

    \I__4103\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27594\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__27603\,
            I => \N__27591\
        );

    \I__4101\ : InMux
    port map (
            O => \N__27602\,
            I => \N__27588\
        );

    \I__4100\ : Span4Mux_v
    port map (
            O => \N__27597\,
            I => \N__27583\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__27594\,
            I => \N__27583\
        );

    \I__4098\ : Odrv12
    port map (
            O => \N__27591\,
            I => \ADC_clk_c\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__27588\,
            I => \ADC_clk_c\
        );

    \I__4096\ : Odrv4
    port map (
            O => \N__27583\,
            I => \ADC_clk_c\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__27576\,
            I => \N__27572\
        );

    \I__4094\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27569\
        );

    \I__4093\ : InMux
    port map (
            O => \N__27572\,
            I => \N__27565\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__27569\,
            I => \N__27562\
        );

    \I__4091\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27559\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__27565\,
            I => \N__27556\
        );

    \I__4089\ : Span4Mux_h
    port map (
            O => \N__27562\,
            I => \N__27553\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__27559\,
            I => \N__27546\
        );

    \I__4087\ : Span4Mux_v
    port map (
            O => \N__27556\,
            I => \N__27546\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__27553\,
            I => \N__27546\
        );

    \I__4085\ : Odrv4
    port map (
            O => \N__27546\,
            I => \N_127\
        );

    \I__4084\ : SRMux
    port map (
            O => \N__27543\,
            I => \N__27537\
        );

    \I__4083\ : SRMux
    port map (
            O => \N__27542\,
            I => \N__27533\
        );

    \I__4082\ : SRMux
    port map (
            O => \N__27541\,
            I => \N__27530\
        );

    \I__4081\ : SRMux
    port map (
            O => \N__27540\,
            I => \N__27527\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__27537\,
            I => \N__27524\
        );

    \I__4079\ : SRMux
    port map (
            O => \N__27536\,
            I => \N__27521\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__27533\,
            I => \N__27518\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__27530\,
            I => \N__27515\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__27527\,
            I => \N__27512\
        );

    \I__4075\ : Span4Mux_h
    port map (
            O => \N__27524\,
            I => \N__27505\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__27521\,
            I => \N__27505\
        );

    \I__4073\ : Span4Mux_v
    port map (
            O => \N__27518\,
            I => \N__27505\
        );

    \I__4072\ : Span4Mux_v
    port map (
            O => \N__27515\,
            I => \N__27502\
        );

    \I__4071\ : Span4Mux_h
    port map (
            O => \N__27512\,
            I => \N__27499\
        );

    \I__4070\ : Span4Mux_v
    port map (
            O => \N__27505\,
            I => \N__27496\
        );

    \I__4069\ : Span4Mux_h
    port map (
            O => \N__27502\,
            I => \N__27491\
        );

    \I__4068\ : Span4Mux_v
    port map (
            O => \N__27499\,
            I => \N__27491\
        );

    \I__4067\ : Odrv4
    port map (
            O => \N__27496\,
            I => \N_1470_i\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__27491\,
            I => \N_1470_i\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__27486\,
            I => \N__27483\
        );

    \I__4064\ : InMux
    port map (
            O => \N__27483\,
            I => \N__27480\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__27480\,
            I => \N__27477\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__27477\,
            I => \N_86\
        );

    \I__4061\ : InMux
    port map (
            O => \N__27474\,
            I => \N__27471\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__27471\,
            I => \N__27467\
        );

    \I__4059\ : InMux
    port map (
            O => \N__27470\,
            I => \N__27464\
        );

    \I__4058\ : Span4Mux_h
    port map (
            O => \N__27467\,
            I => \N__27461\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__27464\,
            I => \sRead_dataZ0\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__27461\,
            I => \sRead_dataZ0\
        );

    \I__4055\ : InMux
    port map (
            O => \N__27456\,
            I => \N__27453\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__27453\,
            I => \N__27449\
        );

    \I__4053\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27446\
        );

    \I__4052\ : Span4Mux_h
    port map (
            O => \N__27449\,
            I => \N__27443\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__27446\,
            I => \sCounterRAMZ0Z_5\
        );

    \I__4050\ : Odrv4
    port map (
            O => \N__27443\,
            I => \sCounterRAMZ0Z_5\
        );

    \I__4049\ : InMux
    port map (
            O => \N__27438\,
            I => \N__27434\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__27437\,
            I => \N__27431\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__27434\,
            I => \N__27428\
        );

    \I__4046\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27425\
        );

    \I__4045\ : Span4Mux_h
    port map (
            O => \N__27428\,
            I => \N__27422\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__27425\,
            I => \sCounterRAMZ0Z_4\
        );

    \I__4043\ : Odrv4
    port map (
            O => \N__27422\,
            I => \sCounterRAMZ0Z_4\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__27417\,
            I => \N__27414\
        );

    \I__4041\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27411\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__27411\,
            I => \N__27407\
        );

    \I__4039\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27404\
        );

    \I__4038\ : Span4Mux_h
    port map (
            O => \N__27407\,
            I => \N__27401\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__27404\,
            I => \sCounterRAMZ0Z_7\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__27401\,
            I => \sCounterRAMZ0Z_7\
        );

    \I__4035\ : InMux
    port map (
            O => \N__27396\,
            I => \N__27393\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__27393\,
            I => \N__27389\
        );

    \I__4033\ : InMux
    port map (
            O => \N__27392\,
            I => \N__27386\
        );

    \I__4032\ : Span4Mux_v
    port map (
            O => \N__27389\,
            I => \N__27383\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__27386\,
            I => \sCounterRAMZ0Z_0\
        );

    \I__4030\ : Odrv4
    port map (
            O => \N__27383\,
            I => \sCounterRAMZ0Z_0\
        );

    \I__4029\ : InMux
    port map (
            O => \N__27378\,
            I => \N__27375\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__27375\,
            I => \N__27372\
        );

    \I__4027\ : Span12Mux_s10_v
    port map (
            O => \N__27372\,
            I => \N__27369\
        );

    \I__4026\ : Odrv12
    port map (
            O => \N__27369\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_5\
        );

    \I__4025\ : InMux
    port map (
            O => \N__27366\,
            I => \N__27363\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__27363\,
            I => \N__27360\
        );

    \I__4023\ : Odrv12
    port map (
            O => \N__27360\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_6\
        );

    \I__4022\ : InMux
    port map (
            O => \N__27357\,
            I => \N__27354\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__27354\,
            I => \N__27351\
        );

    \I__4020\ : Odrv12
    port map (
            O => \N__27351\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_7\
        );

    \I__4019\ : CEMux
    port map (
            O => \N__27348\,
            I => \N__27345\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__27345\,
            I => \spi_slave_inst.un4_i_wr\
        );

    \I__4017\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27336\
        );

    \I__4016\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27336\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__27336\,
            I => \spi_mosi_ready64_prevZ0Z2\
        );

    \I__4014\ : InMux
    port map (
            O => \N__27333\,
            I => \N__27327\
        );

    \I__4013\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27327\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__27327\,
            I => \spi_mosi_ready64_prevZ0\
        );

    \I__4011\ : CascadeMux
    port map (
            O => \N__27324\,
            I => \N__27321\
        );

    \I__4010\ : InMux
    port map (
            O => \N__27321\,
            I => \N__27318\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__27318\,
            I => \spi_mosi_ready64_prevZ0Z3\
        );

    \I__4008\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27306\
        );

    \I__4007\ : InMux
    port map (
            O => \N__27314\,
            I => \N__27306\
        );

    \I__4006\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27303\
        );

    \I__4005\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27298\
        );

    \I__4004\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27298\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__27306\,
            I => spi_mosi_ready
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__27303\,
            I => spi_mosi_ready
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__27298\,
            I => spi_mosi_ready
        );

    \I__4000\ : CascadeMux
    port map (
            O => \N__27291\,
            I => \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_\
        );

    \I__3999\ : IoInMux
    port map (
            O => \N__27288\,
            I => \N__27285\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__27285\,
            I => \N__27282\
        );

    \I__3997\ : Span12Mux_s3_v
    port map (
            O => \N__27282\,
            I => \N__27279\
        );

    \I__3996\ : Span12Mux_v
    port map (
            O => \N__27279\,
            I => \N__27276\
        );

    \I__3995\ : Odrv12
    port map (
            O => \N__27276\,
            I => \LED3_c_i\
        );

    \I__3994\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27270\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__27270\,
            I => \N__27267\
        );

    \I__3992\ : Odrv12
    port map (
            O => \N__27267\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_0\
        );

    \I__3991\ : InMux
    port map (
            O => \N__27264\,
            I => \N__27261\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__27261\,
            I => \N__27258\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__27258\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_1\
        );

    \I__3988\ : InMux
    port map (
            O => \N__27255\,
            I => \N__27252\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__27252\,
            I => \N__27249\
        );

    \I__3986\ : Odrv4
    port map (
            O => \N__27249\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_2\
        );

    \I__3985\ : InMux
    port map (
            O => \N__27246\,
            I => \N__27243\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__27243\,
            I => \N__27240\
        );

    \I__3983\ : Odrv12
    port map (
            O => \N__27240\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_3\
        );

    \I__3982\ : InMux
    port map (
            O => \N__27237\,
            I => \N__27234\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__27234\,
            I => \N__27231\
        );

    \I__3980\ : Span4Mux_h
    port map (
            O => \N__27231\,
            I => \N__27228\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__27228\,
            I => \N__27225\
        );

    \I__3978\ : Odrv4
    port map (
            O => \N__27225\,
            I => \spi_slave_inst.data_in_reg_iZ0Z_4\
        );

    \I__3977\ : CascadeMux
    port map (
            O => \N__27222\,
            I => \N_206_cascade_\
        );

    \I__3976\ : CEMux
    port map (
            O => \N__27219\,
            I => \N__27216\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__27216\,
            I => \N__27213\
        );

    \I__3974\ : Span4Mux_v
    port map (
            O => \N__27213\,
            I => \N__27210\
        );

    \I__3973\ : Span4Mux_v
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__3972\ : Odrv4
    port map (
            O => \N__27207\,
            I => \sAddress_RNIA6242_1Z0Z_0\
        );

    \I__3971\ : InMux
    port map (
            O => \N__27204\,
            I => \N__27201\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__27201\,
            I => \N__27198\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__27198\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_3\
        );

    \I__3968\ : InMux
    port map (
            O => \N__27195\,
            I => \N__27192\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__27192\,
            I => \N__27189\
        );

    \I__3966\ : Odrv4
    port map (
            O => \N__27189\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_7\
        );

    \I__3965\ : InMux
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__27183\,
            I => \N__27180\
        );

    \I__3963\ : Odrv12
    port map (
            O => \N__27180\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_5\
        );

    \I__3962\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27174\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__27174\,
            I => \N__27171\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__27171\,
            I => \spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1\
        );

    \I__3959\ : InMux
    port map (
            O => \N__27168\,
            I => \N__27165\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__27165\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_1\
        );

    \I__3957\ : InMux
    port map (
            O => \N__27162\,
            I => \N__27159\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__27159\,
            I => \N__27156\
        );

    \I__3955\ : Odrv4
    port map (
            O => \N__27156\,
            I => \spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2\
        );

    \I__3954\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27150\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__27150\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_2\
        );

    \I__3952\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27144\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__27144\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_6\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__27141\,
            I => \N__27138\
        );

    \I__3949\ : InMux
    port map (
            O => \N__27138\,
            I => \N__27135\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__27135\,
            I => \N__27132\
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__27132\,
            I => \N_206\
        );

    \I__3946\ : CascadeMux
    port map (
            O => \N__27129\,
            I => \spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3_cascade_\
        );

    \I__3945\ : InMux
    port map (
            O => \N__27126\,
            I => \N__27123\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__27123\,
            I => \spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0\
        );

    \I__3943\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27117\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__27117\,
            I => \spi_slave_inst.N_1394\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__27114\,
            I => \spi_slave_inst.N_1397_cascade_\
        );

    \I__3940\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27108\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__27108\,
            I => \spi_slave_inst.tx_done_reg1_iZ0\
        );

    \I__3938\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27101\
        );

    \I__3937\ : InMux
    port map (
            O => \N__27104\,
            I => \N__27098\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__27101\,
            I => \N__27095\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__27098\,
            I => \spi_slave_inst.tx_done_reg2_iZ0\
        );

    \I__3934\ : Odrv4
    port map (
            O => \N__27095\,
            I => \spi_slave_inst.tx_done_reg2_iZ0\
        );

    \I__3933\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27087\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__27087\,
            I => \N__27084\
        );

    \I__3931\ : Span4Mux_v
    port map (
            O => \N__27084\,
            I => \N__27081\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__27081\,
            I => \spi_slave_inst.tx_done_reg3_iZ0\
        );

    \I__3929\ : InMux
    port map (
            O => \N__27078\,
            I => \N__27075\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__27075\,
            I => \N__27072\
        );

    \I__3927\ : Span4Mux_v
    port map (
            O => \N__27072\,
            I => \N__27069\
        );

    \I__3926\ : Odrv4
    port map (
            O => \N__27069\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_0\
        );

    \I__3925\ : InMux
    port map (
            O => \N__27066\,
            I => \N__27062\
        );

    \I__3924\ : InMux
    port map (
            O => \N__27065\,
            I => \N__27059\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__27062\,
            I => \spi_slave_inst.rx_done_neg_sclk_iZ0\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__27059\,
            I => \spi_slave_inst.rx_done_neg_sclk_iZ0\
        );

    \I__3921\ : InMux
    port map (
            O => \N__27054\,
            I => \N__27051\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__27051\,
            I => \spi_slave_inst.rx_done_pos_sclk_iZ0\
        );

    \I__3919\ : InMux
    port map (
            O => \N__27048\,
            I => \N__27045\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__27045\,
            I => \spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0\
        );

    \I__3917\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27036\
        );

    \I__3916\ : InMux
    port map (
            O => \N__27041\,
            I => \N__27036\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__27036\,
            I => \spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0\
        );

    \I__3914\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27030\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__27030\,
            I => \N__27027\
        );

    \I__3912\ : Span4Mux_v
    port map (
            O => \N__27027\,
            I => \N__27023\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__27026\,
            I => \N__27020\
        );

    \I__3910\ : Sp12to4
    port map (
            O => \N__27023\,
            I => \N__27017\
        );

    \I__3909\ : InMux
    port map (
            O => \N__27020\,
            I => \N__27014\
        );

    \I__3908\ : Odrv12
    port map (
            O => \N__27017\,
            I => \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__27014\,
            I => \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0\
        );

    \I__3906\ : InMux
    port map (
            O => \N__27009\,
            I => \N__27006\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__27006\,
            I => \spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0\
        );

    \I__3904\ : InMux
    port map (
            O => \N__27003\,
            I => \N__26995\
        );

    \I__3903\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26995\
        );

    \I__3902\ : InMux
    port map (
            O => \N__27001\,
            I => \N__26989\
        );

    \I__3901\ : InMux
    port map (
            O => \N__27000\,
            I => \N__26989\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__26995\,
            I => \N__26986\
        );

    \I__3899\ : InMux
    port map (
            O => \N__26994\,
            I => \N__26983\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__26989\,
            I => \N__26980\
        );

    \I__3897\ : Span4Mux_v
    port map (
            O => \N__26986\,
            I => \N__26977\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__26983\,
            I => \N__26974\
        );

    \I__3895\ : Span4Mux_v
    port map (
            O => \N__26980\,
            I => \N__26971\
        );

    \I__3894\ : Span4Mux_h
    port map (
            O => \N__26977\,
            I => \N__26966\
        );

    \I__3893\ : Span4Mux_v
    port map (
            O => \N__26974\,
            I => \N__26966\
        );

    \I__3892\ : Span4Mux_h
    port map (
            O => \N__26971\,
            I => \N__26963\
        );

    \I__3891\ : Odrv4
    port map (
            O => \N__26966\,
            I => \spi_master_inst.sclk_gen_u0.spi_start_iZ0\
        );

    \I__3890\ : Odrv4
    port map (
            O => \N__26963\,
            I => \spi_master_inst.sclk_gen_u0.spi_start_iZ0\
        );

    \I__3889\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26955\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__26955\,
            I => \spi_slave_inst.txdata_reg_iZ0Z_4\
        );

    \I__3887\ : InMux
    port map (
            O => \N__26952\,
            I => \N__26949\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__26949\,
            I => \sEEDelayACQZ0Z_9\
        );

    \I__3885\ : CEMux
    port map (
            O => \N__26946\,
            I => \N__26943\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__26943\,
            I => \N__26940\
        );

    \I__3883\ : Span4Mux_v
    port map (
            O => \N__26940\,
            I => \N__26937\
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__26937\,
            I => \sAddress_RNIA6242Z0Z_0\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__26934\,
            I => \N_99_cascade_\
        );

    \I__3880\ : IoInMux
    port map (
            O => \N__26931\,
            I => \N__26928\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__26928\,
            I => \N__26925\
        );

    \I__3878\ : Span4Mux_s2_v
    port map (
            O => \N__26925\,
            I => \N__26922\
        );

    \I__3877\ : Span4Mux_h
    port map (
            O => \N__26922\,
            I => \N__26919\
        );

    \I__3876\ : Span4Mux_h
    port map (
            O => \N__26919\,
            I => \N__26916\
        );

    \I__3875\ : Span4Mux_h
    port map (
            O => \N__26916\,
            I => \N__26913\
        );

    \I__3874\ : Span4Mux_v
    port map (
            O => \N__26913\,
            I => \N__26909\
        );

    \I__3873\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26906\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__26909\,
            I => \RAM_DATA_cl_12Z0Z_15\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__26906\,
            I => \RAM_DATA_cl_12Z0Z_15\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__26901\,
            I => \N_94_cascade_\
        );

    \I__3869\ : IoInMux
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__26895\,
            I => \N__26892\
        );

    \I__3867\ : IoSpan4Mux
    port map (
            O => \N__26892\,
            I => \N__26889\
        );

    \I__3866\ : Span4Mux_s2_h
    port map (
            O => \N__26889\,
            I => \N__26886\
        );

    \I__3865\ : Sp12to4
    port map (
            O => \N__26886\,
            I => \N__26883\
        );

    \I__3864\ : Span12Mux_v
    port map (
            O => \N__26883\,
            I => \N__26880\
        );

    \I__3863\ : Span12Mux_h
    port map (
            O => \N__26880\,
            I => \N__26876\
        );

    \I__3862\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26873\
        );

    \I__3861\ : Odrv12
    port map (
            O => \N__26876\,
            I => \RAM_DATA_cl_11Z0Z_15\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__26873\,
            I => \RAM_DATA_cl_11Z0Z_15\
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__26868\,
            I => \N_104_cascade_\
        );

    \I__3858\ : IoInMux
    port map (
            O => \N__26865\,
            I => \N__26862\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__26862\,
            I => \N__26859\
        );

    \I__3856\ : Span4Mux_s0_v
    port map (
            O => \N__26859\,
            I => \N__26856\
        );

    \I__3855\ : Sp12to4
    port map (
            O => \N__26856\,
            I => \N__26853\
        );

    \I__3854\ : Span12Mux_h
    port map (
            O => \N__26853\,
            I => \N__26849\
        );

    \I__3853\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26846\
        );

    \I__3852\ : Odrv12
    port map (
            O => \N__26849\,
            I => \RAM_DATA_cl_14Z0Z_15\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__26846\,
            I => \RAM_DATA_cl_14Z0Z_15\
        );

    \I__3850\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26838\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__26838\,
            I => \N__26835\
        );

    \I__3848\ : Span4Mux_v
    port map (
            O => \N__26835\,
            I => \N__26832\
        );

    \I__3847\ : Odrv4
    port map (
            O => \N__26832\,
            I => \sDAC_dataZ0Z_2\
        );

    \I__3846\ : InMux
    port map (
            O => \N__26829\,
            I => \N__26823\
        );

    \I__3845\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26820\
        );

    \I__3844\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26815\
        );

    \I__3843\ : InMux
    port map (
            O => \N__26826\,
            I => \N__26815\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__26823\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_i6\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__26820\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_i6\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__26815\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_i6\
        );

    \I__3839\ : InMux
    port map (
            O => \N__26808\,
            I => \N__26805\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__26805\,
            I => \sEEDelayACQZ0Z_6\
        );

    \I__3837\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26799\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__26799\,
            I => \sEEDelayACQZ0Z_7\
        );

    \I__3835\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26793\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__26793\,
            I => \sEEDelayACQZ0Z_10\
        );

    \I__3833\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26787\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__26787\,
            I => \sEEDelayACQZ0Z_11\
        );

    \I__3831\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26781\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__26781\,
            I => \sEEDelayACQZ0Z_12\
        );

    \I__3829\ : InMux
    port map (
            O => \N__26778\,
            I => \N__26775\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__26775\,
            I => \sEEDelayACQZ0Z_13\
        );

    \I__3827\ : InMux
    port map (
            O => \N__26772\,
            I => \N__26769\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__26769\,
            I => \sEEDelayACQZ0Z_14\
        );

    \I__3825\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26763\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__26763\,
            I => \sEEDelayACQZ0Z_15\
        );

    \I__3823\ : InMux
    port map (
            O => \N__26760\,
            I => \N__26757\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__26757\,
            I => \sEEDelayACQZ0Z_8\
        );

    \I__3821\ : CEMux
    port map (
            O => \N__26754\,
            I => \N__26751\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__26751\,
            I => \N__26748\
        );

    \I__3819\ : Span4Mux_v
    port map (
            O => \N__26748\,
            I => \N__26745\
        );

    \I__3818\ : Odrv4
    port map (
            O => \N__26745\,
            I => \N_76_i\
        );

    \I__3817\ : CascadeMux
    port map (
            O => \N__26742\,
            I => \N_71_cascade_\
        );

    \I__3816\ : InMux
    port map (
            O => \N__26739\,
            I => \N__26736\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__26736\,
            I => \sEEDelayACQZ0Z_0\
        );

    \I__3814\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26730\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__26730\,
            I => \sEEDelayACQZ0Z_1\
        );

    \I__3812\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26724\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__26724\,
            I => \sEEDelayACQZ0Z_2\
        );

    \I__3810\ : InMux
    port map (
            O => \N__26721\,
            I => \N__26718\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__26718\,
            I => \sEEDelayACQZ0Z_3\
        );

    \I__3808\ : InMux
    port map (
            O => \N__26715\,
            I => \N__26712\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__26712\,
            I => \sEEDelayACQZ0Z_4\
        );

    \I__3806\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26706\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__26706\,
            I => \sEEDelayACQZ0Z_5\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__26703\,
            I => \N__26700\
        );

    \I__3803\ : InMux
    port map (
            O => \N__26700\,
            I => \N__26697\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__26697\,
            I => un1_sacqtime_cry_18_sf
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__26694\,
            I => \N__26691\
        );

    \I__3800\ : InMux
    port map (
            O => \N__26691\,
            I => \N__26688\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__26688\,
            I => un1_sacqtime_cry_19_sf
        );

    \I__3798\ : CascadeMux
    port map (
            O => \N__26685\,
            I => \N__26682\
        );

    \I__3797\ : InMux
    port map (
            O => \N__26682\,
            I => \N__26679\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__26679\,
            I => un1_sacqtime_cry_20_sf
        );

    \I__3795\ : CascadeMux
    port map (
            O => \N__26676\,
            I => \N__26673\
        );

    \I__3794\ : InMux
    port map (
            O => \N__26673\,
            I => \N__26670\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__26670\,
            I => un1_sacqtime_cry_21_sf
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__26667\,
            I => \N__26664\
        );

    \I__3791\ : InMux
    port map (
            O => \N__26664\,
            I => \N__26661\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__26661\,
            I => un1_sacqtime_cry_22_sf
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__26658\,
            I => \N__26655\
        );

    \I__3788\ : InMux
    port map (
            O => \N__26655\,
            I => \N__26652\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__26652\,
            I => un1_sacqtime_cry_23_sf
        );

    \I__3786\ : InMux
    port map (
            O => \N__26649\,
            I => \bfn_10_17_0_\
        );

    \I__3785\ : IoInMux
    port map (
            O => \N__26646\,
            I => \N__26643\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__26643\,
            I => \N__26640\
        );

    \I__3783\ : IoSpan4Mux
    port map (
            O => \N__26640\,
            I => \N__26637\
        );

    \I__3782\ : Span4Mux_s2_h
    port map (
            O => \N__26637\,
            I => \N__26634\
        );

    \I__3781\ : Sp12to4
    port map (
            O => \N__26634\,
            I => \N__26631\
        );

    \I__3780\ : Span12Mux_s9_h
    port map (
            O => \N__26631\,
            I => \N__26628\
        );

    \I__3779\ : Span12Mux_h
    port map (
            O => \N__26628\,
            I => \N__26624\
        );

    \I__3778\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26621\
        );

    \I__3777\ : Span12Mux_v
    port map (
            O => \N__26624\,
            I => \N__26618\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__26621\,
            I => \N__26615\
        );

    \I__3775\ : Odrv12
    port map (
            O => \N__26618\,
            I => \RAM_DATA_cl_10Z0Z_15\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__26615\,
            I => \RAM_DATA_cl_10Z0Z_15\
        );

    \I__3773\ : InMux
    port map (
            O => \N__26610\,
            I => \N__26607\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__26607\,
            I => \N__26604\
        );

    \I__3771\ : Odrv12
    port map (
            O => \N__26604\,
            I => \N_106\
        );

    \I__3770\ : IoInMux
    port map (
            O => \N__26601\,
            I => \N__26598\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__26598\,
            I => \N__26595\
        );

    \I__3768\ : IoSpan4Mux
    port map (
            O => \N__26595\,
            I => \N__26592\
        );

    \I__3767\ : Span4Mux_s2_v
    port map (
            O => \N__26592\,
            I => \N__26589\
        );

    \I__3766\ : Span4Mux_v
    port map (
            O => \N__26589\,
            I => \N__26586\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__26586\,
            I => \N_26\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__26583\,
            I => \N__26579\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__26582\,
            I => \N__26576\
        );

    \I__3762\ : InMux
    port map (
            O => \N__26579\,
            I => \N__26573\
        );

    \I__3761\ : InMux
    port map (
            O => \N__26576\,
            I => \N__26570\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__26573\,
            I => \sCounter_i_10\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__26570\,
            I => \sCounter_i_10\
        );

    \I__3758\ : CascadeMux
    port map (
            O => \N__26565\,
            I => \N__26561\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__26564\,
            I => \N__26558\
        );

    \I__3756\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26555\
        );

    \I__3755\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26552\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__26555\,
            I => \sCounter_i_11\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__26552\,
            I => \sCounter_i_11\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__26547\,
            I => \N__26543\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__26546\,
            I => \N__26540\
        );

    \I__3750\ : InMux
    port map (
            O => \N__26543\,
            I => \N__26537\
        );

    \I__3749\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26534\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__26537\,
            I => \sCounter_i_12\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__26534\,
            I => \sCounter_i_12\
        );

    \I__3746\ : CascadeMux
    port map (
            O => \N__26529\,
            I => \N__26525\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__26528\,
            I => \N__26522\
        );

    \I__3744\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26519\
        );

    \I__3743\ : InMux
    port map (
            O => \N__26522\,
            I => \N__26516\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__26519\,
            I => \sCounter_i_13\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__26516\,
            I => \sCounter_i_13\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__26511\,
            I => \N__26507\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__26510\,
            I => \N__26504\
        );

    \I__3738\ : InMux
    port map (
            O => \N__26507\,
            I => \N__26501\
        );

    \I__3737\ : InMux
    port map (
            O => \N__26504\,
            I => \N__26498\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__26501\,
            I => \sCounter_i_14\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__26498\,
            I => \sCounter_i_14\
        );

    \I__3734\ : CascadeMux
    port map (
            O => \N__26493\,
            I => \N__26489\
        );

    \I__3733\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26486\
        );

    \I__3732\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26483\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__26486\,
            I => \sCounter_i_15\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__26483\,
            I => \sCounter_i_15\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__26478\,
            I => \N__26475\
        );

    \I__3728\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26472\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__26472\,
            I => un1_sacqtime_cry_16_sf
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__26469\,
            I => \N__26466\
        );

    \I__3725\ : InMux
    port map (
            O => \N__26466\,
            I => \N__26463\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__26463\,
            I => un1_sacqtime_cry_17_sf
        );

    \I__3723\ : CascadeMux
    port map (
            O => \N__26460\,
            I => \N__26456\
        );

    \I__3722\ : CascadeMux
    port map (
            O => \N__26459\,
            I => \N__26453\
        );

    \I__3721\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26450\
        );

    \I__3720\ : InMux
    port map (
            O => \N__26453\,
            I => \N__26447\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__26450\,
            I => \sCounter_i_2\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__26447\,
            I => \sCounter_i_2\
        );

    \I__3717\ : CascadeMux
    port map (
            O => \N__26442\,
            I => \N__26438\
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__26441\,
            I => \N__26435\
        );

    \I__3715\ : InMux
    port map (
            O => \N__26438\,
            I => \N__26432\
        );

    \I__3714\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26429\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__26432\,
            I => \sCounter_i_3\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__26429\,
            I => \sCounter_i_3\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__26424\,
            I => \N__26420\
        );

    \I__3710\ : CascadeMux
    port map (
            O => \N__26423\,
            I => \N__26417\
        );

    \I__3709\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26414\
        );

    \I__3708\ : InMux
    port map (
            O => \N__26417\,
            I => \N__26411\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__26414\,
            I => \sCounter_i_4\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__26411\,
            I => \sCounter_i_4\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__26406\,
            I => \N__26402\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__26405\,
            I => \N__26399\
        );

    \I__3703\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26396\
        );

    \I__3702\ : InMux
    port map (
            O => \N__26399\,
            I => \N__26393\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__26396\,
            I => \sCounter_i_5\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__26393\,
            I => \sCounter_i_5\
        );

    \I__3699\ : CascadeMux
    port map (
            O => \N__26388\,
            I => \N__26384\
        );

    \I__3698\ : CascadeMux
    port map (
            O => \N__26387\,
            I => \N__26381\
        );

    \I__3697\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26378\
        );

    \I__3696\ : InMux
    port map (
            O => \N__26381\,
            I => \N__26375\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__26378\,
            I => \sCounter_i_6\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__26375\,
            I => \sCounter_i_6\
        );

    \I__3693\ : CascadeMux
    port map (
            O => \N__26370\,
            I => \N__26367\
        );

    \I__3692\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26363\
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__26366\,
            I => \N__26360\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__26363\,
            I => \N__26357\
        );

    \I__3689\ : InMux
    port map (
            O => \N__26360\,
            I => \N__26354\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__26357\,
            I => \sCounter_i_7\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__26354\,
            I => \sCounter_i_7\
        );

    \I__3686\ : CascadeMux
    port map (
            O => \N__26349\,
            I => \N__26345\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__26348\,
            I => \N__26342\
        );

    \I__3684\ : InMux
    port map (
            O => \N__26345\,
            I => \N__26339\
        );

    \I__3683\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26336\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__26339\,
            I => \sCounter_i_8\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__26336\,
            I => \sCounter_i_8\
        );

    \I__3680\ : CascadeMux
    port map (
            O => \N__26331\,
            I => \N__26327\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__26330\,
            I => \N__26324\
        );

    \I__3678\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26321\
        );

    \I__3677\ : InMux
    port map (
            O => \N__26324\,
            I => \N__26318\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__26321\,
            I => \sCounter_i_9\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__26318\,
            I => \sCounter_i_9\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__26313\,
            I => \N__26310\
        );

    \I__3673\ : InMux
    port map (
            O => \N__26310\,
            I => \N__26306\
        );

    \I__3672\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26303\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__26306\,
            I => \N__26300\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__26303\,
            I => \N__26295\
        );

    \I__3669\ : Span4Mux_h
    port map (
            O => \N__26300\,
            I => \N__26292\
        );

    \I__3668\ : InMux
    port map (
            O => \N__26299\,
            I => \N__26287\
        );

    \I__3667\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26287\
        );

    \I__3666\ : Sp12to4
    port map (
            O => \N__26295\,
            I => \N__26284\
        );

    \I__3665\ : Span4Mux_v
    port map (
            O => \N__26292\,
            I => \N__26281\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__26287\,
            I => \button_debounce_counterZ0Z_0\
        );

    \I__3663\ : Odrv12
    port map (
            O => \N__26284\,
            I => \button_debounce_counterZ0Z_0\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__26281\,
            I => \button_debounce_counterZ0Z_0\
        );

    \I__3661\ : InMux
    port map (
            O => \N__26274\,
            I => \N__26271\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__26271\,
            I => \N__26268\
        );

    \I__3659\ : Span4Mux_v
    port map (
            O => \N__26268\,
            I => \N__26264\
        );

    \I__3658\ : InMux
    port map (
            O => \N__26267\,
            I => \N__26261\
        );

    \I__3657\ : Span4Mux_v
    port map (
            O => \N__26264\,
            I => \N__26258\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__26261\,
            I => \N__26253\
        );

    \I__3655\ : Span4Mux_h
    port map (
            O => \N__26258\,
            I => \N__26253\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__26253\,
            I => \button_debounce_counterZ0Z_1\
        );

    \I__3653\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26247\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__26247\,
            I => \N__26244\
        );

    \I__3651\ : Glb2LocalMux
    port map (
            O => \N__26244\,
            I => \N__26226\
        );

    \I__3650\ : SRMux
    port map (
            O => \N__26243\,
            I => \N__26226\
        );

    \I__3649\ : SRMux
    port map (
            O => \N__26242\,
            I => \N__26226\
        );

    \I__3648\ : SRMux
    port map (
            O => \N__26241\,
            I => \N__26226\
        );

    \I__3647\ : SRMux
    port map (
            O => \N__26240\,
            I => \N__26226\
        );

    \I__3646\ : SRMux
    port map (
            O => \N__26239\,
            I => \N__26226\
        );

    \I__3645\ : GlobalMux
    port map (
            O => \N__26226\,
            I => \N__26223\
        );

    \I__3644\ : gio2CtrlBuf
    port map (
            O => \N__26223\,
            I => \N_3089_g\
        );

    \I__3643\ : InMux
    port map (
            O => \N__26220\,
            I => \N__26216\
        );

    \I__3642\ : InMux
    port map (
            O => \N__26219\,
            I => \N__26213\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__26216\,
            I => \spi_mosi_ready_prevZ0Z2\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__26213\,
            I => \spi_mosi_ready_prevZ0Z2\
        );

    \I__3639\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26204\
        );

    \I__3638\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26201\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__26204\,
            I => \spi_mosi_ready_prevZ0\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__26201\,
            I => \spi_mosi_ready_prevZ0\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__26196\,
            I => \N__26193\
        );

    \I__3634\ : InMux
    port map (
            O => \N__26193\,
            I => \N__26190\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__26190\,
            I => \spi_mosi_ready_prevZ0Z3\
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__26187\,
            I => \spi_mosi_ready_prev3_RNILKERZ0_cascade_\
        );

    \I__3631\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26180\
        );

    \I__3630\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26177\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__26180\,
            I => \N__26174\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__26177\,
            I => \spi_slave_inst.tx_ready_iZ0\
        );

    \I__3627\ : Odrv4
    port map (
            O => \N__26174\,
            I => \spi_slave_inst.tx_ready_iZ0\
        );

    \I__3626\ : CascadeMux
    port map (
            O => \N__26169\,
            I => \N__26165\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__26168\,
            I => \N__26162\
        );

    \I__3624\ : InMux
    port map (
            O => \N__26165\,
            I => \N__26159\
        );

    \I__3623\ : InMux
    port map (
            O => \N__26162\,
            I => \N__26156\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__26159\,
            I => \sCounter_i_0\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__26156\,
            I => \sCounter_i_0\
        );

    \I__3620\ : InMux
    port map (
            O => \N__26151\,
            I => \N__26147\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__26150\,
            I => \N__26144\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__26147\,
            I => \N__26141\
        );

    \I__3617\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26138\
        );

    \I__3616\ : Odrv4
    port map (
            O => \N__26141\,
            I => \sCounter_i_1\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__26138\,
            I => \sCounter_i_1\
        );

    \I__3614\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26130\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__26130\,
            I => \spi_slave_inst.rx_done_reg3_iZ0\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__26127\,
            I => \spi_slave_inst.rx_ready_i_RNOZ0Z_0_cascade_\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__26124\,
            I => \spi_slave_inst.un4_tx_done_reg2_i_cascade_\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__26121\,
            I => \N__26117\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__26120\,
            I => \N__26112\
        );

    \I__3608\ : InMux
    port map (
            O => \N__26117\,
            I => \N__26108\
        );

    \I__3607\ : InMux
    port map (
            O => \N__26116\,
            I => \N__26099\
        );

    \I__3606\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26099\
        );

    \I__3605\ : InMux
    port map (
            O => \N__26112\,
            I => \N__26099\
        );

    \I__3604\ : InMux
    port map (
            O => \N__26111\,
            I => \N__26099\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__26108\,
            I => \sEETrigCounterZ0Z_3\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__26099\,
            I => \sEETrigCounterZ0Z_3\
        );

    \I__3601\ : CascadeMux
    port map (
            O => \N__26094\,
            I => \N__26091\
        );

    \I__3600\ : InMux
    port map (
            O => \N__26091\,
            I => \N__26088\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__26088\,
            I => \N__26085\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__26085\,
            I => un10_trig_prev_3
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__26082\,
            I => \N__26077\
        );

    \I__3596\ : InMux
    port map (
            O => \N__26081\,
            I => \N__26071\
        );

    \I__3595\ : InMux
    port map (
            O => \N__26080\,
            I => \N__26071\
        );

    \I__3594\ : InMux
    port map (
            O => \N__26077\,
            I => \N__26066\
        );

    \I__3593\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26066\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__26071\,
            I => \sEETrigCounterZ0Z_2\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__26066\,
            I => \sEETrigCounterZ0Z_2\
        );

    \I__3590\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26058\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__26058\,
            I => un10_trig_prev_2
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__26055\,
            I => \N__26052\
        );

    \I__3587\ : InMux
    port map (
            O => \N__26052\,
            I => \N__26049\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__26049\,
            I => \N__26046\
        );

    \I__3585\ : Odrv4
    port map (
            O => \N__26046\,
            I => un10_trig_prev_0
        );

    \I__3584\ : CascadeMux
    port map (
            O => \N__26043\,
            I => \N__26039\
        );

    \I__3583\ : InMux
    port map (
            O => \N__26042\,
            I => \N__26026\
        );

    \I__3582\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26026\
        );

    \I__3581\ : InMux
    port map (
            O => \N__26038\,
            I => \N__26026\
        );

    \I__3580\ : InMux
    port map (
            O => \N__26037\,
            I => \N__26026\
        );

    \I__3579\ : InMux
    port map (
            O => \N__26036\,
            I => \N__26021\
        );

    \I__3578\ : InMux
    port map (
            O => \N__26035\,
            I => \N__26021\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__26026\,
            I => \sEETrigCounterZ0Z_0\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__26021\,
            I => \sEETrigCounterZ0Z_0\
        );

    \I__3575\ : InMux
    port map (
            O => \N__26016\,
            I => \N__26005\
        );

    \I__3574\ : InMux
    port map (
            O => \N__26015\,
            I => \N__26005\
        );

    \I__3573\ : InMux
    port map (
            O => \N__26014\,
            I => \N__26005\
        );

    \I__3572\ : InMux
    port map (
            O => \N__26013\,
            I => \N__26000\
        );

    \I__3571\ : InMux
    port map (
            O => \N__26012\,
            I => \N__26000\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__26005\,
            I => \sEETrigCounterZ0Z_1\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__26000\,
            I => \sEETrigCounterZ0Z_1\
        );

    \I__3568\ : CascadeMux
    port map (
            O => \N__25995\,
            I => \N__25992\
        );

    \I__3567\ : InMux
    port map (
            O => \N__25992\,
            I => \N__25989\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__25989\,
            I => un10_trig_prev_1
        );

    \I__3565\ : InMux
    port map (
            O => \N__25986\,
            I => \N__25983\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__25983\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_15\
        );

    \I__3563\ : InMux
    port map (
            O => \N__25980\,
            I => \N__25976\
        );

    \I__3562\ : InMux
    port map (
            O => \N__25979\,
            I => \N__25973\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__25976\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__25973\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0\
        );

    \I__3559\ : InMux
    port map (
            O => \N__25968\,
            I => \bfn_10_6_0_\
        );

    \I__3558\ : InMux
    port map (
            O => \N__25965\,
            I => \N__25961\
        );

    \I__3557\ : InMux
    port map (
            O => \N__25964\,
            I => \N__25958\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__25961\,
            I => \N__25953\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__25958\,
            I => \N__25953\
        );

    \I__3554\ : Odrv4
    port map (
            O => \N__25953\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1\
        );

    \I__3553\ : InMux
    port map (
            O => \N__25950\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0\
        );

    \I__3552\ : CascadeMux
    port map (
            O => \N__25947\,
            I => \N__25943\
        );

    \I__3551\ : InMux
    port map (
            O => \N__25946\,
            I => \N__25940\
        );

    \I__3550\ : InMux
    port map (
            O => \N__25943\,
            I => \N__25937\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__25940\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__25937\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2\
        );

    \I__3547\ : InMux
    port map (
            O => \N__25932\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1\
        );

    \I__3546\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25925\
        );

    \I__3545\ : InMux
    port map (
            O => \N__25928\,
            I => \N__25922\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__25925\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__25922\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3\
        );

    \I__3542\ : InMux
    port map (
            O => \N__25917\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2\
        );

    \I__3541\ : InMux
    port map (
            O => \N__25914\,
            I => \N__25910\
        );

    \I__3540\ : InMux
    port map (
            O => \N__25913\,
            I => \N__25907\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__25910\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__25907\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4\
        );

    \I__3537\ : InMux
    port map (
            O => \N__25902\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3\
        );

    \I__3536\ : InMux
    port map (
            O => \N__25899\,
            I => \N__25895\
        );

    \I__3535\ : InMux
    port map (
            O => \N__25898\,
            I => \N__25892\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__25895\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__25892\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5\
        );

    \I__3532\ : InMux
    port map (
            O => \N__25887\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4\
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__25884\,
            I => \N__25880\
        );

    \I__3530\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25877\
        );

    \I__3529\ : InMux
    port map (
            O => \N__25880\,
            I => \N__25874\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__25877\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__25874\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6\
        );

    \I__3526\ : InMux
    port map (
            O => \N__25869\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5\
        );

    \I__3525\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25848\
        );

    \I__3524\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25848\
        );

    \I__3523\ : InMux
    port map (
            O => \N__25864\,
            I => \N__25848\
        );

    \I__3522\ : InMux
    port map (
            O => \N__25863\,
            I => \N__25848\
        );

    \I__3521\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25848\
        );

    \I__3520\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25841\
        );

    \I__3519\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25841\
        );

    \I__3518\ : InMux
    port map (
            O => \N__25859\,
            I => \N__25841\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__25848\,
            I => \N__25836\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__25841\,
            I => \N__25836\
        );

    \I__3515\ : Odrv4
    port map (
            O => \N__25836\,
            I => \spi_master_inst.sclk_gen_u0.falling_count_start_i_i\
        );

    \I__3514\ : InMux
    port map (
            O => \N__25833\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6\
        );

    \I__3513\ : InMux
    port map (
            O => \N__25830\,
            I => \N__25826\
        );

    \I__3512\ : InMux
    port map (
            O => \N__25829\,
            I => \N__25823\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__25826\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__25823\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7\
        );

    \I__3509\ : CEMux
    port map (
            O => \N__25818\,
            I => \N__25815\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__25815\,
            I => \N__25812\
        );

    \I__3507\ : Span4Mux_h
    port map (
            O => \N__25812\,
            I => \N__25809\
        );

    \I__3506\ : Sp12to4
    port map (
            O => \N__25809\,
            I => \N__25806\
        );

    \I__3505\ : Odrv12
    port map (
            O => \N__25806\,
            I => \spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i\
        );

    \I__3504\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25800\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__25800\,
            I => \spi_slave_inst.un23_i_ssn_3\
        );

    \I__3502\ : InMux
    port map (
            O => \N__25797\,
            I => \N__25792\
        );

    \I__3501\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25789\
        );

    \I__3500\ : InMux
    port map (
            O => \N__25795\,
            I => \N__25786\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__25792\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__25789\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__25786\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5\
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__25779\,
            I => \N__25775\
        );

    \I__3495\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25770\
        );

    \I__3494\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25767\
        );

    \I__3493\ : InMux
    port map (
            O => \N__25774\,
            I => \N__25764\
        );

    \I__3492\ : InMux
    port map (
            O => \N__25773\,
            I => \N__25761\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__25770\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__25767\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__25764\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__25761\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2\
        );

    \I__3487\ : InMux
    port map (
            O => \N__25752\,
            I => \N__25749\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__25749\,
            I => \N__25746\
        );

    \I__3485\ : Span12Mux_s9_h
    port map (
            O => \N__25746\,
            I => \N__25743\
        );

    \I__3484\ : Odrv12
    port map (
            O => \N__25743\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_6\
        );

    \I__3483\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25737\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__25737\,
            I => \N__25734\
        );

    \I__3481\ : Span4Mux_v
    port map (
            O => \N__25734\,
            I => \N__25731\
        );

    \I__3480\ : Odrv4
    port map (
            O => \N__25731\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_1\
        );

    \I__3479\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25725\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__25725\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_2\
        );

    \I__3477\ : InMux
    port map (
            O => \N__25722\,
            I => \N__25719\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__25719\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_11\
        );

    \I__3475\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25713\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__25713\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_12\
        );

    \I__3473\ : InMux
    port map (
            O => \N__25710\,
            I => \N__25707\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__25707\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_3\
        );

    \I__3471\ : InMux
    port map (
            O => \N__25704\,
            I => \N__25701\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__25701\,
            I => \N__25698\
        );

    \I__3469\ : Span4Mux_h
    port map (
            O => \N__25698\,
            I => \N__25695\
        );

    \I__3468\ : Odrv4
    port map (
            O => \N__25695\,
            I => \spi_master_inst.spi_data_path_u1.data_inZ0Z_14\
        );

    \I__3467\ : InMux
    port map (
            O => \N__25692\,
            I => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3\
        );

    \I__3466\ : InMux
    port map (
            O => \N__25689\,
            I => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4\
        );

    \I__3465\ : InMux
    port map (
            O => \N__25686\,
            I => \N__25682\
        );

    \I__3464\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25679\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__25682\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__25679\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__3461\ : InMux
    port map (
            O => \N__25674\,
            I => \N__25670\
        );

    \I__3460\ : InMux
    port map (
            O => \N__25673\,
            I => \N__25667\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__25670\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__25667\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__25662\,
            I => \N__25658\
        );

    \I__3456\ : InMux
    port map (
            O => \N__25661\,
            I => \N__25655\
        );

    \I__3455\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25652\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__25655\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__25652\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__3452\ : InMux
    port map (
            O => \N__25647\,
            I => \N__25643\
        );

    \I__3451\ : InMux
    port map (
            O => \N__25646\,
            I => \N__25640\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__25643\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__25640\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__3448\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25631\
        );

    \I__3447\ : InMux
    port map (
            O => \N__25634\,
            I => \N__25628\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__25631\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__25628\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__25623\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_i6_3_cascade_\
        );

    \I__3443\ : InMux
    port map (
            O => \N__25620\,
            I => \N__25616\
        );

    \I__3442\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25613\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__25616\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__25613\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__25608\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__25605\,
            I => \N__25601\
        );

    \I__3437\ : InMux
    port map (
            O => \N__25604\,
            I => \N__25598\
        );

    \I__3436\ : InMux
    port map (
            O => \N__25601\,
            I => \N__25595\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__25598\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_5\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__25595\,
            I => \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_5\
        );

    \I__3433\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25586\
        );

    \I__3432\ : InMux
    port map (
            O => \N__25589\,
            I => \N__25583\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__25586\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__25583\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3\
        );

    \I__3429\ : CascadeMux
    port map (
            O => \N__25578\,
            I => \N__25575\
        );

    \I__3428\ : InMux
    port map (
            O => \N__25575\,
            I => \N__25570\
        );

    \I__3427\ : InMux
    port map (
            O => \N__25574\,
            I => \N__25567\
        );

    \I__3426\ : InMux
    port map (
            O => \N__25573\,
            I => \N__25564\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__25570\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__25567\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__25564\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__25557\,
            I => \N__25553\
        );

    \I__3421\ : CascadeMux
    port map (
            O => \N__25556\,
            I => \N__25549\
        );

    \I__3420\ : InMux
    port map (
            O => \N__25553\,
            I => \N__25546\
        );

    \I__3419\ : InMux
    port map (
            O => \N__25552\,
            I => \N__25543\
        );

    \I__3418\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25540\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__25546\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__25543\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__25540\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0\
        );

    \I__3414\ : InMux
    port map (
            O => \N__25533\,
            I => \N__25529\
        );

    \I__3413\ : InMux
    port map (
            O => \N__25532\,
            I => \N__25526\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__25529\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__25526\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4\
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__25521\,
            I => \spi_slave_inst.un23_i_ssn_3_cascade_\
        );

    \I__3409\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25509\
        );

    \I__3408\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25509\
        );

    \I__3407\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25509\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__25509\,
            I => \spi_slave_inst.un23_i_ssn\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__25506\,
            I => \spi_slave_inst.un23_i_ssn_cascade_\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__25503\,
            I => \N__25499\
        );

    \I__3403\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25496\
        );

    \I__3402\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25493\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__25496\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__25493\,
            I => \spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa\
        );

    \I__3399\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25485\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__25485\,
            I => \N__25482\
        );

    \I__3397\ : Span4Mux_h
    port map (
            O => \N__25482\,
            I => \N__25479\
        );

    \I__3396\ : Span4Mux_h
    port map (
            O => \N__25479\,
            I => \N__25476\
        );

    \I__3395\ : Odrv4
    port map (
            O => \N__25476\,
            I => op_gt_op_gt_un13_striginternallto23_8
        );

    \I__3394\ : InMux
    port map (
            O => \N__25473\,
            I => \bfn_9_20_0_\
        );

    \I__3393\ : CEMux
    port map (
            O => \N__25470\,
            I => \N__25467\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__25467\,
            I => \N__25464\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__25464\,
            I => \LED3_c_0\
        );

    \I__3390\ : InMux
    port map (
            O => \N__25461\,
            I => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0\
        );

    \I__3389\ : InMux
    port map (
            O => \N__25458\,
            I => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1\
        );

    \I__3388\ : InMux
    port map (
            O => \N__25455\,
            I => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__25452\,
            I => \N__25449\
        );

    \I__3386\ : InMux
    port map (
            O => \N__25449\,
            I => \N__25446\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__25446\,
            I => \sEEDelayACQ_i_12\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__25443\,
            I => \N__25440\
        );

    \I__3383\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25437\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__25437\,
            I => \sEEDelayACQ_i_13\
        );

    \I__3381\ : CascadeMux
    port map (
            O => \N__25434\,
            I => \N__25431\
        );

    \I__3380\ : InMux
    port map (
            O => \N__25431\,
            I => \N__25428\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__25428\,
            I => \sEEDelayACQ_i_14\
        );

    \I__3378\ : InMux
    port map (
            O => \N__25425\,
            I => \N__25422\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__25422\,
            I => \sEEDelayACQ_i_15\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__25419\,
            I => \N__25416\
        );

    \I__3375\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25413\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__25413\,
            I => \sEEDelayACQ_i_4\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__25410\,
            I => \N__25407\
        );

    \I__3372\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25404\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__25404\,
            I => \sEEDelayACQ_i_5\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__25401\,
            I => \N__25398\
        );

    \I__3369\ : InMux
    port map (
            O => \N__25398\,
            I => \N__25395\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__25395\,
            I => \sEEDelayACQ_i_6\
        );

    \I__3367\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25389\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__25389\,
            I => \sEEDelayACQ_i_7\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__25386\,
            I => \N__25383\
        );

    \I__3364\ : InMux
    port map (
            O => \N__25383\,
            I => \N__25380\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__25380\,
            I => \sEEDelayACQ_i_8\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__25377\,
            I => \N__25374\
        );

    \I__3361\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25371\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__25371\,
            I => \sEEDelayACQ_i_9\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__25368\,
            I => \N__25365\
        );

    \I__3358\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25362\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__25362\,
            I => \sEEDelayACQ_i_10\
        );

    \I__3356\ : CascadeMux
    port map (
            O => \N__25359\,
            I => \N__25356\
        );

    \I__3355\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25353\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__25353\,
            I => \sEEDelayACQ_i_11\
        );

    \I__3353\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25347\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__25347\,
            I => \N__25344\
        );

    \I__3351\ : Span4Mux_v
    port map (
            O => \N__25344\,
            I => \N__25341\
        );

    \I__3350\ : Odrv4
    port map (
            O => \N__25341\,
            I => \un4_spoff_cry_23_THRU_CO\
        );

    \I__3349\ : InMux
    port map (
            O => \N__25338\,
            I => \bfn_9_16_0_\
        );

    \I__3348\ : IoInMux
    port map (
            O => \N__25335\,
            I => \N__25332\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__25332\,
            I => \N__25329\
        );

    \I__3346\ : Span12Mux_s8_h
    port map (
            O => \N__25329\,
            I => \N__25326\
        );

    \I__3345\ : Odrv12
    port map (
            O => \N__25326\,
            I => \N_1612_i\
        );

    \I__3344\ : InMux
    port map (
            O => \N__25323\,
            I => \N__25319\
        );

    \I__3343\ : InMux
    port map (
            O => \N__25322\,
            I => \N__25316\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__25319\,
            I => \N__25311\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__25316\,
            I => \N__25311\
        );

    \I__3340\ : Odrv4
    port map (
            O => \N__25311\,
            I => \sCounterRAMZ0Z_6\
        );

    \I__3339\ : InMux
    port map (
            O => \N__25308\,
            I => \N__25304\
        );

    \I__3338\ : InMux
    port map (
            O => \N__25307\,
            I => \N__25301\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__25304\,
            I => \N__25298\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__25301\,
            I => \sCounterRAMZ0Z_3\
        );

    \I__3335\ : Odrv4
    port map (
            O => \N__25298\,
            I => \sCounterRAMZ0Z_3\
        );

    \I__3334\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25290\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__25290\,
            I => \N__25287\
        );

    \I__3332\ : Span4Mux_v
    port map (
            O => \N__25287\,
            I => \N__25283\
        );

    \I__3331\ : InMux
    port map (
            O => \N__25286\,
            I => \N__25280\
        );

    \I__3330\ : Odrv4
    port map (
            O => \N__25283\,
            I => \button_debounce_counterZ0Z_21\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__25280\,
            I => \button_debounce_counterZ0Z_21\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__25275\,
            I => \N__25272\
        );

    \I__3327\ : InMux
    port map (
            O => \N__25272\,
            I => \N__25269\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__25269\,
            I => \N__25266\
        );

    \I__3325\ : Span4Mux_v
    port map (
            O => \N__25266\,
            I => \N__25262\
        );

    \I__3324\ : InMux
    port map (
            O => \N__25265\,
            I => \N__25259\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__25262\,
            I => \button_debounce_counterZ0Z_22\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__25259\,
            I => \button_debounce_counterZ0Z_22\
        );

    \I__3321\ : InMux
    port map (
            O => \N__25254\,
            I => \N__25251\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__25251\,
            I => \sbuttonModeStatus_0_sqmuxa_0\
        );

    \I__3319\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25245\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__25245\,
            I => \N__25242\
        );

    \I__3317\ : Span4Mux_h
    port map (
            O => \N__25242\,
            I => \N__25239\
        );

    \I__3316\ : Odrv4
    port map (
            O => \N__25239\,
            I => \sbuttonModeStatus_0_sqmuxa_18\
        );

    \I__3315\ : InMux
    port map (
            O => \N__25236\,
            I => \N__25232\
        );

    \I__3314\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25229\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__25232\,
            I => \button_debounce_counterZ0Z_4\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__25229\,
            I => \button_debounce_counterZ0Z_4\
        );

    \I__3311\ : InMux
    port map (
            O => \N__25224\,
            I => \N__25220\
        );

    \I__3310\ : InMux
    port map (
            O => \N__25223\,
            I => \N__25217\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__25220\,
            I => \button_debounce_counterZ0Z_3\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__25217\,
            I => \button_debounce_counterZ0Z_3\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__25212\,
            I => \N__25208\
        );

    \I__3306\ : InMux
    port map (
            O => \N__25211\,
            I => \N__25205\
        );

    \I__3305\ : InMux
    port map (
            O => \N__25208\,
            I => \N__25202\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__25205\,
            I => \button_debounce_counterZ0Z_5\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__25202\,
            I => \button_debounce_counterZ0Z_5\
        );

    \I__3302\ : InMux
    port map (
            O => \N__25197\,
            I => \N__25193\
        );

    \I__3301\ : InMux
    port map (
            O => \N__25196\,
            I => \N__25190\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__25193\,
            I => \button_debounce_counterZ0Z_2\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__25190\,
            I => \button_debounce_counterZ0Z_2\
        );

    \I__3298\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25182\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__25182\,
            I => \N__25179\
        );

    \I__3296\ : Span4Mux_h
    port map (
            O => \N__25179\,
            I => \N__25176\
        );

    \I__3295\ : Odrv4
    port map (
            O => \N__25176\,
            I => \sbuttonModeStatus_0_sqmuxa_13\
        );

    \I__3294\ : CascadeMux
    port map (
            O => \N__25173\,
            I => \N__25170\
        );

    \I__3293\ : InMux
    port map (
            O => \N__25170\,
            I => \N__25167\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__25167\,
            I => \sEEDelayACQ_i_0\
        );

    \I__3291\ : CascadeMux
    port map (
            O => \N__25164\,
            I => \N__25161\
        );

    \I__3290\ : InMux
    port map (
            O => \N__25161\,
            I => \N__25158\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__25158\,
            I => \sEEDelayACQ_i_1\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__25155\,
            I => \N__25152\
        );

    \I__3287\ : InMux
    port map (
            O => \N__25152\,
            I => \N__25149\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__25149\,
            I => \sEEDelayACQ_i_2\
        );

    \I__3285\ : CascadeMux
    port map (
            O => \N__25146\,
            I => \N__25143\
        );

    \I__3284\ : InMux
    port map (
            O => \N__25143\,
            I => \N__25140\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__25140\,
            I => \sEEDelayACQ_i_3\
        );

    \I__3282\ : InMux
    port map (
            O => \N__25137\,
            I => \N__25134\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__25134\,
            I => \sCounter_i_16\
        );

    \I__3280\ : InMux
    port map (
            O => \N__25131\,
            I => \N__25128\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__25128\,
            I => \sCounter_i_17\
        );

    \I__3278\ : InMux
    port map (
            O => \N__25125\,
            I => \N__25122\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__25122\,
            I => \sCounter_i_18\
        );

    \I__3276\ : InMux
    port map (
            O => \N__25119\,
            I => \N__25116\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__25116\,
            I => \sCounter_i_19\
        );

    \I__3274\ : InMux
    port map (
            O => \N__25113\,
            I => \N__25110\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__25110\,
            I => \sCounter_i_20\
        );

    \I__3272\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25104\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__25104\,
            I => \sCounter_i_21\
        );

    \I__3270\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25098\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__25098\,
            I => \sCounter_i_22\
        );

    \I__3268\ : InMux
    port map (
            O => \N__25095\,
            I => \N__25092\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__25092\,
            I => \sCounter_i_23\
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__25089\,
            I => \un1_reset_rpi_inv_2_i_1_cascade_\
        );

    \I__3265\ : InMux
    port map (
            O => \N__25086\,
            I => \N__25083\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__25083\,
            I => \N__25080\
        );

    \I__3263\ : Odrv4
    port map (
            O => \N__25080\,
            I => \un1_sTrigCounter_ac0_0_4\
        );

    \I__3262\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25072\
        );

    \I__3261\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25069\
        );

    \I__3260\ : InMux
    port map (
            O => \N__25075\,
            I => \N__25066\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__25072\,
            I => \N__25061\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__25069\,
            I => \N__25061\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__25066\,
            I => \sTrigCounterZ0Z_6\
        );

    \I__3256\ : Odrv12
    port map (
            O => \N__25061\,
            I => \sTrigCounterZ0Z_6\
        );

    \I__3255\ : InMux
    port map (
            O => \N__25056\,
            I => \N__25053\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__25053\,
            I => \N__25050\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__25050\,
            I => \un1_sTrigCounter_axbxc7_m7_0_a2_2\
        );

    \I__3252\ : InMux
    port map (
            O => \N__25047\,
            I => \N__25044\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__25044\,
            I => un1_reset_rpi_inv_2_i_1
        );

    \I__3250\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25038\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__25038\,
            I => \N__25035\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__25035\,
            I => \N_123\
        );

    \I__3247\ : InMux
    port map (
            O => \N__25032\,
            I => \N__25028\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__25031\,
            I => \N__25025\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__25028\,
            I => \N__25022\
        );

    \I__3244\ : InMux
    port map (
            O => \N__25025\,
            I => \N__25019\
        );

    \I__3243\ : Span4Mux_v
    port map (
            O => \N__25022\,
            I => \N__25016\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__25019\,
            I => \sTrigCounterZ0Z_7\
        );

    \I__3241\ : Odrv4
    port map (
            O => \N__25016\,
            I => \sTrigCounterZ0Z_7\
        );

    \I__3240\ : InMux
    port map (
            O => \N__25011\,
            I => \N__25008\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__25008\,
            I => \sEEPeriodZ0Z_14\
        );

    \I__3238\ : InMux
    port map (
            O => \N__25005\,
            I => \N__25002\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__25002\,
            I => \sEEPeriodZ0Z_15\
        );

    \I__3236\ : InMux
    port map (
            O => \N__24999\,
            I => \N__24996\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__24996\,
            I => \sEEPeriodZ0Z_8\
        );

    \I__3234\ : InMux
    port map (
            O => \N__24993\,
            I => \N__24990\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__24990\,
            I => \sEEPeriodZ0Z_9\
        );

    \I__3232\ : InMux
    port map (
            O => \N__24987\,
            I => \N__24984\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__24984\,
            I => \N__24981\
        );

    \I__3230\ : Span4Mux_v
    port map (
            O => \N__24981\,
            I => \N__24978\
        );

    \I__3229\ : Span4Mux_h
    port map (
            O => \N__24978\,
            I => \N__24975\
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__24975\,
            I => op_gt_op_gt_un13_striginternallto23_12
        );

    \I__3227\ : InMux
    port map (
            O => \N__24972\,
            I => \N__24969\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__24969\,
            I => \N__24966\
        );

    \I__3225\ : Span4Mux_h
    port map (
            O => \N__24966\,
            I => \N__24963\
        );

    \I__3224\ : Odrv4
    port map (
            O => \N__24963\,
            I => un1_reset_rpi_inv_2_i_o3_12
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__24960\,
            I => \N__24957\
        );

    \I__3222\ : InMux
    port map (
            O => \N__24957\,
            I => \N__24954\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__24954\,
            I => \N__24951\
        );

    \I__3220\ : Span4Mux_h
    port map (
            O => \N__24951\,
            I => \N__24948\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__24948\,
            I => op_gt_op_gt_un13_striginternallto23_15
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__24945\,
            I => \N__24935\
        );

    \I__3217\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24931\
        );

    \I__3216\ : InMux
    port map (
            O => \N__24943\,
            I => \N__24928\
        );

    \I__3215\ : InMux
    port map (
            O => \N__24942\,
            I => \N__24924\
        );

    \I__3214\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24921\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__24940\,
            I => \N__24918\
        );

    \I__3212\ : CascadeMux
    port map (
            O => \N__24939\,
            I => \N__24915\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__24938\,
            I => \N__24912\
        );

    \I__3210\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24904\
        );

    \I__3209\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24904\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__24931\,
            I => \N__24901\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__24928\,
            I => \N__24898\
        );

    \I__3206\ : InMux
    port map (
            O => \N__24927\,
            I => \N__24895\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__24924\,
            I => \N__24890\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__24921\,
            I => \N__24890\
        );

    \I__3203\ : InMux
    port map (
            O => \N__24918\,
            I => \N__24879\
        );

    \I__3202\ : InMux
    port map (
            O => \N__24915\,
            I => \N__24879\
        );

    \I__3201\ : InMux
    port map (
            O => \N__24912\,
            I => \N__24879\
        );

    \I__3200\ : InMux
    port map (
            O => \N__24911\,
            I => \N__24879\
        );

    \I__3199\ : InMux
    port map (
            O => \N__24910\,
            I => \N__24879\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__24909\,
            I => \N__24875\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__24904\,
            I => \N__24871\
        );

    \I__3196\ : Span4Mux_v
    port map (
            O => \N__24901\,
            I => \N__24866\
        );

    \I__3195\ : Span4Mux_v
    port map (
            O => \N__24898\,
            I => \N__24866\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__24895\,
            I => \N__24859\
        );

    \I__3193\ : Span4Mux_h
    port map (
            O => \N__24890\,
            I => \N__24859\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__24879\,
            I => \N__24859\
        );

    \I__3191\ : InMux
    port map (
            O => \N__24878\,
            I => \N__24852\
        );

    \I__3190\ : InMux
    port map (
            O => \N__24875\,
            I => \N__24852\
        );

    \I__3189\ : InMux
    port map (
            O => \N__24874\,
            I => \N__24852\
        );

    \I__3188\ : Odrv4
    port map (
            O => \N__24871\,
            I => \sEETrigInternal_prevZ0\
        );

    \I__3187\ : Odrv4
    port map (
            O => \N__24866\,
            I => \sEETrigInternal_prevZ0\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__24859\,
            I => \sEETrigInternal_prevZ0\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__24852\,
            I => \sEETrigInternal_prevZ0\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__24843\,
            I => \N__24840\
        );

    \I__3183\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24837\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__24837\,
            I => \N__24834\
        );

    \I__3181\ : Span4Mux_h
    port map (
            O => \N__24834\,
            I => \N__24831\
        );

    \I__3180\ : Span4Mux_v
    port map (
            O => \N__24831\,
            I => \N__24828\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__24828\,
            I => \N_5_0\
        );

    \I__3178\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24819\
        );

    \I__3177\ : InMux
    port map (
            O => \N__24824\,
            I => \N__24811\
        );

    \I__3176\ : InMux
    port map (
            O => \N__24823\,
            I => \N__24811\
        );

    \I__3175\ : InMux
    port map (
            O => \N__24822\,
            I => \N__24808\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__24819\,
            I => \N__24805\
        );

    \I__3173\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24800\
        );

    \I__3172\ : InMux
    port map (
            O => \N__24817\,
            I => \N__24800\
        );

    \I__3171\ : InMux
    port map (
            O => \N__24816\,
            I => \N__24794\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__24811\,
            I => \N__24791\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__24808\,
            I => \N__24787\
        );

    \I__3168\ : Span4Mux_v
    port map (
            O => \N__24805\,
            I => \N__24782\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__24800\,
            I => \N__24782\
        );

    \I__3166\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24779\
        );

    \I__3165\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24776\
        );

    \I__3164\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24773\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__24794\,
            I => \N__24768\
        );

    \I__3162\ : Span4Mux_v
    port map (
            O => \N__24791\,
            I => \N__24768\
        );

    \I__3161\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24765\
        );

    \I__3160\ : Span4Mux_h
    port map (
            O => \N__24787\,
            I => \N__24758\
        );

    \I__3159\ : Span4Mux_v
    port map (
            O => \N__24782\,
            I => \N__24758\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__24779\,
            I => \N__24758\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__24776\,
            I => \un4_speriod_cry_23_THRU_CO\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__24773\,
            I => \un4_speriod_cry_23_THRU_CO\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__24768\,
            I => \un4_speriod_cry_23_THRU_CO\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__24765\,
            I => \un4_speriod_cry_23_THRU_CO\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__24758\,
            I => \un4_speriod_cry_23_THRU_CO\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__24747\,
            I => \un1_reset_rpi_inv_2_i_1_1_0_cascade_\
        );

    \I__3151\ : CascadeMux
    port map (
            O => \N__24744\,
            I => \un1_sTrigCounter_ac0_0_0_cascade_\
        );

    \I__3150\ : InMux
    port map (
            O => \N__24741\,
            I => \N__24737\
        );

    \I__3149\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24734\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__24737\,
            I => \N__24731\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__24734\,
            I => \N__24726\
        );

    \I__3146\ : Span4Mux_h
    port map (
            O => \N__24731\,
            I => \N__24726\
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__24726\,
            I => un1_reset_rpi_inv_2_i_o3_0_0
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__24723\,
            I => \un1_sTrigCounter_ac0_0_2_0_cascade_\
        );

    \I__3143\ : InMux
    port map (
            O => \N__24720\,
            I => \N__24715\
        );

    \I__3142\ : InMux
    port map (
            O => \N__24719\,
            I => \N__24710\
        );

    \I__3141\ : InMux
    port map (
            O => \N__24718\,
            I => \N__24707\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__24715\,
            I => \N__24704\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__24714\,
            I => \N__24700\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__24713\,
            I => \N__24695\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__24710\,
            I => \N__24691\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__24707\,
            I => \N__24686\
        );

    \I__3135\ : Span4Mux_v
    port map (
            O => \N__24704\,
            I => \N__24686\
        );

    \I__3134\ : InMux
    port map (
            O => \N__24703\,
            I => \N__24683\
        );

    \I__3133\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24680\
        );

    \I__3132\ : InMux
    port map (
            O => \N__24699\,
            I => \N__24677\
        );

    \I__3131\ : InMux
    port map (
            O => \N__24698\,
            I => \N__24674\
        );

    \I__3130\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24669\
        );

    \I__3129\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24669\
        );

    \I__3128\ : Span4Mux_v
    port map (
            O => \N__24691\,
            I => \N__24664\
        );

    \I__3127\ : Span4Mux_v
    port map (
            O => \N__24686\,
            I => \N__24664\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__24683\,
            I => \un10_trig_prev_cry_7_THRU_CO\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__24680\,
            I => \un10_trig_prev_cry_7_THRU_CO\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__24677\,
            I => \un10_trig_prev_cry_7_THRU_CO\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__24674\,
            I => \un10_trig_prev_cry_7_THRU_CO\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__24669\,
            I => \un10_trig_prev_cry_7_THRU_CO\
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__24664\,
            I => \un10_trig_prev_cry_7_THRU_CO\
        );

    \I__3120\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24648\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__24648\,
            I => \N__24642\
        );

    \I__3118\ : InMux
    port map (
            O => \N__24647\,
            I => \N__24637\
        );

    \I__3117\ : InMux
    port map (
            O => \N__24646\,
            I => \N__24637\
        );

    \I__3116\ : InMux
    port map (
            O => \N__24645\,
            I => \N__24634\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__24642\,
            I => \sTrigCounterZ0Z_5\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__24637\,
            I => \sTrigCounterZ0Z_5\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__24634\,
            I => \sTrigCounterZ0Z_5\
        );

    \I__3112\ : InMux
    port map (
            O => \N__24627\,
            I => \N__24621\
        );

    \I__3111\ : InMux
    port map (
            O => \N__24626\,
            I => \N__24621\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__24621\,
            I => \un1_sTrigCounter_ac0_0_2\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__24618\,
            I => \un1_sTrigCounter_ac0_3_out_cascade_\
        );

    \I__3108\ : InMux
    port map (
            O => \N__24615\,
            I => \N__24603\
        );

    \I__3107\ : InMux
    port map (
            O => \N__24614\,
            I => \N__24603\
        );

    \I__3106\ : InMux
    port map (
            O => \N__24613\,
            I => \N__24603\
        );

    \I__3105\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24599\
        );

    \I__3104\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24594\
        );

    \I__3103\ : InMux
    port map (
            O => \N__24610\,
            I => \N__24594\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__24603\,
            I => \N__24591\
        );

    \I__3101\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24588\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__24599\,
            I => \N__24585\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__24594\,
            I => \sTrigCounterZ0Z_2\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__24591\,
            I => \sTrigCounterZ0Z_2\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__24588\,
            I => \sTrigCounterZ0Z_2\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__24585\,
            I => \sTrigCounterZ0Z_2\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__24576\,
            I => \N__24573\
        );

    \I__3094\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24570\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__24570\,
            I => g1_0_1_0
        );

    \I__3092\ : InMux
    port map (
            O => \N__24567\,
            I => \N__24564\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__24564\,
            I => g1_3_0
        );

    \I__3090\ : InMux
    port map (
            O => \N__24561\,
            I => \N__24558\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__24558\,
            I => \sEEPeriodZ0Z_10\
        );

    \I__3088\ : InMux
    port map (
            O => \N__24555\,
            I => \N__24552\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__24552\,
            I => \sEEPeriodZ0Z_11\
        );

    \I__3086\ : InMux
    port map (
            O => \N__24549\,
            I => \N__24546\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__24546\,
            I => \sEEPeriodZ0Z_12\
        );

    \I__3084\ : InMux
    port map (
            O => \N__24543\,
            I => \N__24540\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__24540\,
            I => \sEEPeriodZ0Z_13\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__24537\,
            I => \N__24534\
        );

    \I__3081\ : InMux
    port map (
            O => \N__24534\,
            I => \N__24531\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__24531\,
            I => un10_trig_prev_7
        );

    \I__3079\ : InMux
    port map (
            O => \N__24528\,
            I => \N__24525\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__24525\,
            I => \sTrigCounter_i_7\
        );

    \I__3077\ : InMux
    port map (
            O => \N__24522\,
            I => \bfn_9_9_0_\
        );

    \I__3076\ : CEMux
    port map (
            O => \N__24519\,
            I => \N__24516\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__24516\,
            I => \N__24513\
        );

    \I__3074\ : Odrv4
    port map (
            O => \N__24513\,
            I => \sAddress_RNI9IH12_1Z0Z_1\
        );

    \I__3073\ : InMux
    port map (
            O => \N__24510\,
            I => \N__24503\
        );

    \I__3072\ : InMux
    port map (
            O => \N__24509\,
            I => \N__24498\
        );

    \I__3071\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24498\
        );

    \I__3070\ : InMux
    port map (
            O => \N__24507\,
            I => \N__24495\
        );

    \I__3069\ : InMux
    port map (
            O => \N__24506\,
            I => \N__24492\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__24503\,
            I => \N__24485\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__24498\,
            I => \N__24482\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__24495\,
            I => \N__24477\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__24492\,
            I => \N__24477\
        );

    \I__3064\ : InMux
    port map (
            O => \N__24491\,
            I => \N__24470\
        );

    \I__3063\ : InMux
    port map (
            O => \N__24490\,
            I => \N__24470\
        );

    \I__3062\ : InMux
    port map (
            O => \N__24489\,
            I => \N__24470\
        );

    \I__3061\ : InMux
    port map (
            O => \N__24488\,
            I => \N__24461\
        );

    \I__3060\ : Span4Mux_v
    port map (
            O => \N__24485\,
            I => \N__24458\
        );

    \I__3059\ : Span4Mux_v
    port map (
            O => \N__24482\,
            I => \N__24451\
        );

    \I__3058\ : Span4Mux_h
    port map (
            O => \N__24477\,
            I => \N__24451\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__24470\,
            I => \N__24451\
        );

    \I__3056\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24438\
        );

    \I__3055\ : InMux
    port map (
            O => \N__24468\,
            I => \N__24438\
        );

    \I__3054\ : InMux
    port map (
            O => \N__24467\,
            I => \N__24438\
        );

    \I__3053\ : InMux
    port map (
            O => \N__24466\,
            I => \N__24438\
        );

    \I__3052\ : InMux
    port map (
            O => \N__24465\,
            I => \N__24438\
        );

    \I__3051\ : InMux
    port map (
            O => \N__24464\,
            I => \N__24438\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__24461\,
            I => \trig_prevZ0\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__24458\,
            I => \trig_prevZ0\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__24451\,
            I => \trig_prevZ0\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__24438\,
            I => \trig_prevZ0\
        );

    \I__3046\ : InMux
    port map (
            O => \N__24429\,
            I => \N__24425\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__24428\,
            I => \N__24422\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__24425\,
            I => \N__24419\
        );

    \I__3043\ : InMux
    port map (
            O => \N__24422\,
            I => \N__24416\
        );

    \I__3042\ : Span4Mux_v
    port map (
            O => \N__24419\,
            I => \N__24413\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__24416\,
            I => \N__24410\
        );

    \I__3040\ : Odrv4
    port map (
            O => \N__24413\,
            I => un3_trig_0_3
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__24410\,
            I => un3_trig_0_3
        );

    \I__3038\ : InMux
    port map (
            O => \N__24405\,
            I => \N__24402\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__24402\,
            I => g1_0_0_2
        );

    \I__3036\ : InMux
    port map (
            O => \N__24399\,
            I => \N__24396\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__24396\,
            I => \N__24393\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__24393\,
            I => g1_0_0
        );

    \I__3033\ : InMux
    port map (
            O => \N__24390\,
            I => \N__24387\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__24387\,
            I => g1_0
        );

    \I__3031\ : InMux
    port map (
            O => \N__24384\,
            I => \N__24381\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__24381\,
            I => \N__24373\
        );

    \I__3029\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24370\
        );

    \I__3028\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24365\
        );

    \I__3027\ : InMux
    port map (
            O => \N__24378\,
            I => \N__24365\
        );

    \I__3026\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24362\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__24376\,
            I => \N__24358\
        );

    \I__3024\ : Span4Mux_v
    port map (
            O => \N__24373\,
            I => \N__24352\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__24370\,
            I => \N__24352\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__24365\,
            I => \N__24347\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__24362\,
            I => \N__24347\
        );

    \I__3020\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24344\
        );

    \I__3019\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24339\
        );

    \I__3018\ : InMux
    port map (
            O => \N__24357\,
            I => \N__24339\
        );

    \I__3017\ : Span4Mux_v
    port map (
            O => \N__24352\,
            I => \N__24332\
        );

    \I__3016\ : Span4Mux_h
    port map (
            O => \N__24347\,
            I => \N__24332\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__24344\,
            I => \N__24332\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__24339\,
            I => \N__24329\
        );

    \I__3013\ : Span4Mux_v
    port map (
            O => \N__24332\,
            I => \N__24326\
        );

    \I__3012\ : Odrv12
    port map (
            O => \N__24329\,
            I => \sPeriod_prevZ0\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__24326\,
            I => \sPeriod_prevZ0\
        );

    \I__3010\ : IoInMux
    port map (
            O => \N__24321\,
            I => \N__24318\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__24318\,
            I => \N__24315\
        );

    \I__3008\ : Span4Mux_s1_h
    port map (
            O => \N__24315\,
            I => \N__24311\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__24314\,
            I => \N__24306\
        );

    \I__3006\ : Span4Mux_h
    port map (
            O => \N__24311\,
            I => \N__24303\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__24310\,
            I => \N__24300\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__24309\,
            I => \N__24297\
        );

    \I__3003\ : InMux
    port map (
            O => \N__24306\,
            I => \N__24294\
        );

    \I__3002\ : Span4Mux_h
    port map (
            O => \N__24303\,
            I => \N__24291\
        );

    \I__3001\ : InMux
    port map (
            O => \N__24300\,
            I => \N__24288\
        );

    \I__3000\ : InMux
    port map (
            O => \N__24297\,
            I => \N__24285\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__24294\,
            I => \N__24282\
        );

    \I__2998\ : Span4Mux_v
    port map (
            O => \N__24291\,
            I => \N__24277\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__24288\,
            I => \N__24277\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__24285\,
            I => \N__24274\
        );

    \I__2995\ : Span4Mux_h
    port map (
            O => \N__24282\,
            I => \N__24265\
        );

    \I__2994\ : Span4Mux_v
    port map (
            O => \N__24277\,
            I => \N__24265\
        );

    \I__2993\ : Span4Mux_h
    port map (
            O => \N__24274\,
            I => \N__24265\
        );

    \I__2992\ : InMux
    port map (
            O => \N__24273\,
            I => \N__24260\
        );

    \I__2991\ : InMux
    port map (
            O => \N__24272\,
            I => \N__24260\
        );

    \I__2990\ : Span4Mux_v
    port map (
            O => \N__24265\,
            I => \N__24252\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__24260\,
            I => \N__24252\
        );

    \I__2988\ : InMux
    port map (
            O => \N__24259\,
            I => \N__24247\
        );

    \I__2987\ : InMux
    port map (
            O => \N__24258\,
            I => \N__24247\
        );

    \I__2986\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24244\
        );

    \I__2985\ : Span4Mux_h
    port map (
            O => \N__24252\,
            I => \N__24241\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__24247\,
            I => \N__24236\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__24244\,
            I => \N__24236\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__24241\,
            I => \LED_MODE_c\
        );

    \I__2981\ : Odrv12
    port map (
            O => \N__24236\,
            I => \LED_MODE_c\
        );

    \I__2980\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24225\
        );

    \I__2979\ : InMux
    port map (
            O => \N__24230\,
            I => \N__24222\
        );

    \I__2978\ : InMux
    port map (
            O => \N__24229\,
            I => \N__24219\
        );

    \I__2977\ : InMux
    port map (
            O => \N__24228\,
            I => \N__24216\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__24225\,
            I => \N__24213\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__24222\,
            I => \sTrigCounterZ0Z_4\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__24219\,
            I => \sTrigCounterZ0Z_4\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__24216\,
            I => \sTrigCounterZ0Z_4\
        );

    \I__2972\ : Odrv4
    port map (
            O => \N__24213\,
            I => \sTrigCounterZ0Z_4\
        );

    \I__2971\ : InMux
    port map (
            O => \N__24204\,
            I => \N__24197\
        );

    \I__2970\ : InMux
    port map (
            O => \N__24203\,
            I => \N__24194\
        );

    \I__2969\ : InMux
    port map (
            O => \N__24202\,
            I => \N__24189\
        );

    \I__2968\ : InMux
    port map (
            O => \N__24201\,
            I => \N__24189\
        );

    \I__2967\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24186\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__24197\,
            I => \sTrigCounterZ0Z_3\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__24194\,
            I => \sTrigCounterZ0Z_3\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__24189\,
            I => \sTrigCounterZ0Z_3\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__24186\,
            I => \sTrigCounterZ0Z_3\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__24177\,
            I => \N__24173\
        );

    \I__2961\ : InMux
    port map (
            O => \N__24176\,
            I => \N__24168\
        );

    \I__2960\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24168\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__24168\,
            I => \sEETrigCounterZ0Z_4\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__24165\,
            I => \N__24160\
        );

    \I__2957\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24155\
        );

    \I__2956\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24155\
        );

    \I__2955\ : InMux
    port map (
            O => \N__24160\,
            I => \N__24152\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__24155\,
            I => un8_trig_prev_0_c5_a0_0
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__24152\,
            I => un8_trig_prev_0_c5_a0_0
        );

    \I__2952\ : InMux
    port map (
            O => \N__24147\,
            I => \N__24144\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__24144\,
            I => \sTrigCounter_i_0\
        );

    \I__2950\ : InMux
    port map (
            O => \N__24141\,
            I => \N__24138\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__24138\,
            I => \sTrigCounter_i_1\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__24135\,
            I => \N__24132\
        );

    \I__2947\ : InMux
    port map (
            O => \N__24132\,
            I => \N__24129\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__24129\,
            I => \sTrigCounter_i_2\
        );

    \I__2945\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24123\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__24123\,
            I => \sTrigCounter_i_3\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__24120\,
            I => \N__24117\
        );

    \I__2942\ : InMux
    port map (
            O => \N__24117\,
            I => \N__24114\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__24114\,
            I => un10_trig_prev_4
        );

    \I__2940\ : InMux
    port map (
            O => \N__24111\,
            I => \N__24108\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__24108\,
            I => \sTrigCounter_i_4\
        );

    \I__2938\ : CascadeMux
    port map (
            O => \N__24105\,
            I => \N__24102\
        );

    \I__2937\ : InMux
    port map (
            O => \N__24102\,
            I => \N__24099\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__24099\,
            I => un10_trig_prev_5
        );

    \I__2935\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24093\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__24093\,
            I => \sTrigCounter_i_5\
        );

    \I__2933\ : CascadeMux
    port map (
            O => \N__24090\,
            I => \N__24087\
        );

    \I__2932\ : InMux
    port map (
            O => \N__24087\,
            I => \N__24084\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__24084\,
            I => un10_trig_prev_6
        );

    \I__2930\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24078\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__24078\,
            I => \N__24075\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__24075\,
            I => \sTrigCounter_i_6\
        );

    \I__2927\ : InMux
    port map (
            O => \N__24072\,
            I => \N__24069\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__24069\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2\
        );

    \I__2925\ : InMux
    port map (
            O => \N__24066\,
            I => \N__24060\
        );

    \I__2924\ : InMux
    port map (
            O => \N__24065\,
            I => \N__24060\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__24060\,
            I => \N__24053\
        );

    \I__2922\ : InMux
    port map (
            O => \N__24059\,
            I => \N__24048\
        );

    \I__2921\ : InMux
    port map (
            O => \N__24058\,
            I => \N__24048\
        );

    \I__2920\ : InMux
    port map (
            O => \N__24057\,
            I => \N__24045\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__24056\,
            I => \N__24042\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__24053\,
            I => \N__24033\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__24048\,
            I => \N__24033\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__24045\,
            I => \N__24033\
        );

    \I__2915\ : InMux
    port map (
            O => \N__24042\,
            I => \N__24028\
        );

    \I__2914\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24028\
        );

    \I__2913\ : InMux
    port map (
            O => \N__24040\,
            I => \N__24025\
        );

    \I__2912\ : Span4Mux_v
    port map (
            O => \N__24033\,
            I => \N__24021\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__24028\,
            I => \N__24018\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__24025\,
            I => \N__24015\
        );

    \I__2909\ : InMux
    port map (
            O => \N__24024\,
            I => \N__24012\
        );

    \I__2908\ : Span4Mux_v
    port map (
            O => \N__24021\,
            I => \N__24009\
        );

    \I__2907\ : Span4Mux_v
    port map (
            O => \N__24018\,
            I => \N__24006\
        );

    \I__2906\ : Span4Mux_v
    port map (
            O => \N__24015\,
            I => \N__24001\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__24012\,
            I => \N__24001\
        );

    \I__2904\ : Span4Mux_h
    port map (
            O => \N__24009\,
            I => \N__23998\
        );

    \I__2903\ : Span4Mux_v
    port map (
            O => \N__24006\,
            I => \N__23995\
        );

    \I__2902\ : Span4Mux_h
    port map (
            O => \N__24001\,
            I => \N__23992\
        );

    \I__2901\ : Sp12to4
    port map (
            O => \N__23998\,
            I => \N__23987\
        );

    \I__2900\ : Sp12to4
    port map (
            O => \N__23995\,
            I => \N__23987\
        );

    \I__2899\ : Span4Mux_v
    port map (
            O => \N__23992\,
            I => \N__23984\
        );

    \I__2898\ : Odrv12
    port map (
            O => \N__23987\,
            I => trig_ext_c
        );

    \I__2897\ : Odrv4
    port map (
            O => \N__23984\,
            I => trig_ext_c
        );

    \I__2896\ : InMux
    port map (
            O => \N__23979\,
            I => \N__23973\
        );

    \I__2895\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23973\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__23973\,
            I => \N__23967\
        );

    \I__2893\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23959\
        );

    \I__2892\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23959\
        );

    \I__2891\ : InMux
    port map (
            O => \N__23970\,
            I => \N__23956\
        );

    \I__2890\ : Span4Mux_h
    port map (
            O => \N__23967\,
            I => \N__23953\
        );

    \I__2889\ : InMux
    port map (
            O => \N__23966\,
            I => \N__23948\
        );

    \I__2888\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23948\
        );

    \I__2887\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23945\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__23959\,
            I => \N__23940\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__23956\,
            I => \N__23940\
        );

    \I__2884\ : Span4Mux_h
    port map (
            O => \N__23953\,
            I => \N__23935\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__23948\,
            I => \N__23935\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__23945\,
            I => \N__23932\
        );

    \I__2881\ : Span4Mux_v
    port map (
            O => \N__23940\,
            I => \N__23928\
        );

    \I__2880\ : Span4Mux_v
    port map (
            O => \N__23935\,
            I => \N__23925\
        );

    \I__2879\ : Span4Mux_v
    port map (
            O => \N__23932\,
            I => \N__23922\
        );

    \I__2878\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23919\
        );

    \I__2877\ : Sp12to4
    port map (
            O => \N__23928\,
            I => \N__23910\
        );

    \I__2876\ : Sp12to4
    port map (
            O => \N__23925\,
            I => \N__23910\
        );

    \I__2875\ : Sp12to4
    port map (
            O => \N__23922\,
            I => \N__23910\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__23919\,
            I => \N__23910\
        );

    \I__2873\ : Odrv12
    port map (
            O => \N__23910\,
            I => trig_rpi_c
        );

    \I__2872\ : InMux
    port map (
            O => \N__23907\,
            I => \N__23903\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__23906\,
            I => \N__23896\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__23903\,
            I => \N__23893\
        );

    \I__2869\ : InMux
    port map (
            O => \N__23902\,
            I => \N__23887\
        );

    \I__2868\ : InMux
    port map (
            O => \N__23901\,
            I => \N__23887\
        );

    \I__2867\ : InMux
    port map (
            O => \N__23900\,
            I => \N__23884\
        );

    \I__2866\ : InMux
    port map (
            O => \N__23899\,
            I => \N__23879\
        );

    \I__2865\ : InMux
    port map (
            O => \N__23896\,
            I => \N__23879\
        );

    \I__2864\ : Span4Mux_v
    port map (
            O => \N__23893\,
            I => \N__23874\
        );

    \I__2863\ : InMux
    port map (
            O => \N__23892\,
            I => \N__23871\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__23887\,
            I => \N__23864\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__23884\,
            I => \N__23864\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__23879\,
            I => \N__23864\
        );

    \I__2859\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23859\
        );

    \I__2858\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23859\
        );

    \I__2857\ : Span4Mux_h
    port map (
            O => \N__23874\,
            I => \N__23856\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__23871\,
            I => \N__23853\
        );

    \I__2855\ : Span4Mux_h
    port map (
            O => \N__23864\,
            I => \N__23848\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__23859\,
            I => \N__23848\
        );

    \I__2853\ : Sp12to4
    port map (
            O => \N__23856\,
            I => \N__23845\
        );

    \I__2852\ : Span12Mux_h
    port map (
            O => \N__23853\,
            I => \N__23840\
        );

    \I__2851\ : Sp12to4
    port map (
            O => \N__23848\,
            I => \N__23840\
        );

    \I__2850\ : Span12Mux_h
    port map (
            O => \N__23845\,
            I => \N__23837\
        );

    \I__2849\ : Span12Mux_v
    port map (
            O => \N__23840\,
            I => \N__23834\
        );

    \I__2848\ : Span12Mux_v
    port map (
            O => \N__23837\,
            I => \N__23829\
        );

    \I__2847\ : Span12Mux_h
    port map (
            O => \N__23834\,
            I => \N__23829\
        );

    \I__2846\ : Odrv12
    port map (
            O => \N__23829\,
            I => trig_ft_c
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__23826\,
            I => \un8_trig_prev_0_c5_a0_0_0_cascade_\
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__23823\,
            I => \un8_trig_prev_0_c4_a0_1_cascade_\
        );

    \I__2843\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23811\
        );

    \I__2842\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23811\
        );

    \I__2841\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23811\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__23811\,
            I => \sEETrigCounterZ0Z_5\
        );

    \I__2839\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23802\
        );

    \I__2838\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23802\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__23802\,
            I => \sEETrigCounterZ0Z_6\
        );

    \I__2836\ : InMux
    port map (
            O => \N__23799\,
            I => \N__23796\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__23796\,
            I => \sEETrigCounterZ0Z_7\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__23793\,
            I => \un8_trig_prev_0_c7_a0_1_cascade_\
        );

    \I__2833\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23784\
        );

    \I__2832\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23784\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__23784\,
            I => un8_trig_prev_0_c4_a0_1
        );

    \I__2830\ : InMux
    port map (
            O => \N__23781\,
            I => \N__23778\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__23778\,
            I => \N__23775\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__23775\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15\
        );

    \I__2827\ : InMux
    port map (
            O => \N__23772\,
            I => \N__23769\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__23769\,
            I => \N__23766\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__23766\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11\
        );

    \I__2824\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23760\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__23760\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10\
        );

    \I__2822\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23751\
        );

    \I__2821\ : InMux
    port map (
            O => \N__23756\,
            I => \N__23751\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__23751\,
            I => \N__23747\
        );

    \I__2819\ : InMux
    port map (
            O => \N__23750\,
            I => \N__23744\
        );

    \I__2818\ : Odrv12
    port map (
            O => \N__23747\,
            I => \spi_master_inst.sclk_gen_u0.N_158_7\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__23744\,
            I => \spi_master_inst.sclk_gen_u0.N_158_7\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__23739\,
            I => \N__23736\
        );

    \I__2815\ : InMux
    port map (
            O => \N__23736\,
            I => \N__23732\
        );

    \I__2814\ : InMux
    port map (
            O => \N__23735\,
            I => \N__23729\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__23732\,
            I => \N__23721\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__23729\,
            I => \N__23721\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__23728\,
            I => \N__23718\
        );

    \I__2810\ : InMux
    port map (
            O => \N__23727\,
            I => \N__23712\
        );

    \I__2809\ : InMux
    port map (
            O => \N__23726\,
            I => \N__23712\
        );

    \I__2808\ : Span4Mux_h
    port map (
            O => \N__23721\,
            I => \N__23709\
        );

    \I__2807\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23704\
        );

    \I__2806\ : InMux
    port map (
            O => \N__23717\,
            I => \N__23704\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__23712\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__23709\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__23704\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__23697\,
            I => \spi_master_inst.sclk_gen_u0.N_158_7_cascade_\
        );

    \I__2801\ : InMux
    port map (
            O => \N__23694\,
            I => \N__23689\
        );

    \I__2800\ : InMux
    port map (
            O => \N__23693\,
            I => \N__23683\
        );

    \I__2799\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23683\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__23689\,
            I => \N__23679\
        );

    \I__2797\ : InMux
    port map (
            O => \N__23688\,
            I => \N__23675\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__23683\,
            I => \N__23672\
        );

    \I__2795\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23669\
        );

    \I__2794\ : Span12Mux_s11_h
    port map (
            O => \N__23679\,
            I => \N__23666\
        );

    \I__2793\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23663\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__23675\,
            I => \N__23660\
        );

    \I__2791\ : Odrv4
    port map (
            O => \N__23672\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__23669\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\
        );

    \I__2789\ : Odrv12
    port map (
            O => \N__23666\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__23663\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\
        );

    \I__2787\ : Odrv12
    port map (
            O => \N__23660\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\
        );

    \I__2786\ : InMux
    port map (
            O => \N__23649\,
            I => \N__23646\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__23646\,
            I => \spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0\
        );

    \I__2784\ : InMux
    port map (
            O => \N__23643\,
            I => \N__23636\
        );

    \I__2783\ : InMux
    port map (
            O => \N__23642\,
            I => \N__23636\
        );

    \I__2782\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23633\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__23636\,
            I => \spi_master_inst.sclk_gen_u0.falling_count_start_iZ0\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__23633\,
            I => \spi_master_inst.sclk_gen_u0.falling_count_start_iZ0\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__23628\,
            I => \N__23625\
        );

    \I__2778\ : InMux
    port map (
            O => \N__23625\,
            I => \N__23622\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__23622\,
            I => \N__23619\
        );

    \I__2776\ : Odrv4
    port map (
            O => \N__23619\,
            I => un3_trig_0_0
        );

    \I__2775\ : CascadeMux
    port map (
            O => \N__23616\,
            I => \un3_trig_0_0_cascade_\
        );

    \I__2774\ : InMux
    port map (
            O => \N__23613\,
            I => \N__23610\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__23610\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2\
        );

    \I__2772\ : InMux
    port map (
            O => \N__23607\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4\
        );

    \I__2771\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23601\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__23601\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO\
        );

    \I__2769\ : InMux
    port map (
            O => \N__23598\,
            I => \N__23595\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__23595\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO\
        );

    \I__2767\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23589\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__23589\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12\
        );

    \I__2765\ : InMux
    port map (
            O => \N__23586\,
            I => \N__23583\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__23583\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2\
        );

    \I__2763\ : InMux
    port map (
            O => \N__23580\,
            I => \N__23577\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__23577\,
            I => \N__23574\
        );

    \I__2761\ : Odrv12
    port map (
            O => \N__23574\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3\
        );

    \I__2760\ : InMux
    port map (
            O => \N__23571\,
            I => \N__23568\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__23568\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4\
        );

    \I__2758\ : InMux
    port map (
            O => \N__23565\,
            I => \N__23562\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__23562\,
            I => \N__23559\
        );

    \I__2756\ : Span4Mux_h
    port map (
            O => \N__23559\,
            I => \N__23556\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__23556\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5\
        );

    \I__2754\ : InMux
    port map (
            O => \N__23553\,
            I => un1_button_debounce_counter_cry_21
        );

    \I__2753\ : InMux
    port map (
            O => \N__23550\,
            I => \bfn_8_20_0_\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__23547\,
            I => \N__23544\
        );

    \I__2751\ : InMux
    port map (
            O => \N__23544\,
            I => \N__23540\
        );

    \I__2750\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23537\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__23540\,
            I => \N__23534\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__23537\,
            I => \button_debounce_counterZ0Z_23\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__23534\,
            I => \button_debounce_counterZ0Z_23\
        );

    \I__2746\ : InMux
    port map (
            O => \N__23529\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0\
        );

    \I__2745\ : InMux
    port map (
            O => \N__23526\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1\
        );

    \I__2744\ : InMux
    port map (
            O => \N__23523\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2\
        );

    \I__2743\ : InMux
    port map (
            O => \N__23520\,
            I => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__23517\,
            I => \N__23513\
        );

    \I__2741\ : InMux
    port map (
            O => \N__23516\,
            I => \N__23510\
        );

    \I__2740\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23507\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__23510\,
            I => \button_debounce_counterZ0Z_13\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__23507\,
            I => \button_debounce_counterZ0Z_13\
        );

    \I__2737\ : InMux
    port map (
            O => \N__23502\,
            I => un1_button_debounce_counter_cry_12
        );

    \I__2736\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23495\
        );

    \I__2735\ : InMux
    port map (
            O => \N__23498\,
            I => \N__23492\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__23495\,
            I => \button_debounce_counterZ0Z_14\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__23492\,
            I => \button_debounce_counterZ0Z_14\
        );

    \I__2732\ : InMux
    port map (
            O => \N__23487\,
            I => un1_button_debounce_counter_cry_13
        );

    \I__2731\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23480\
        );

    \I__2730\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23477\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__23480\,
            I => \button_debounce_counterZ0Z_15\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__23477\,
            I => \button_debounce_counterZ0Z_15\
        );

    \I__2727\ : InMux
    port map (
            O => \N__23472\,
            I => un1_button_debounce_counter_cry_14
        );

    \I__2726\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23465\
        );

    \I__2725\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23462\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__23465\,
            I => \button_debounce_counterZ0Z_16\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__23462\,
            I => \button_debounce_counterZ0Z_16\
        );

    \I__2722\ : InMux
    port map (
            O => \N__23457\,
            I => un1_button_debounce_counter_cry_15
        );

    \I__2721\ : InMux
    port map (
            O => \N__23454\,
            I => \N__23451\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__23451\,
            I => \N__23447\
        );

    \I__2719\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23444\
        );

    \I__2718\ : Odrv12
    port map (
            O => \N__23447\,
            I => \button_debounce_counterZ0Z_17\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__23444\,
            I => \button_debounce_counterZ0Z_17\
        );

    \I__2716\ : InMux
    port map (
            O => \N__23439\,
            I => \bfn_8_19_0_\
        );

    \I__2715\ : InMux
    port map (
            O => \N__23436\,
            I => \N__23433\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__23433\,
            I => \N__23430\
        );

    \I__2713\ : Span4Mux_v
    port map (
            O => \N__23430\,
            I => \N__23426\
        );

    \I__2712\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23423\
        );

    \I__2711\ : Odrv4
    port map (
            O => \N__23426\,
            I => \button_debounce_counterZ0Z_18\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__23423\,
            I => \button_debounce_counterZ0Z_18\
        );

    \I__2709\ : InMux
    port map (
            O => \N__23418\,
            I => un1_button_debounce_counter_cry_17
        );

    \I__2708\ : InMux
    port map (
            O => \N__23415\,
            I => \N__23412\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__23412\,
            I => \N__23408\
        );

    \I__2706\ : InMux
    port map (
            O => \N__23411\,
            I => \N__23405\
        );

    \I__2705\ : Odrv12
    port map (
            O => \N__23408\,
            I => \button_debounce_counterZ0Z_19\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__23405\,
            I => \button_debounce_counterZ0Z_19\
        );

    \I__2703\ : InMux
    port map (
            O => \N__23400\,
            I => un1_button_debounce_counter_cry_18
        );

    \I__2702\ : CascadeMux
    port map (
            O => \N__23397\,
            I => \N__23394\
        );

    \I__2701\ : InMux
    port map (
            O => \N__23394\,
            I => \N__23391\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__23391\,
            I => \N__23388\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__23388\,
            I => \N__23384\
        );

    \I__2698\ : InMux
    port map (
            O => \N__23387\,
            I => \N__23381\
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__23384\,
            I => \button_debounce_counterZ0Z_20\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__23381\,
            I => \button_debounce_counterZ0Z_20\
        );

    \I__2695\ : InMux
    port map (
            O => \N__23376\,
            I => un1_button_debounce_counter_cry_19
        );

    \I__2694\ : InMux
    port map (
            O => \N__23373\,
            I => un1_button_debounce_counter_cry_20
        );

    \I__2693\ : InMux
    port map (
            O => \N__23370\,
            I => un1_button_debounce_counter_cry_4
        );

    \I__2692\ : InMux
    port map (
            O => \N__23367\,
            I => \N__23363\
        );

    \I__2691\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23360\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__23363\,
            I => \button_debounce_counterZ0Z_6\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__23360\,
            I => \button_debounce_counterZ0Z_6\
        );

    \I__2688\ : InMux
    port map (
            O => \N__23355\,
            I => un1_button_debounce_counter_cry_5
        );

    \I__2687\ : InMux
    port map (
            O => \N__23352\,
            I => \N__23348\
        );

    \I__2686\ : InMux
    port map (
            O => \N__23351\,
            I => \N__23345\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__23348\,
            I => \button_debounce_counterZ0Z_7\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__23345\,
            I => \button_debounce_counterZ0Z_7\
        );

    \I__2683\ : InMux
    port map (
            O => \N__23340\,
            I => un1_button_debounce_counter_cry_6
        );

    \I__2682\ : InMux
    port map (
            O => \N__23337\,
            I => \N__23333\
        );

    \I__2681\ : InMux
    port map (
            O => \N__23336\,
            I => \N__23330\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__23333\,
            I => \button_debounce_counterZ0Z_8\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__23330\,
            I => \button_debounce_counterZ0Z_8\
        );

    \I__2678\ : InMux
    port map (
            O => \N__23325\,
            I => un1_button_debounce_counter_cry_7
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__23322\,
            I => \N__23318\
        );

    \I__2676\ : InMux
    port map (
            O => \N__23321\,
            I => \N__23315\
        );

    \I__2675\ : InMux
    port map (
            O => \N__23318\,
            I => \N__23312\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__23315\,
            I => \button_debounce_counterZ0Z_9\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__23312\,
            I => \button_debounce_counterZ0Z_9\
        );

    \I__2672\ : InMux
    port map (
            O => \N__23307\,
            I => \bfn_8_18_0_\
        );

    \I__2671\ : InMux
    port map (
            O => \N__23304\,
            I => \N__23300\
        );

    \I__2670\ : InMux
    port map (
            O => \N__23303\,
            I => \N__23297\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__23300\,
            I => \button_debounce_counterZ0Z_10\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__23297\,
            I => \button_debounce_counterZ0Z_10\
        );

    \I__2667\ : InMux
    port map (
            O => \N__23292\,
            I => un1_button_debounce_counter_cry_9
        );

    \I__2666\ : InMux
    port map (
            O => \N__23289\,
            I => \N__23285\
        );

    \I__2665\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23282\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__23285\,
            I => \button_debounce_counterZ0Z_11\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__23282\,
            I => \button_debounce_counterZ0Z_11\
        );

    \I__2662\ : InMux
    port map (
            O => \N__23277\,
            I => un1_button_debounce_counter_cry_10
        );

    \I__2661\ : InMux
    port map (
            O => \N__23274\,
            I => \N__23270\
        );

    \I__2660\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23267\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__23270\,
            I => \button_debounce_counterZ0Z_12\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__23267\,
            I => \button_debounce_counterZ0Z_12\
        );

    \I__2657\ : InMux
    port map (
            O => \N__23262\,
            I => un1_button_debounce_counter_cry_11
        );

    \I__2656\ : InMux
    port map (
            O => \N__23259\,
            I => \sCounter_cry_18\
        );

    \I__2655\ : InMux
    port map (
            O => \N__23256\,
            I => \sCounter_cry_19\
        );

    \I__2654\ : InMux
    port map (
            O => \N__23253\,
            I => \sCounter_cry_20\
        );

    \I__2653\ : InMux
    port map (
            O => \N__23250\,
            I => \sCounter_cry_21\
        );

    \I__2652\ : InMux
    port map (
            O => \N__23247\,
            I => \N__23231\
        );

    \I__2651\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23231\
        );

    \I__2650\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23231\
        );

    \I__2649\ : InMux
    port map (
            O => \N__23244\,
            I => \N__23231\
        );

    \I__2648\ : InMux
    port map (
            O => \N__23243\,
            I => \N__23206\
        );

    \I__2647\ : InMux
    port map (
            O => \N__23242\,
            I => \N__23206\
        );

    \I__2646\ : InMux
    port map (
            O => \N__23241\,
            I => \N__23206\
        );

    \I__2645\ : InMux
    port map (
            O => \N__23240\,
            I => \N__23206\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__23231\,
            I => \N__23203\
        );

    \I__2643\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23194\
        );

    \I__2642\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23194\
        );

    \I__2641\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23194\
        );

    \I__2640\ : InMux
    port map (
            O => \N__23227\,
            I => \N__23194\
        );

    \I__2639\ : InMux
    port map (
            O => \N__23226\,
            I => \N__23185\
        );

    \I__2638\ : InMux
    port map (
            O => \N__23225\,
            I => \N__23185\
        );

    \I__2637\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23185\
        );

    \I__2636\ : InMux
    port map (
            O => \N__23223\,
            I => \N__23185\
        );

    \I__2635\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23176\
        );

    \I__2634\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23176\
        );

    \I__2633\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23176\
        );

    \I__2632\ : InMux
    port map (
            O => \N__23219\,
            I => \N__23176\
        );

    \I__2631\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23167\
        );

    \I__2630\ : InMux
    port map (
            O => \N__23217\,
            I => \N__23167\
        );

    \I__2629\ : InMux
    port map (
            O => \N__23216\,
            I => \N__23167\
        );

    \I__2628\ : InMux
    port map (
            O => \N__23215\,
            I => \N__23167\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__23206\,
            I => \LED_ACQ_c_i\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__23203\,
            I => \LED_ACQ_c_i\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__23194\,
            I => \LED_ACQ_c_i\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__23185\,
            I => \LED_ACQ_c_i\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__23176\,
            I => \LED_ACQ_c_i\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__23167\,
            I => \LED_ACQ_c_i\
        );

    \I__2621\ : InMux
    port map (
            O => \N__23154\,
            I => \sCounter_cry_22\
        );

    \I__2620\ : InMux
    port map (
            O => \N__23151\,
            I => un1_button_debounce_counter_cry_1
        );

    \I__2619\ : InMux
    port map (
            O => \N__23148\,
            I => un1_button_debounce_counter_cry_2
        );

    \I__2618\ : InMux
    port map (
            O => \N__23145\,
            I => un1_button_debounce_counter_cry_3
        );

    \I__2617\ : InMux
    port map (
            O => \N__23142\,
            I => \sCounter_cry_9\
        );

    \I__2616\ : InMux
    port map (
            O => \N__23139\,
            I => \sCounter_cry_10\
        );

    \I__2615\ : InMux
    port map (
            O => \N__23136\,
            I => \sCounter_cry_11\
        );

    \I__2614\ : InMux
    port map (
            O => \N__23133\,
            I => \sCounter_cry_12\
        );

    \I__2613\ : InMux
    port map (
            O => \N__23130\,
            I => \sCounter_cry_13\
        );

    \I__2612\ : InMux
    port map (
            O => \N__23127\,
            I => \sCounter_cry_14\
        );

    \I__2611\ : InMux
    port map (
            O => \N__23124\,
            I => \bfn_8_16_0_\
        );

    \I__2610\ : InMux
    port map (
            O => \N__23121\,
            I => \sCounter_cry_16\
        );

    \I__2609\ : InMux
    port map (
            O => \N__23118\,
            I => \sCounter_cry_17\
        );

    \I__2608\ : InMux
    port map (
            O => \N__23115\,
            I => \sCounter_cry_0\
        );

    \I__2607\ : InMux
    port map (
            O => \N__23112\,
            I => \sCounter_cry_1\
        );

    \I__2606\ : InMux
    port map (
            O => \N__23109\,
            I => \sCounter_cry_2\
        );

    \I__2605\ : InMux
    port map (
            O => \N__23106\,
            I => \sCounter_cry_3\
        );

    \I__2604\ : InMux
    port map (
            O => \N__23103\,
            I => \sCounter_cry_4\
        );

    \I__2603\ : InMux
    port map (
            O => \N__23100\,
            I => \sCounter_cry_5\
        );

    \I__2602\ : InMux
    port map (
            O => \N__23097\,
            I => \sCounter_cry_6\
        );

    \I__2601\ : InMux
    port map (
            O => \N__23094\,
            I => \bfn_8_15_0_\
        );

    \I__2600\ : InMux
    port map (
            O => \N__23091\,
            I => \sCounter_cry_8\
        );

    \I__2599\ : InMux
    port map (
            O => \N__23088\,
            I => \N__23085\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__23085\,
            I => \sEEPeriodZ0Z_20\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__23082\,
            I => \N__23079\
        );

    \I__2596\ : InMux
    port map (
            O => \N__23079\,
            I => \N__23076\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__23076\,
            I => \sEEPeriod_i_20\
        );

    \I__2594\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23070\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__23070\,
            I => \sEEPeriodZ0Z_21\
        );

    \I__2592\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23064\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__23064\,
            I => \sEEPeriod_i_21\
        );

    \I__2590\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23058\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__23058\,
            I => \sEEPeriodZ0Z_22\
        );

    \I__2588\ : InMux
    port map (
            O => \N__23055\,
            I => \N__23052\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__23052\,
            I => \sEEPeriod_i_22\
        );

    \I__2586\ : InMux
    port map (
            O => \N__23049\,
            I => \N__23046\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__23046\,
            I => \sEEPeriodZ0Z_23\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__23043\,
            I => \N__23040\
        );

    \I__2583\ : InMux
    port map (
            O => \N__23040\,
            I => \N__23037\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__23037\,
            I => \sEEPeriod_i_23\
        );

    \I__2581\ : InMux
    port map (
            O => \N__23034\,
            I => \bfn_8_13_0_\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__23031\,
            I => \N__23028\
        );

    \I__2579\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23025\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__23025\,
            I => un1_reset_rpi_inv_2_i_o3_15
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__23022\,
            I => \N__23019\
        );

    \I__2576\ : InMux
    port map (
            O => \N__23019\,
            I => \N__23016\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__23016\,
            I => un1_reset_rpi_inv_2_i_o3_11
        );

    \I__2574\ : InMux
    port map (
            O => \N__23013\,
            I => \N__23010\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__23010\,
            I => \sbuttonModeStatus_0_sqmuxa_17\
        );

    \I__2572\ : InMux
    port map (
            O => \N__23007\,
            I => \bfn_8_14_0_\
        );

    \I__2571\ : CascadeMux
    port map (
            O => \N__23004\,
            I => \N__23001\
        );

    \I__2570\ : InMux
    port map (
            O => \N__23001\,
            I => \N__22998\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__22998\,
            I => \sEEPeriod_i_12\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__22995\,
            I => \N__22992\
        );

    \I__2567\ : InMux
    port map (
            O => \N__22992\,
            I => \N__22989\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__22989\,
            I => \sEEPeriod_i_13\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__22986\,
            I => \N__22983\
        );

    \I__2564\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22980\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__22980\,
            I => \sEEPeriod_i_14\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__22977\,
            I => \N__22974\
        );

    \I__2561\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22971\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__22971\,
            I => \sEEPeriod_i_15\
        );

    \I__2559\ : InMux
    port map (
            O => \N__22968\,
            I => \N__22965\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__22965\,
            I => \sEEPeriodZ0Z_16\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__22962\,
            I => \N__22959\
        );

    \I__2556\ : InMux
    port map (
            O => \N__22959\,
            I => \N__22956\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__22956\,
            I => \sEEPeriod_i_16\
        );

    \I__2554\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22950\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__22950\,
            I => \sEEPeriodZ0Z_17\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__22947\,
            I => \N__22944\
        );

    \I__2551\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22941\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__22941\,
            I => \sEEPeriod_i_17\
        );

    \I__2549\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22935\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__22935\,
            I => \sEEPeriodZ0Z_18\
        );

    \I__2547\ : CascadeMux
    port map (
            O => \N__22932\,
            I => \N__22929\
        );

    \I__2546\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22926\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__22926\,
            I => \sEEPeriod_i_18\
        );

    \I__2544\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22920\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__22920\,
            I => \sEEPeriodZ0Z_19\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__22917\,
            I => \N__22914\
        );

    \I__2541\ : InMux
    port map (
            O => \N__22914\,
            I => \N__22911\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__22911\,
            I => \sEEPeriod_i_19\
        );

    \I__2539\ : InMux
    port map (
            O => \N__22908\,
            I => \N__22905\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__22905\,
            I => \sEEPeriodZ0Z_4\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__22902\,
            I => \N__22899\
        );

    \I__2536\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22896\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__22896\,
            I => \sEEPeriod_i_4\
        );

    \I__2534\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22890\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__22890\,
            I => \sEEPeriodZ0Z_5\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__22887\,
            I => \N__22884\
        );

    \I__2531\ : InMux
    port map (
            O => \N__22884\,
            I => \N__22881\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__22881\,
            I => \sEEPeriod_i_5\
        );

    \I__2529\ : InMux
    port map (
            O => \N__22878\,
            I => \N__22875\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__22875\,
            I => \sEEPeriodZ0Z_6\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__22872\,
            I => \N__22869\
        );

    \I__2526\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22866\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__22866\,
            I => \sEEPeriod_i_6\
        );

    \I__2524\ : InMux
    port map (
            O => \N__22863\,
            I => \N__22860\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__22860\,
            I => \sEEPeriodZ0Z_7\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__22857\,
            I => \N__22854\
        );

    \I__2521\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22851\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__22851\,
            I => \sEEPeriod_i_7\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__22848\,
            I => \N__22845\
        );

    \I__2518\ : InMux
    port map (
            O => \N__22845\,
            I => \N__22842\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__22842\,
            I => \sEEPeriod_i_8\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__22839\,
            I => \N__22836\
        );

    \I__2515\ : InMux
    port map (
            O => \N__22836\,
            I => \N__22833\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__22833\,
            I => \sEEPeriod_i_9\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__22830\,
            I => \N__22827\
        );

    \I__2512\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22824\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__22824\,
            I => \sEEPeriod_i_10\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__22821\,
            I => \N__22818\
        );

    \I__2509\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22815\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__22815\,
            I => \sEEPeriod_i_11\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__22812\,
            I => \g2_0_0_cascade_\
        );

    \I__2506\ : InMux
    port map (
            O => \N__22809\,
            I => \N__22806\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__22806\,
            I => \N__22803\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__22803\,
            I => g1_0_0_0
        );

    \I__2503\ : InMux
    port map (
            O => \N__22800\,
            I => \N__22797\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__22797\,
            I => g1_0_1
        );

    \I__2501\ : InMux
    port map (
            O => \N__22794\,
            I => \N__22791\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__22791\,
            I => \N__22788\
        );

    \I__2499\ : Span4Mux_v
    port map (
            O => \N__22788\,
            I => \N__22785\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__22785\,
            I => g0_2_0
        );

    \I__2497\ : InMux
    port map (
            O => \N__22782\,
            I => \N__22779\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__22779\,
            I => g1_4
        );

    \I__2495\ : CascadeMux
    port map (
            O => \N__22776\,
            I => \g2_0_cascade_\
        );

    \I__2494\ : InMux
    port map (
            O => \N__22773\,
            I => \N__22770\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__22770\,
            I => \sEEPeriodZ0Z_0\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__22767\,
            I => \N__22764\
        );

    \I__2491\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22761\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__22761\,
            I => \sEEPeriod_i_0\
        );

    \I__2489\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22755\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__22755\,
            I => \sEEPeriodZ0Z_1\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__22752\,
            I => \N__22749\
        );

    \I__2486\ : InMux
    port map (
            O => \N__22749\,
            I => \N__22746\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__22746\,
            I => \sEEPeriod_i_1\
        );

    \I__2484\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22740\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__22740\,
            I => \sEEPeriodZ0Z_2\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__22737\,
            I => \N__22734\
        );

    \I__2481\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22731\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__22731\,
            I => \sEEPeriod_i_2\
        );

    \I__2479\ : InMux
    port map (
            O => \N__22728\,
            I => \N__22725\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__22725\,
            I => \sEEPeriodZ0Z_3\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__22722\,
            I => \N__22719\
        );

    \I__2476\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22716\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__22716\,
            I => \sEEPeriod_i_3\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__22713\,
            I => \N__22710\
        );

    \I__2473\ : InMux
    port map (
            O => \N__22710\,
            I => \N__22707\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__22707\,
            I => g0_2_0_2
        );

    \I__2471\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22701\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__22701\,
            I => \N__22698\
        );

    \I__2469\ : Span4Mux_v
    port map (
            O => \N__22698\,
            I => \N__22695\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__22695\,
            I => g1_1
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__22692\,
            I => \g2_0_2_cascade_\
        );

    \I__2466\ : InMux
    port map (
            O => \N__22689\,
            I => \N__22686\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__22686\,
            I => g1_0_3
        );

    \I__2464\ : InMux
    port map (
            O => \N__22683\,
            I => \N__22680\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__22680\,
            I => g0_2_0_1
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__22677\,
            I => \g2_0_1_cascade_\
        );

    \I__2461\ : InMux
    port map (
            O => \N__22674\,
            I => \N__22671\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__22671\,
            I => \N__22668\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__22668\,
            I => g1_2
        );

    \I__2458\ : InMux
    port map (
            O => \N__22665\,
            I => \N__22662\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__22662\,
            I => g1_0_0_1
        );

    \I__2456\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22656\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__22656\,
            I => g1_0_2
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__22653\,
            I => \N__22650\
        );

    \I__2453\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22647\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__22647\,
            I => \N__22644\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__22644\,
            I => g0_2_0_0
        );

    \I__2450\ : InMux
    port map (
            O => \N__22641\,
            I => \N__22631\
        );

    \I__2449\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22631\
        );

    \I__2448\ : InMux
    port map (
            O => \N__22639\,
            I => \N__22624\
        );

    \I__2447\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22619\
        );

    \I__2446\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22619\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__22636\,
            I => \N__22614\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__22631\,
            I => \N__22611\
        );

    \I__2443\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22606\
        );

    \I__2442\ : InMux
    port map (
            O => \N__22629\,
            I => \N__22606\
        );

    \I__2441\ : InMux
    port map (
            O => \N__22628\,
            I => \N__22601\
        );

    \I__2440\ : InMux
    port map (
            O => \N__22627\,
            I => \N__22601\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__22624\,
            I => \N__22598\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__22619\,
            I => \N__22595\
        );

    \I__2437\ : InMux
    port map (
            O => \N__22618\,
            I => \N__22590\
        );

    \I__2436\ : InMux
    port map (
            O => \N__22617\,
            I => \N__22590\
        );

    \I__2435\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22587\
        );

    \I__2434\ : Span4Mux_v
    port map (
            O => \N__22611\,
            I => \N__22576\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__22606\,
            I => \N__22576\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22576\
        );

    \I__2431\ : Span4Mux_h
    port map (
            O => \N__22598\,
            I => \N__22576\
        );

    \I__2430\ : Span4Mux_h
    port map (
            O => \N__22595\,
            I => \N__22576\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__22590\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__22587\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__2427\ : Odrv4
    port map (
            O => \N__22576\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\
        );

    \I__2426\ : InMux
    port map (
            O => \N__22569\,
            I => \N__22566\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__22566\,
            I => \N__22563\
        );

    \I__2424\ : Span4Mux_v
    port map (
            O => \N__22563\,
            I => \N__22560\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__22560\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12\
        );

    \I__2422\ : InMux
    port map (
            O => \N__22557\,
            I => \N__22548\
        );

    \I__2421\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22548\
        );

    \I__2420\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22548\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__22548\,
            I => \spi_master_inst.sclk_gen_u0.N_150_0\
        );

    \I__2418\ : InMux
    port map (
            O => \N__22545\,
            I => \N__22542\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__22542\,
            I => \N__22539\
        );

    \I__2416\ : Odrv4
    port map (
            O => \N__22539\,
            I => \spi_master_inst.sclk_gen_u0.N_36\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__22536\,
            I => \N__22533\
        );

    \I__2414\ : InMux
    port map (
            O => \N__22533\,
            I => \N__22526\
        );

    \I__2413\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22526\
        );

    \I__2412\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22523\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__22526\,
            I => \N__22520\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__22523\,
            I => \N__22517\
        );

    \I__2409\ : Span4Mux_v
    port map (
            O => \N__22520\,
            I => \N__22514\
        );

    \I__2408\ : Span4Mux_h
    port map (
            O => \N__22517\,
            I => \N__22510\
        );

    \I__2407\ : Span4Mux_h
    port map (
            O => \N__22514\,
            I => \N__22507\
        );

    \I__2406\ : InMux
    port map (
            O => \N__22513\,
            I => \N__22504\
        );

    \I__2405\ : Span4Mux_h
    port map (
            O => \N__22510\,
            I => \N__22501\
        );

    \I__2404\ : Odrv4
    port map (
            O => \N__22507\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__22504\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__22501\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0\
        );

    \I__2401\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22487\
        );

    \I__2400\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22487\
        );

    \I__2399\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22484\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__22487\,
            I => \N__22480\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22477\
        );

    \I__2396\ : InMux
    port map (
            O => \N__22483\,
            I => \N__22474\
        );

    \I__2395\ : Span4Mux_v
    port map (
            O => \N__22480\,
            I => \N__22469\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__22477\,
            I => \N__22469\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__22474\,
            I => \spi_master_inst.sclk_gen_u0.div_clk_iZ0\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__22469\,
            I => \spi_master_inst.sclk_gen_u0.div_clk_iZ0\
        );

    \I__2391\ : InMux
    port map (
            O => \N__22464\,
            I => \N__22461\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__22461\,
            I => \spi_master_inst.sclk_gen_u0.delay_clk_iZ0\
        );

    \I__2389\ : InMux
    port map (
            O => \N__22458\,
            I => \N__22455\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__22455\,
            I => \N__22452\
        );

    \I__2387\ : Span4Mux_v
    port map (
            O => \N__22452\,
            I => \N__22449\
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__22449\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14\
        );

    \I__2385\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22443\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__22443\,
            I => \N__22440\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__22440\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0\
        );

    \I__2382\ : InMux
    port map (
            O => \N__22437\,
            I => \N__22434\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__22434\,
            I => \N__22431\
        );

    \I__2380\ : Odrv4
    port map (
            O => \N__22431\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8\
        );

    \I__2379\ : InMux
    port map (
            O => \N__22428\,
            I => \N__22425\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__22425\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9\
        );

    \I__2377\ : InMux
    port map (
            O => \N__22422\,
            I => \N__22419\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__22419\,
            I => \N__22416\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__22416\,
            I => \N__22413\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__22413\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7\
        );

    \I__2373\ : InMux
    port map (
            O => \N__22410\,
            I => \N__22407\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__22407\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1\
        );

    \I__2371\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22401\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__22401\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13\
        );

    \I__2369\ : InMux
    port map (
            O => \N__22398\,
            I => \N__22395\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__22395\,
            I => \N__22392\
        );

    \I__2367\ : Span4Mux_h
    port map (
            O => \N__22392\,
            I => \N__22389\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__22389\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10\
        );

    \I__2365\ : InMux
    port map (
            O => \N__22386\,
            I => \sCounterRAM_cry_4\
        );

    \I__2364\ : InMux
    port map (
            O => \N__22383\,
            I => \sCounterRAM_cry_5\
        );

    \I__2363\ : InMux
    port map (
            O => \N__22380\,
            I => \N__22364\
        );

    \I__2362\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22364\
        );

    \I__2361\ : InMux
    port map (
            O => \N__22378\,
            I => \N__22364\
        );

    \I__2360\ : InMux
    port map (
            O => \N__22377\,
            I => \N__22364\
        );

    \I__2359\ : InMux
    port map (
            O => \N__22376\,
            I => \N__22355\
        );

    \I__2358\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22355\
        );

    \I__2357\ : InMux
    port map (
            O => \N__22374\,
            I => \N__22355\
        );

    \I__2356\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22355\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__22364\,
            I => \un1_spi_data_miso_0_sqmuxa_1_i_0_N_3_0\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__22355\,
            I => \un1_spi_data_miso_0_sqmuxa_1_i_0_N_3_0\
        );

    \I__2353\ : InMux
    port map (
            O => \N__22350\,
            I => \sCounterRAM_cry_6\
        );

    \I__2352\ : InMux
    port map (
            O => \N__22347\,
            I => \N__22344\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__22344\,
            I => \sSPI_MSB0LSB1_RNIO3VPZ0Z1\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__22341\,
            I => \N__22338\
        );

    \I__2349\ : InMux
    port map (
            O => \N__22338\,
            I => \N__22335\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__22335\,
            I => \N__22332\
        );

    \I__2347\ : Span4Mux_v
    port map (
            O => \N__22332\,
            I => \N__22329\
        );

    \I__2346\ : Span4Mux_h
    port map (
            O => \N__22329\,
            I => \N__22326\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__22326\,
            I => \sbuttonModeStatus_0_sqmuxa_16\
        );

    \I__2344\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22320\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__22320\,
            I => \N__22317\
        );

    \I__2342\ : Span4Mux_v
    port map (
            O => \N__22317\,
            I => \N__22314\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__22314\,
            I => \sbuttonModeStatus_0_sqmuxa_14\
        );

    \I__2340\ : InMux
    port map (
            O => \N__22311\,
            I => \N__22308\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__22308\,
            I => \N__22305\
        );

    \I__2338\ : Sp12to4
    port map (
            O => \N__22305\,
            I => \N__22302\
        );

    \I__2337\ : Odrv12
    port map (
            O => \N__22302\,
            I => \sbuttonModeStatus_0_sqmuxa_15\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__22299\,
            I => \op_gt_op_gt_un13_striginternallto23_11_cascade_\
        );

    \I__2335\ : InMux
    port map (
            O => \N__22296\,
            I => \N__22293\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__22293\,
            I => op_gt_op_gt_un13_striginternallto23_16
        );

    \I__2333\ : InMux
    port map (
            O => \N__22290\,
            I => \N__22284\
        );

    \I__2332\ : InMux
    port map (
            O => \N__22289\,
            I => \N__22284\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__22284\,
            I => \N__22281\
        );

    \I__2330\ : Span4Mux_v
    port map (
            O => \N__22281\,
            I => \N__22277\
        );

    \I__2329\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22274\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__22277\,
            I => \sTrigInternalZ0\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__22274\,
            I => \sTrigInternalZ0\
        );

    \I__2326\ : CascadeMux
    port map (
            O => \N__22269\,
            I => \N__22266\
        );

    \I__2325\ : InMux
    port map (
            O => \N__22266\,
            I => \N__22263\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__22263\,
            I => op_gt_op_gt_un13_striginternal_0
        );

    \I__2323\ : IoInMux
    port map (
            O => \N__22260\,
            I => \N__22257\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__22257\,
            I => \N__22254\
        );

    \I__2321\ : IoSpan4Mux
    port map (
            O => \N__22254\,
            I => \N__22251\
        );

    \I__2320\ : Span4Mux_s2_h
    port map (
            O => \N__22251\,
            I => \N__22248\
        );

    \I__2319\ : Sp12to4
    port map (
            O => \N__22248\,
            I => \N__22245\
        );

    \I__2318\ : Span12Mux_s11_v
    port map (
            O => \N__22245\,
            I => \N__22242\
        );

    \I__2317\ : Odrv12
    port map (
            O => \N__22242\,
            I => \LED_ACQ_obuf_RNOZ0\
        );

    \I__2316\ : InMux
    port map (
            O => \N__22239\,
            I => \N__22236\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__22236\,
            I => op_gt_op_gt_un13_striginternallto23_18
        );

    \I__2314\ : InMux
    port map (
            O => \N__22233\,
            I => \bfn_7_16_0_\
        );

    \I__2313\ : InMux
    port map (
            O => \N__22230\,
            I => \sCounterRAM_cry_0\
        );

    \I__2312\ : InMux
    port map (
            O => \N__22227\,
            I => \sCounterRAM_cry_1\
        );

    \I__2311\ : InMux
    port map (
            O => \N__22224\,
            I => \sCounterRAM_cry_2\
        );

    \I__2310\ : InMux
    port map (
            O => \N__22221\,
            I => \sCounterRAM_cry_3\
        );

    \I__2309\ : CascadeMux
    port map (
            O => \N__22218\,
            I => \sbuttonModeStatus_0_sqmuxa_22_cascade_\
        );

    \I__2308\ : InMux
    port map (
            O => \N__22215\,
            I => \N__22212\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__22212\,
            I => \N__22209\
        );

    \I__2306\ : Span4Mux_v
    port map (
            O => \N__22209\,
            I => \N__22206\
        );

    \I__2305\ : Span4Mux_v
    port map (
            O => \N__22206\,
            I => \N__22202\
        );

    \I__2304\ : InMux
    port map (
            O => \N__22205\,
            I => \N__22199\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__22202\,
            I => \sbuttonModeStatusZ0\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__22199\,
            I => \sbuttonModeStatusZ0\
        );

    \I__2301\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22191\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__22191\,
            I => \N__22188\
        );

    \I__2299\ : Odrv12
    port map (
            O => \N__22188\,
            I => g1_0_0_3
        );

    \I__2298\ : InMux
    port map (
            O => \N__22185\,
            I => \N__22182\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__22182\,
            I => un1_reset_rpi_inv_2_i_o3_16
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__22179\,
            I => \N__22176\
        );

    \I__2295\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22173\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__22173\,
            I => \N__22170\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__22170\,
            I => g0_2_0_4
        );

    \I__2292\ : InMux
    port map (
            O => \N__22167\,
            I => \N__22164\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__22164\,
            I => g2_0_4
        );

    \I__2290\ : InMux
    port map (
            O => \N__22161\,
            I => \N__22158\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__22158\,
            I => g2_0_3
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__22155\,
            I => \g1_0_1_1_cascade_\
        );

    \I__2287\ : InMux
    port map (
            O => \N__22152\,
            I => \N__22149\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__22149\,
            I => g1_0_4
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__22146\,
            I => \N__22143\
        );

    \I__2284\ : InMux
    port map (
            O => \N__22143\,
            I => \N__22140\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__22140\,
            I => op_gt_op_gt_un13_striginternallto23_13
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__22137\,
            I => \op_gt_op_gt_un13_striginternal_0_cascade_\
        );

    \I__2281\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22130\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__22133\,
            I => \N__22127\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__22130\,
            I => \N__22124\
        );

    \I__2278\ : InMux
    port map (
            O => \N__22127\,
            I => \N__22121\
        );

    \I__2277\ : Span4Mux_v
    port map (
            O => \N__22124\,
            I => \N__22118\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__22121\,
            I => \N__22115\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__22118\,
            I => un3_trig_0_4
        );

    \I__2274\ : Odrv12
    port map (
            O => \N__22115\,
            I => un3_trig_0_4
        );

    \I__2273\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22107\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__22107\,
            I => \N__22104\
        );

    \I__2271\ : Odrv12
    port map (
            O => \N__22104\,
            I => un1_reset_rpi_inv_2_i_o3_8
        );

    \I__2270\ : CascadeMux
    port map (
            O => \N__22101\,
            I => \un1_reset_rpi_inv_2_i_o3_18_cascade_\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__22098\,
            I => \N__22095\
        );

    \I__2268\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22092\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__22092\,
            I => \N__22088\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__22091\,
            I => \N__22085\
        );

    \I__2265\ : Span4Mux_v
    port map (
            O => \N__22088\,
            I => \N__22082\
        );

    \I__2264\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22079\
        );

    \I__2263\ : Span4Mux_h
    port map (
            O => \N__22082\,
            I => \N__22076\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__22079\,
            I => \N__22073\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__22076\,
            I => un3_trig_0_5
        );

    \I__2260\ : Odrv12
    port map (
            O => \N__22073\,
            I => un3_trig_0_5
        );

    \I__2259\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22065\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__22065\,
            I => un1_reset_rpi_inv_2_i_o3_13
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__22062\,
            I => \N__22059\
        );

    \I__2256\ : InMux
    port map (
            O => \N__22059\,
            I => \N__22056\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__22056\,
            I => g0_2_0_3
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__22053\,
            I => \sTrigInternal_RNIOMLDZ0Z1_cascade_\
        );

    \I__2253\ : InMux
    port map (
            O => \N__22050\,
            I => \N__22047\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__22047\,
            I => \sTrigInternal_RNIOMLDZ0Z1\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__22044\,
            I => \sTrigInternal_RNOZ0Z_0_cascade_\
        );

    \I__2250\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22037\
        );

    \I__2249\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22034\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__22037\,
            I => \N__22029\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__22034\,
            I => \N__22029\
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__22029\,
            I => un3_trig_0
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__22026\,
            I => \sEETrigInternal_prev_RNISEUGZ0_cascade_\
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__22023\,
            I => \N__22019\
        );

    \I__2243\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22014\
        );

    \I__2242\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22014\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__22014\,
            I => \N__22011\
        );

    \I__2240\ : Odrv12
    port map (
            O => \N__22011\,
            I => un3_trig_0_2
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__22008\,
            I => \N__22004\
        );

    \I__2238\ : InMux
    port map (
            O => \N__22007\,
            I => \N__21999\
        );

    \I__2237\ : InMux
    port map (
            O => \N__22004\,
            I => \N__21999\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__21999\,
            I => \N__21996\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__21996\,
            I => un3_trig_0_1
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__21993\,
            I => \g1_3_cascade_\
        );

    \I__2233\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21987\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__21987\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13\
        );

    \I__2231\ : InMux
    port map (
            O => \N__21984\,
            I => \N__21981\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__21981\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1\
        );

    \I__2229\ : InMux
    port map (
            O => \N__21978\,
            I => \N__21975\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__21975\,
            I => \N__21972\
        );

    \I__2227\ : Span4Mux_h
    port map (
            O => \N__21972\,
            I => \N__21969\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__21969\,
            I => \sEESingleContZ0\
        );

    \I__2225\ : InMux
    port map (
            O => \N__21966\,
            I => \N__21961\
        );

    \I__2224\ : InMux
    port map (
            O => \N__21965\,
            I => \N__21956\
        );

    \I__2223\ : InMux
    port map (
            O => \N__21964\,
            I => \N__21956\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__21961\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__21956\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3\
        );

    \I__2220\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21943\
        );

    \I__2219\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21943\
        );

    \I__2218\ : InMux
    port map (
            O => \N__21949\,
            I => \N__21940\
        );

    \I__2217\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21937\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__21943\,
            I => \spi_master_inst.sclk_gen_u0.N_1515\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__21940\,
            I => \spi_master_inst.sclk_gen_u0.N_1515\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__21937\,
            I => \spi_master_inst.sclk_gen_u0.N_1515\
        );

    \I__2213\ : CEMux
    port map (
            O => \N__21930\,
            I => \N__21927\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__21927\,
            I => \N__21924\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__21924\,
            I => \sEESingleCont_1_sqmuxa\
        );

    \I__2210\ : InMux
    port map (
            O => \N__21921\,
            I => \bfn_6_14_0_\
        );

    \I__2209\ : IoInMux
    port map (
            O => \N__21918\,
            I => \N__21915\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__21915\,
            I => \N__21912\
        );

    \I__2207\ : Span4Mux_s1_h
    port map (
            O => \N__21912\,
            I => \N__21909\
        );

    \I__2206\ : Span4Mux_h
    port map (
            O => \N__21909\,
            I => \N__21906\
        );

    \I__2205\ : Span4Mux_h
    port map (
            O => \N__21906\,
            I => \N__21903\
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__21903\,
            I => \pon_obuf_RNOZ0\
        );

    \I__2203\ : InMux
    port map (
            O => \N__21900\,
            I => \N__21897\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__21897\,
            I => \N__21894\
        );

    \I__2201\ : Odrv12
    port map (
            O => \N__21894\,
            I => g1_0_5
        );

    \I__2200\ : InMux
    port map (
            O => \N__21891\,
            I => \N__21888\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__21888\,
            I => g1
        );

    \I__2198\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21882\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__21882\,
            I => \sEEPon_i_1\
        );

    \I__2196\ : InMux
    port map (
            O => \N__21879\,
            I => \N__21876\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21873\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__21873\,
            I => \sEEPonZ0Z_2\
        );

    \I__2193\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21867\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__21867\,
            I => \sEEPon_i_2\
        );

    \I__2191\ : InMux
    port map (
            O => \N__21864\,
            I => \N__21861\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__21861\,
            I => \N__21858\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__21858\,
            I => \sEEPonZ0Z_3\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__21855\,
            I => \N__21852\
        );

    \I__2187\ : InMux
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__21849\,
            I => \sEEPon_i_3\
        );

    \I__2185\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21843\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__21843\,
            I => \N__21840\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__21840\,
            I => \sEEPonZ0Z_4\
        );

    \I__2182\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21834\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__21834\,
            I => \sEEPon_i_4\
        );

    \I__2180\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21828\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__21828\,
            I => \N__21825\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__21825\,
            I => \sEEPonZ0Z_5\
        );

    \I__2177\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21819\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__21819\,
            I => \sEEPon_i_5\
        );

    \I__2175\ : InMux
    port map (
            O => \N__21816\,
            I => \N__21813\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__21813\,
            I => \N__21810\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__21810\,
            I => \N__21807\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__21807\,
            I => \sEEPonZ0Z_6\
        );

    \I__2171\ : InMux
    port map (
            O => \N__21804\,
            I => \N__21801\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__21801\,
            I => \sEEPon_i_6\
        );

    \I__2169\ : InMux
    port map (
            O => \N__21798\,
            I => \N__21795\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__21795\,
            I => \N__21792\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__21792\,
            I => \sEEPonZ0Z_7\
        );

    \I__2166\ : InMux
    port map (
            O => \N__21789\,
            I => \N__21786\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__21786\,
            I => \sEEPon_i_7\
        );

    \I__2164\ : InMux
    port map (
            O => \N__21783\,
            I => \N__21780\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__21780\,
            I => \sEEPonPoffZ0Z_1\
        );

    \I__2162\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21774\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__21774\,
            I => \sEEPonPoffZ0Z_2\
        );

    \I__2160\ : InMux
    port map (
            O => \N__21771\,
            I => \N__21768\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__21768\,
            I => \sEEPonPoffZ0Z_3\
        );

    \I__2158\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21762\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__21762\,
            I => \sEEPonPoffZ0Z_4\
        );

    \I__2156\ : InMux
    port map (
            O => \N__21759\,
            I => \N__21756\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__21756\,
            I => \sEEPonPoffZ0Z_5\
        );

    \I__2154\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21750\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__21750\,
            I => \sEEPonPoffZ0Z_6\
        );

    \I__2152\ : InMux
    port map (
            O => \N__21747\,
            I => \N__21744\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__21744\,
            I => \sEEPonPoffZ0Z_7\
        );

    \I__2150\ : InMux
    port map (
            O => \N__21741\,
            I => \N__21738\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__21738\,
            I => \N__21735\
        );

    \I__2148\ : Odrv12
    port map (
            O => \N__21735\,
            I => \sEEPonZ0Z_0\
        );

    \I__2147\ : InMux
    port map (
            O => \N__21732\,
            I => \N__21729\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__21729\,
            I => \sEEPon_i_0\
        );

    \I__2145\ : InMux
    port map (
            O => \N__21726\,
            I => \N__21723\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__21723\,
            I => \N__21720\
        );

    \I__2143\ : Odrv12
    port map (
            O => \N__21720\,
            I => \sEEPonZ0Z_1\
        );

    \I__2142\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21714\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__21714\,
            I => \sEEPonPoffZ0Z_0\
        );

    \I__2140\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21708\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__21708\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11\
        );

    \I__2138\ : CascadeMux
    port map (
            O => \N__21705\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15_cascade_\
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__21702\,
            I => \N__21697\
        );

    \I__2136\ : InMux
    port map (
            O => \N__21701\,
            I => \N__21689\
        );

    \I__2135\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21686\
        );

    \I__2134\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21683\
        );

    \I__2133\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21680\
        );

    \I__2132\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21673\
        );

    \I__2131\ : InMux
    port map (
            O => \N__21694\,
            I => \N__21673\
        );

    \I__2130\ : InMux
    port map (
            O => \N__21693\,
            I => \N__21673\
        );

    \I__2129\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21670\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__21689\,
            I => \N__21667\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__21686\,
            I => \N__21662\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__21683\,
            I => \N__21662\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__21680\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__21673\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__21670\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__21667\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2121\ : Odrv12
    port map (
            O => \N__21662\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\
        );

    \I__2120\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21648\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__21648\,
            I => \N__21645\
        );

    \I__2118\ : Odrv4
    port map (
            O => \N__21645\,
            I => \spi_master_inst.spi_data_path_u1.N_1412\
        );

    \I__2117\ : InMux
    port map (
            O => \N__21642\,
            I => \N__21637\
        );

    \I__2116\ : InMux
    port map (
            O => \N__21641\,
            I => \N__21634\
        );

    \I__2115\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21631\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__21637\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__21634\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__21631\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3\
        );

    \I__2111\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21619\
        );

    \I__2110\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21616\
        );

    \I__2109\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21613\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__21619\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__21616\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__21613\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__21606\,
            I => \N__21602\
        );

    \I__2104\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21598\
        );

    \I__2103\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21595\
        );

    \I__2102\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21592\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__21598\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__21595\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__21592\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2\
        );

    \I__2098\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21581\
        );

    \I__2097\ : InMux
    port map (
            O => \N__21584\,
            I => \N__21578\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__21581\,
            I => \spi_master_inst.sclk_gen_u0.N_1666\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__21578\,
            I => \spi_master_inst.sclk_gen_u0.N_1666\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__21573\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3_cascade_\
        );

    \I__2093\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21565\
        );

    \I__2092\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21562\
        );

    \I__2091\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21559\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__21565\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__21562\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__21559\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__21552\,
            I => \spi_master_inst.sclk_gen_u0.N_1515_cascade_\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__21549\,
            I => \spi_master_inst.sclk_gen_u0.N_36_cascade_\
        );

    \I__2085\ : InMux
    port map (
            O => \N__21546\,
            I => \N__21543\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__21543\,
            I => \spi_master_inst.sclk_gen_u0.N_48\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__21540\,
            I => \spi_master_inst.sclk_gen_u0.N_5_cascade_\
        );

    \I__2082\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21533\
        );

    \I__2081\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21530\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__21533\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_start_iZ0\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__21530\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_start_iZ0\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__21525\,
            I => \N__21521\
        );

    \I__2077\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21517\
        );

    \I__2076\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21512\
        );

    \I__2075\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21512\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__21517\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__21512\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1\
        );

    \I__2072\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21504\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__21504\,
            I => \spi_master_inst.spi_data_path_u1.N_1415\
        );

    \I__2070\ : InMux
    port map (
            O => \N__21501\,
            I => \N__21498\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__21498\,
            I => \N__21495\
        );

    \I__2068\ : Span4Mux_h
    port map (
            O => \N__21495\,
            I => \N__21492\
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__21492\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__21489\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14_cascade_\
        );

    \I__2065\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21483\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__21483\,
            I => \spi_master_inst.spi_data_path_u1.N_1419\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__21480\,
            I => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_\
        );

    \I__2062\ : InMux
    port map (
            O => \N__21477\,
            I => \N__21474\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__21474\,
            I => \spi_master_inst.spi_data_path_u1.N_1422\
        );

    \I__2060\ : InMux
    port map (
            O => \N__21471\,
            I => \N__21465\
        );

    \I__2059\ : InMux
    port map (
            O => \N__21470\,
            I => \N__21465\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__21465\,
            I => \spi_master_inst.sclk_gen_u0.N_1520\
        );

    \I__2057\ : InMux
    port map (
            O => \N__21462\,
            I => \N__21444\
        );

    \I__2056\ : InMux
    port map (
            O => \N__21461\,
            I => \N__21444\
        );

    \I__2055\ : InMux
    port map (
            O => \N__21460\,
            I => \N__21444\
        );

    \I__2054\ : InMux
    port map (
            O => \N__21459\,
            I => \N__21444\
        );

    \I__2053\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21444\
        );

    \I__2052\ : InMux
    port map (
            O => \N__21457\,
            I => \N__21437\
        );

    \I__2051\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21437\
        );

    \I__2050\ : InMux
    port map (
            O => \N__21455\,
            I => \N__21437\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__21444\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_start_i_i\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__21437\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_start_i_i\
        );

    \I__2047\ : InMux
    port map (
            O => \N__21432\,
            I => \bfn_5_13_0_\
        );

    \I__2046\ : InMux
    port map (
            O => \N__21429\,
            I => \N__21426\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__21426\,
            I => \spi_master_inst.spi_data_path_u1.N_1423\
        );

    \I__2044\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21417\
        );

    \I__2043\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21417\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__21417\,
            I => \N__21413\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__21416\,
            I => \N__21410\
        );

    \I__2040\ : Span4Mux_v
    port map (
            O => \N__21413\,
            I => \N__21405\
        );

    \I__2039\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21402\
        );

    \I__2038\ : InMux
    port map (
            O => \N__21409\,
            I => \N__21399\
        );

    \I__2037\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21396\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__21405\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__21402\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__21399\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__21396\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__21387\,
            I => \N__21384\
        );

    \I__2031\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21381\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__21381\,
            I => \spi_master_inst.spi_data_path_u1.N_1416\
        );

    \I__2029\ : InMux
    port map (
            O => \N__21378\,
            I => \N__21375\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__21375\,
            I => \sEEPonPoff_i_0\
        );

    \I__2027\ : InMux
    port map (
            O => \N__21372\,
            I => \N__21369\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__21369\,
            I => \sEEPonPoff_i_1\
        );

    \I__2025\ : InMux
    port map (
            O => \N__21366\,
            I => \N__21363\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__21363\,
            I => \sEEPonPoff_i_2\
        );

    \I__2023\ : CascadeMux
    port map (
            O => \N__21360\,
            I => \N__21357\
        );

    \I__2022\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21354\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__21354\,
            I => \sEEPonPoff_i_3\
        );

    \I__2020\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21348\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__21348\,
            I => \sEEPonPoff_i_4\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__21345\,
            I => \N__21342\
        );

    \I__2017\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21339\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__21339\,
            I => \sEEPonPoff_i_5\
        );

    \I__2015\ : InMux
    port map (
            O => \N__21336\,
            I => \N__21333\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__21333\,
            I => \sEEPonPoff_i_6\
        );

    \I__2013\ : InMux
    port map (
            O => \N__21330\,
            I => \N__21327\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__21327\,
            I => \sEEPonPoff_i_7\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__21324\,
            I => \spi_master_inst.sclk_gen_u0.N_1666_cascade_\
        );

    \I__2010\ : InMux
    port map (
            O => \N__21321\,
            I => \N__21318\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__21318\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4\
        );

    \I__2008\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21309\
        );

    \I__2007\ : InMux
    port map (
            O => \N__21314\,
            I => \N__21309\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__21309\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__21306\,
            I => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__21303\,
            I => \spi_master_inst.sclk_gen_u0.N_48_cascade_\
        );

    \I__2003\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21293\
        );

    \I__2002\ : InMux
    port map (
            O => \N__21299\,
            I => \N__21290\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__21298\,
            I => \N__21287\
        );

    \I__2000\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21284\
        );

    \I__1999\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21281\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__21293\,
            I => \N__21278\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__21290\,
            I => \N__21275\
        );

    \I__1996\ : InMux
    port map (
            O => \N__21287\,
            I => \N__21272\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__21284\,
            I => \N__21265\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__21281\,
            I => \N__21265\
        );

    \I__1993\ : Span4Mux_h
    port map (
            O => \N__21278\,
            I => \N__21265\
        );

    \I__1992\ : Span4Mux_h
    port map (
            O => \N__21275\,
            I => \N__21262\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__21272\,
            I => \spi_master_inst.ss_start_i\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__21265\,
            I => \spi_master_inst.ss_start_i\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__21262\,
            I => \spi_master_inst.ss_start_i\
        );

    \I__1988\ : InMux
    port map (
            O => \N__21255\,
            I => \bfn_5_5_0_\
        );

    \I__1987\ : InMux
    port map (
            O => \N__21252\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_0\
        );

    \I__1986\ : InMux
    port map (
            O => \N__21249\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_1\
        );

    \I__1985\ : InMux
    port map (
            O => \N__21246\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_2\
        );

    \I__1984\ : InMux
    port map (
            O => \N__21243\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_3\
        );

    \I__1983\ : InMux
    port map (
            O => \N__21240\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_4\
        );

    \I__1982\ : InMux
    port map (
            O => \N__21237\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_5\
        );

    \I__1981\ : InMux
    port map (
            O => \N__21234\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_6\
        );

    \I__1980\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21227\
        );

    \I__1979\ : InMux
    port map (
            O => \N__21230\,
            I => \N__21224\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__21227\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__21224\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6\
        );

    \I__1976\ : InMux
    port map (
            O => \N__21219\,
            I => \N__21215\
        );

    \I__1975\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21212\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__21215\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__21212\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__21207\,
            I => \N__21203\
        );

    \I__1971\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21200\
        );

    \I__1970\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21197\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__21200\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__21197\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7\
        );

    \I__1967\ : InMux
    port map (
            O => \N__21192\,
            I => \N__21188\
        );

    \I__1966\ : InMux
    port map (
            O => \N__21191\,
            I => \N__21185\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__21188\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__21185\,
            I => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4\
        );

    \I__1963\ : InMux
    port map (
            O => \N__21180\,
            I => \N__21177\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__21177\,
            I => \N__21173\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__21176\,
            I => \N__21169\
        );

    \I__1960\ : Span4Mux_v
    port map (
            O => \N__21173\,
            I => \N__21165\
        );

    \I__1959\ : InMux
    port map (
            O => \N__21172\,
            I => \N__21162\
        );

    \I__1958\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21159\
        );

    \I__1957\ : InMux
    port map (
            O => \N__21168\,
            I => \N__21156\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__21165\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__21162\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__21159\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__21156\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0\
        );

    \I__1952\ : IoInMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__21144\,
            I => \N__21141\
        );

    \I__1950\ : Span4Mux_s0_v
    port map (
            O => \N__21141\,
            I => \N__21138\
        );

    \I__1949\ : Span4Mux_v
    port map (
            O => \N__21138\,
            I => \N__21135\
        );

    \I__1948\ : Span4Mux_v
    port map (
            O => \N__21135\,
            I => \N__21132\
        );

    \I__1947\ : Odrv4
    port map (
            O => \N__21132\,
            I => \DAC_mosi_c\
        );

    \I__1946\ : InMux
    port map (
            O => \N__21129\,
            I => \N__21126\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__21126\,
            I => \N__21123\
        );

    \I__1944\ : Span4Mux_h
    port map (
            O => \N__21123\,
            I => \N__21120\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__21120\,
            I => \spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1\
        );

    \I__1942\ : InMux
    port map (
            O => \N__21117\,
            I => \N__21114\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__21114\,
            I => \N__21111\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__21111\,
            I => \N__21106\
        );

    \I__1939\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21103\
        );

    \I__1938\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21100\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__21106\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__21103\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__21100\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5\
        );

    \I__1934\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21090\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__21090\,
            I => \N__21087\
        );

    \I__1932\ : Span4Mux_v
    port map (
            O => \N__21087\,
            I => \N__21082\
        );

    \I__1931\ : InMux
    port map (
            O => \N__21086\,
            I => \N__21079\
        );

    \I__1930\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21076\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__21082\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__21079\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__21076\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4\
        );

    \I__1926\ : IoInMux
    port map (
            O => \N__21069\,
            I => \N__21066\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__21066\,
            I => \N__21063\
        );

    \I__1924\ : Span4Mux_s1_v
    port map (
            O => \N__21063\,
            I => \N__21060\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__21060\,
            I => \N__21056\
        );

    \I__1922\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21053\
        );

    \I__1921\ : Span4Mux_v
    port map (
            O => \N__21056\,
            I => \N__21050\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__21053\,
            I => \N__21047\
        );

    \I__1919\ : Span4Mux_h
    port map (
            O => \N__21050\,
            I => \N__21042\
        );

    \I__1918\ : Span4Mux_v
    port map (
            O => \N__21047\,
            I => \N__21042\
        );

    \I__1917\ : Odrv4
    port map (
            O => \N__21042\,
            I => \DAC_sclk_c\
        );

    \I__1916\ : InMux
    port map (
            O => \N__21039\,
            I => \N__21036\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__21036\,
            I => \N__21033\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__21033\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO\
        );

    \I__1913\ : InMux
    port map (
            O => \N__21030\,
            I => \N__21023\
        );

    \I__1912\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21018\
        );

    \I__1911\ : InMux
    port map (
            O => \N__21028\,
            I => \N__21018\
        );

    \I__1910\ : InMux
    port map (
            O => \N__21027\,
            I => \N__21015\
        );

    \I__1909\ : InMux
    port map (
            O => \N__21026\,
            I => \N__21012\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__21023\,
            I => \N__21007\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__21018\,
            I => \N__21007\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__21015\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__21012\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__21007\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__21000\,
            I => \N__20996\
        );

    \I__1902\ : InMux
    port map (
            O => \N__20999\,
            I => \N__20987\
        );

    \I__1901\ : InMux
    port map (
            O => \N__20996\,
            I => \N__20987\
        );

    \I__1900\ : InMux
    port map (
            O => \N__20995\,
            I => \N__20987\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__20994\,
            I => \N__20981\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__20987\,
            I => \N__20978\
        );

    \I__1897\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20975\
        );

    \I__1896\ : CEMux
    port map (
            O => \N__20985\,
            I => \N__20972\
        );

    \I__1895\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20967\
        );

    \I__1894\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20967\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__20978\,
            I => \N__20964\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20961\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__20972\,
            I => \spi_master_inst.o_sclk_RNIH6AC\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__20967\,
            I => \spi_master_inst.o_sclk_RNIH6AC\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__20964\,
            I => \spi_master_inst.o_sclk_RNIH6AC\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__20961\,
            I => \spi_master_inst.o_sclk_RNIH6AC\
        );

    \I__1887\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20949\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__20949\,
            I => \N__20946\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__20946\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO\
        );

    \I__1884\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20940\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__20940\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO\
        );

    \I__1882\ : InMux
    port map (
            O => \N__20937\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0\
        );

    \I__1881\ : InMux
    port map (
            O => \N__20934\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1\
        );

    \I__1880\ : InMux
    port map (
            O => \N__20931\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2\
        );

    \I__1879\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20924\
        );

    \I__1878\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20921\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__20924\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__20921\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4\
        );

    \I__1875\ : InMux
    port map (
            O => \N__20916\,
            I => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3\
        );

    \I__1874\ : InMux
    port map (
            O => \N__20913\,
            I => \bfn_3_5_0_\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__20910\,
            I => \N__20906\
        );

    \I__1872\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20903\
        );

    \I__1871\ : InMux
    port map (
            O => \N__20906\,
            I => \N__20900\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__20903\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__20900\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5\
        );

    \I__1868\ : InMux
    port map (
            O => \N__20895\,
            I => \bfn_3_3_0_\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__20892\,
            I => \N__20889\
        );

    \I__1866\ : InMux
    port map (
            O => \N__20889\,
            I => \N__20885\
        );

    \I__1865\ : InMux
    port map (
            O => \N__20888\,
            I => \N__20882\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__20885\,
            I => \N__20879\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__20882\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1\
        );

    \I__1862\ : Odrv12
    port map (
            O => \N__20879\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1\
        );

    \I__1861\ : InMux
    port map (
            O => \N__20874\,
            I => \N__20871\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__20871\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_s_1\
        );

    \I__1859\ : InMux
    port map (
            O => \N__20868\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0\
        );

    \I__1858\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20860\
        );

    \I__1857\ : InMux
    port map (
            O => \N__20864\,
            I => \N__20857\
        );

    \I__1856\ : InMux
    port map (
            O => \N__20863\,
            I => \N__20854\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__20860\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__20857\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__20854\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2\
        );

    \I__1852\ : InMux
    port map (
            O => \N__20847\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__20844\,
            I => \N__20841\
        );

    \I__1850\ : InMux
    port map (
            O => \N__20841\,
            I => \N__20836\
        );

    \I__1849\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20833\
        );

    \I__1848\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20830\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__20836\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__20833\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__20830\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3\
        );

    \I__1844\ : InMux
    port map (
            O => \N__20823\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2\
        );

    \I__1843\ : InMux
    port map (
            O => \N__20820\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3\
        );

    \I__1842\ : InMux
    port map (
            O => \N__20817\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4\
        );

    \I__1841\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20809\
        );

    \I__1840\ : InMux
    port map (
            O => \N__20813\,
            I => \N__20806\
        );

    \I__1839\ : InMux
    port map (
            O => \N__20812\,
            I => \N__20803\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__20809\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__20806\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__20803\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6\
        );

    \I__1835\ : InMux
    port map (
            O => \N__20796\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5\
        );

    \I__1834\ : InMux
    port map (
            O => \N__20793\,
            I => \N__20779\
        );

    \I__1833\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20779\
        );

    \I__1832\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20779\
        );

    \I__1831\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20774\
        );

    \I__1830\ : InMux
    port map (
            O => \N__20789\,
            I => \N__20774\
        );

    \I__1829\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20767\
        );

    \I__1828\ : InMux
    port map (
            O => \N__20787\,
            I => \N__20767\
        );

    \I__1827\ : InMux
    port map (
            O => \N__20786\,
            I => \N__20767\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__20779\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__20774\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__20767\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i\
        );

    \I__1823\ : InMux
    port map (
            O => \N__20760\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__20757\,
            I => \N__20752\
        );

    \I__1821\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20749\
        );

    \I__1820\ : InMux
    port map (
            O => \N__20755\,
            I => \N__20746\
        );

    \I__1819\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20743\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__20749\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__20746\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__20743\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7\
        );

    \I__1815\ : InMux
    port map (
            O => \N__20736\,
            I => \N__20732\
        );

    \I__1814\ : InMux
    port map (
            O => \N__20735\,
            I => \N__20729\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__20732\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__20729\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2\
        );

    \I__1811\ : InMux
    port map (
            O => \N__20724\,
            I => \sRAM_pointer_read_cry_11\
        );

    \I__1810\ : InMux
    port map (
            O => \N__20721\,
            I => \sRAM_pointer_read_cry_12\
        );

    \I__1809\ : InMux
    port map (
            O => \N__20718\,
            I => \sRAM_pointer_read_cry_13\
        );

    \I__1808\ : InMux
    port map (
            O => \N__20715\,
            I => \sRAM_pointer_read_cry_14\
        );

    \I__1807\ : InMux
    port map (
            O => \N__20712\,
            I => \bfn_2_13_0_\
        );

    \I__1806\ : InMux
    port map (
            O => \N__20709\,
            I => \sRAM_pointer_read_cry_16\
        );

    \I__1805\ : InMux
    port map (
            O => \N__20706\,
            I => \sRAM_pointer_read_cry_17\
        );

    \I__1804\ : CEMux
    port map (
            O => \N__20703\,
            I => \N__20694\
        );

    \I__1803\ : CEMux
    port map (
            O => \N__20702\,
            I => \N__20694\
        );

    \I__1802\ : CEMux
    port map (
            O => \N__20701\,
            I => \N__20694\
        );

    \I__1801\ : GlobalMux
    port map (
            O => \N__20694\,
            I => \N__20691\
        );

    \I__1800\ : gio2CtrlBuf
    port map (
            O => \N__20691\,
            I => \N_28_g\
        );

    \I__1799\ : InMux
    port map (
            O => \N__20688\,
            I => \N__20685\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__20685\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__20682\,
            I => \N__20679\
        );

    \I__1796\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20676\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__20676\,
            I => \spi_master_inst.sclk_gen_u0.sclk_count_i_s_0\
        );

    \I__1794\ : InMux
    port map (
            O => \N__20673\,
            I => \sRAM_pointer_read_cry_1\
        );

    \I__1793\ : InMux
    port map (
            O => \N__20670\,
            I => \sRAM_pointer_read_cry_2\
        );

    \I__1792\ : InMux
    port map (
            O => \N__20667\,
            I => \sRAM_pointer_read_cry_3\
        );

    \I__1791\ : InMux
    port map (
            O => \N__20664\,
            I => \sRAM_pointer_read_cry_4\
        );

    \I__1790\ : InMux
    port map (
            O => \N__20661\,
            I => \sRAM_pointer_read_cry_5\
        );

    \I__1789\ : InMux
    port map (
            O => \N__20658\,
            I => \sRAM_pointer_read_cry_6\
        );

    \I__1788\ : InMux
    port map (
            O => \N__20655\,
            I => \bfn_2_12_0_\
        );

    \I__1787\ : InMux
    port map (
            O => \N__20652\,
            I => \sRAM_pointer_read_cry_8\
        );

    \I__1786\ : InMux
    port map (
            O => \N__20649\,
            I => \sRAM_pointer_read_cry_9\
        );

    \I__1785\ : InMux
    port map (
            O => \N__20646\,
            I => \sRAM_pointer_read_cry_10\
        );

    \I__1784\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20640\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__20640\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__20637\,
            I => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3_cascade_\
        );

    \I__1781\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20631\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__20631\,
            I => \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1\
        );

    \I__1779\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20622\
        );

    \I__1778\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20622\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__20622\,
            I => \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__20619\,
            I => \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i_cascade_\
        );

    \I__1775\ : InMux
    port map (
            O => \N__20616\,
            I => \bfn_2_11_0_\
        );

    \I__1774\ : InMux
    port map (
            O => \N__20613\,
            I => \sRAM_pointer_read_cry_0\
        );

    \I__1773\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20607\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__20607\,
            I => \N__20604\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__20604\,
            I => \N__20601\
        );

    \I__1770\ : Span4Mux_h
    port map (
            O => \N__20601\,
            I => \N__20598\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__20598\,
            I => button_mode_c
        );

    \I__1768\ : IoInMux
    port map (
            O => \N__20595\,
            I => \N__20592\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__20592\,
            I => \N__20589\
        );

    \I__1766\ : Span4Mux_s0_h
    port map (
            O => \N__20589\,
            I => \N__20586\
        );

    \I__1765\ : Span4Mux_v
    port map (
            O => \N__20586\,
            I => \N__20583\
        );

    \I__1764\ : Span4Mux_v
    port map (
            O => \N__20583\,
            I => \N__20580\
        );

    \I__1763\ : Span4Mux_h
    port map (
            O => \N__20580\,
            I => \N__20577\
        );

    \I__1762\ : Odrv4
    port map (
            O => \N__20577\,
            I => \button_mode_ibuf_RNIN5KZ0Z7\
        );

    \I__1761\ : IoInMux
    port map (
            O => \N__20574\,
            I => \N__20571\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__20571\,
            I => \N__20568\
        );

    \I__1759\ : Span12Mux_s7_v
    port map (
            O => \N__20568\,
            I => \N__20565\
        );

    \I__1758\ : Odrv12
    port map (
            O => \N__20565\,
            I => \DAC_cs_c\
        );

    \I__1757\ : IoInMux
    port map (
            O => \N__20562\,
            I => \N__20559\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__20559\,
            I => \N__20556\
        );

    \I__1755\ : Span4Mux_s0_h
    port map (
            O => \N__20556\,
            I => \N__20553\
        );

    \I__1754\ : Span4Mux_h
    port map (
            O => \N__20553\,
            I => \N__20550\
        );

    \I__1753\ : Sp12to4
    port map (
            O => \N__20550\,
            I => \N__20547\
        );

    \I__1752\ : Span12Mux_v
    port map (
            O => \N__20547\,
            I => \N__20544\
        );

    \I__1751\ : Span12Mux_h
    port map (
            O => \N__20544\,
            I => \N__20541\
        );

    \I__1750\ : Odrv12
    port map (
            O => \N__20541\,
            I => \pll128M2_inst.pll_clk128\
        );

    \I__1749\ : IoInMux
    port map (
            O => \N__20538\,
            I => \N__20535\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__20535\,
            I => \N__20532\
        );

    \I__1747\ : Span4Mux_s3_v
    port map (
            O => \N__20532\,
            I => \N__20529\
        );

    \I__1746\ : Sp12to4
    port map (
            O => \N__20529\,
            I => \N__20526\
        );

    \I__1745\ : Span12Mux_h
    port map (
            O => \N__20526\,
            I => \N__20523\
        );

    \I__1744\ : Span12Mux_v
    port map (
            O => \N__20523\,
            I => \N__20520\
        );

    \I__1743\ : Odrv12
    port map (
            O => \N__20520\,
            I => clk_c
        );

    \I__1742\ : IoInMux
    port map (
            O => \N__20517\,
            I => \N__20514\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__20514\,
            I => \N__20511\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__20511\,
            I => \pll128M2_inst.pll_clk64_0\
        );

    \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C\ : INV
    port map (
            O => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            I => \N__30702\
        );

    \INVspi_slave_inst.tx_done_neg_sclk_iC\ : INV
    port map (
            O => \INVspi_slave_inst.tx_done_neg_sclk_iC_net\,
            I => \N__30701\
        );

    \INVspi_slave_inst.rx_done_neg_sclk_iC\ : INV
    port map (
            O => \INVspi_slave_inst.rx_done_neg_sclk_iC_net\,
            I => \N__30699\
        );

    \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C\ : INV
    port map (
            O => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            I => \N__30698\
        );

    \IN_MUX_bfv_22_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_10_0_\
        );

    \IN_MUX_bfv_22_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_scounterdac_cry_8,
            carryinitout => \bfn_22_11_0_\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_sacqtime_cry_7,
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_sacqtime_cry_15,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_sacqtime_cry_23,
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_9_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_3_0_\
        );

    \IN_MUX_bfv_3_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_4_0_\
        );

    \IN_MUX_bfv_3_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO\,
            carryinitout => \bfn_3_5_0_\
        );

    \IN_MUX_bfv_15_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_10_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_6_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un7_spon_cry_7,
            carryinitout => \bfn_6_12_0_\
        );

    \IN_MUX_bfv_6_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un7_spon_cry_15,
            carryinitout => \bfn_6_13_0_\
        );

    \IN_MUX_bfv_6_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un7_spon_cry_23,
            carryinitout => \bfn_6_14_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_sdacdyn_cry_7,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_sdacdyn_cry_15,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_sdacdyn_cry_23,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_spoff_cry_7,
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_spoff_cry_15,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_spoff_cry_23,
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_speriod_cry_7,
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_speriod_cry_15,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_speriod_cry_23,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_sacqtime_cry_7,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_sacqtime_cry_15,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un4_sacqtime_cry_23,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_spoff_cry_7,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_spoff_cry_15,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_spoff_cry_23,
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un10_trig_prev_cry_7,
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_15_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_2_0_\
        );

    \IN_MUX_bfv_10_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_2_0_\
        );

    \IN_MUX_bfv_3_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_3_0_\
        );

    \IN_MUX_bfv_5_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_5_0_\
        );

    \IN_MUX_bfv_10_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_6_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_button_debounce_counter_cry_8,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un1_button_debounce_counter_cry_16,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO\,
            carryinitout => \bfn_8_20_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sRAM_pointer_write_cry_7\,
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sRAM_pointer_write_cry_15\,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sRAM_pointer_read_cry_7\,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sRAM_pointer_read_cry_15\,
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sCounter_cry_7\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sCounter_cry_15\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_15_0_\
        );

    \reset_rpi_ibuf_RNIIUT3_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__27288\,
            GLOBALBUFFEROUTPUT => \LED3_c_i_g\
        );

    \sEEPointerReset_RNI2CQM_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__26601\,
            GLOBALBUFFEROUTPUT => \N_26_g\
        );

    \pll128M2_inst.PLLOUTCOREB_derived_clock_RNI5L14\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__20517\,
            GLOBALBUFFEROUTPUT => pll_clk64_0_g
        );

    \spi_sclk_inferred_clock_RNIH8F3\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__28701\,
            GLOBALBUFFEROUTPUT => spi_sclk_g
        );

    \sEEPointerReset_RNILL2C1_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__27849\,
            GLOBALBUFFEROUTPUT => \N_28_g\
        );

    \pll128M2_inst.PLLOUTCOREA_derived_clock_RNI4765\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__20562\,
            GLOBALBUFFEROUTPUT => pll_clk128_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \sCounterDAC_RNIBR1C_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__53346\,
            GLOBALBUFFEROUTPUT => op_eq_scounterdac10_g
        );

    \button_mode_ibuf_RNIN5K7_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__20595\,
            GLOBALBUFFEROUTPUT => \N_3089_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \button_mode_ibuf_RNIN5K7_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__32691\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20610\,
            lcout => \button_mode_ibuf_RNIN5KZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.o_slave_csn_0_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21300\,
            lcout => \DAC_cs_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53259\,
            ce => 'H',
            sr => \N__53148\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIIUTC1_7_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20812\,
            in1 => \N__21109\,
            in2 => \N__20757\,
            in3 => \N__21085\,
            lcout => \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_1_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111110101010"
        )
    port map (
            in0 => \N__20874\,
            in1 => \N__20628\,
            in2 => \N__22536\,
            in3 => \N__20790\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53265\,
            ce => 'H',
            sr => \N__53147\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_0_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__22532\,
            in1 => \N__20627\,
            in2 => \N__20682\,
            in3 => \N__20789\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53265\,
            ce => 'H',
            sr => \N__53147\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52_2_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__22637\,
            in1 => \N__21299\,
            in2 => \N__21702\,
            in3 => \N__20643\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_RNI06S51_5_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__20927\,
            in1 => \N__21408\,
            in2 => \N__20910\,
            in3 => \N__21168\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3\,
            ltout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIL1LO1_2_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__22638\,
            in1 => \_gnd_net_\,
            in2 => \N__20637\,
            in3 => \N__21700\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIL2KE2_1_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__20839\,
            in1 => \N__20864\,
            in2 => \N__20892\,
            in3 => \N__20634\,
            lcout => \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i\,
            ltout => \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_start_i_RNIPPNJ2_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20619\,
            in3 => \N__22531\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_0_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001111101000000"
        )
    port map (
            in0 => \N__21026\,
            in1 => \N__20736\,
            in2 => \N__20994\,
            in3 => \N__21172\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53272\,
            ce => 'H',
            sr => \N__53144\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_1_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010011110000"
        )
    port map (
            in0 => \N__21027\,
            in1 => \N__20943\,
            in2 => \N__21416\,
            in3 => \N__20984\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53272\,
            ce => 'H',
            sr => \N__53144\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_6_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25752\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53272\,
            ce => 'H',
            sr => \N__53144\
        );

    \sRAM_pointer_read_0_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33548\,
            in1 => \N__29750\,
            in2 => \_gnd_net_\,
            in3 => \N__20616\,
            lcout => \sRAM_pointer_readZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \sRAM_pointer_read_cry_0\,
            clk => \N__47843\,
            ce => \N__20701\,
            sr => \N__53118\
        );

    \sRAM_pointer_read_1_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33544\,
            in1 => \N__29675\,
            in2 => \_gnd_net_\,
            in3 => \N__20613\,
            lcout => \sRAM_pointer_readZ0Z_1\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_0\,
            carryout => \sRAM_pointer_read_cry_1\,
            clk => \N__47843\,
            ce => \N__20701\,
            sr => \N__53118\
        );

    \sRAM_pointer_read_2_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33549\,
            in1 => \N__28067\,
            in2 => \_gnd_net_\,
            in3 => \N__20673\,
            lcout => \sRAM_pointer_readZ0Z_2\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_1\,
            carryout => \sRAM_pointer_read_cry_2\,
            clk => \N__47843\,
            ce => \N__20701\,
            sr => \N__53118\
        );

    \sRAM_pointer_read_3_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33545\,
            in1 => \N__28673\,
            in2 => \_gnd_net_\,
            in3 => \N__20670\,
            lcout => \sRAM_pointer_readZ0Z_3\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_2\,
            carryout => \sRAM_pointer_read_cry_3\,
            clk => \N__47843\,
            ce => \N__20701\,
            sr => \N__53118\
        );

    \sRAM_pointer_read_4_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33550\,
            in1 => \N__28637\,
            in2 => \_gnd_net_\,
            in3 => \N__20667\,
            lcout => \sRAM_pointer_readZ0Z_4\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_3\,
            carryout => \sRAM_pointer_read_cry_4\,
            clk => \N__47843\,
            ce => \N__20701\,
            sr => \N__53118\
        );

    \sRAM_pointer_read_5_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33546\,
            in1 => \N__28592\,
            in2 => \_gnd_net_\,
            in3 => \N__20664\,
            lcout => \sRAM_pointer_readZ0Z_5\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_4\,
            carryout => \sRAM_pointer_read_cry_5\,
            clk => \N__47843\,
            ce => \N__20701\,
            sr => \N__53118\
        );

    \sRAM_pointer_read_6_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33551\,
            in1 => \N__28547\,
            in2 => \_gnd_net_\,
            in3 => \N__20661\,
            lcout => \sRAM_pointer_readZ0Z_6\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_5\,
            carryout => \sRAM_pointer_read_cry_6\,
            clk => \N__47843\,
            ce => \N__20701\,
            sr => \N__53118\
        );

    \sRAM_pointer_read_7_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33547\,
            in1 => \N__28499\,
            in2 => \_gnd_net_\,
            in3 => \N__20658\,
            lcout => \sRAM_pointer_readZ0Z_7\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_6\,
            carryout => \sRAM_pointer_read_cry_7\,
            clk => \N__47843\,
            ce => \N__20701\,
            sr => \N__53118\
        );

    \sRAM_pointer_read_8_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33459\,
            in1 => \N__28451\,
            in2 => \_gnd_net_\,
            in3 => \N__20655\,
            lcout => \sRAM_pointer_readZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \sRAM_pointer_read_cry_8\,
            clk => \N__47852\,
            ce => \N__20702\,
            sr => \N__53105\
        );

    \sRAM_pointer_read_9_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33446\,
            in1 => \N__28403\,
            in2 => \_gnd_net_\,
            in3 => \N__20652\,
            lcout => \sRAM_pointer_readZ0Z_9\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_8\,
            carryout => \sRAM_pointer_read_cry_9\,
            clk => \N__47852\,
            ce => \N__20702\,
            sr => \N__53105\
        );

    \sRAM_pointer_read_10_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33456\,
            in1 => \N__29630\,
            in2 => \_gnd_net_\,
            in3 => \N__20649\,
            lcout => \sRAM_pointer_readZ0Z_10\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_9\,
            carryout => \sRAM_pointer_read_cry_10\,
            clk => \N__47852\,
            ce => \N__20702\,
            sr => \N__53105\
        );

    \sRAM_pointer_read_11_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33443\,
            in1 => \N__30392\,
            in2 => \_gnd_net_\,
            in3 => \N__20646\,
            lcout => \sRAM_pointer_readZ0Z_11\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_10\,
            carryout => \sRAM_pointer_read_cry_11\,
            clk => \N__47852\,
            ce => \N__20702\,
            sr => \N__53105\
        );

    \sRAM_pointer_read_12_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33457\,
            in1 => \N__30338\,
            in2 => \_gnd_net_\,
            in3 => \N__20724\,
            lcout => \sRAM_pointer_readZ0Z_12\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_11\,
            carryout => \sRAM_pointer_read_cry_12\,
            clk => \N__47852\,
            ce => \N__20702\,
            sr => \N__53105\
        );

    \sRAM_pointer_read_13_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33444\,
            in1 => \N__30302\,
            in2 => \_gnd_net_\,
            in3 => \N__20721\,
            lcout => \sRAM_pointer_readZ0Z_13\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_12\,
            carryout => \sRAM_pointer_read_cry_13\,
            clk => \N__47852\,
            ce => \N__20702\,
            sr => \N__53105\
        );

    \sRAM_pointer_read_14_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33458\,
            in1 => \N__28289\,
            in2 => \_gnd_net_\,
            in3 => \N__20718\,
            lcout => \sRAM_pointer_readZ0Z_14\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_13\,
            carryout => \sRAM_pointer_read_cry_14\,
            clk => \N__47852\,
            ce => \N__20702\,
            sr => \N__53105\
        );

    \sRAM_pointer_read_15_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33445\,
            in1 => \N__28241\,
            in2 => \_gnd_net_\,
            in3 => \N__20715\,
            lcout => \sRAM_pointer_readZ0Z_15\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_14\,
            carryout => \sRAM_pointer_read_cry_15\,
            clk => \N__47852\,
            ce => \N__20702\,
            sr => \N__53105\
        );

    \sRAM_pointer_read_16_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33503\,
            in1 => \N__28199\,
            in2 => \_gnd_net_\,
            in3 => \N__20712\,
            lcout => \sRAM_pointer_readZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \sRAM_pointer_read_cry_16\,
            clk => \N__47853\,
            ce => \N__20703\,
            sr => \N__53089\
        );

    \sRAM_pointer_read_17_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33484\,
            in1 => \N__28151\,
            in2 => \_gnd_net_\,
            in3 => \N__20709\,
            lcout => \sRAM_pointer_readZ0Z_17\,
            ltout => OPEN,
            carryin => \sRAM_pointer_read_cry_16\,
            carryout => \sRAM_pointer_read_cry_17\,
            clk => \N__47853\,
            ce => \N__20703\,
            sr => \N__53089\
        );

    \sRAM_pointer_read_18_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33504\,
            in1 => \N__28109\,
            in2 => \_gnd_net_\,
            in3 => \N__20706\,
            lcout => \sRAM_pointer_readZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47853\,
            ce => \N__20703\,
            sr => \N__53089\
        );

    \spi_master_inst.sclk_gen_u0.div_clk_i_RNO_0_LC_3_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20863\,
            in1 => \N__20755\,
            in2 => \N__20844\,
            in3 => \N__20813\,
            lcout => \spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_0_LC_3_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20688\,
            in2 => \_gnd_net_\,
            in3 => \N__20895\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_i_s_0\,
            ltout => OPEN,
            carryin => \bfn_3_3_0_\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_1_LC_3_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20888\,
            in2 => \_gnd_net_\,
            in3 => \N__20868\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_i_s_1\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_2_LC_3_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20791\,
            in1 => \N__20865\,
            in2 => \_gnd_net_\,
            in3 => \N__20847\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2\,
            clk => \N__53260\,
            ce => 'H',
            sr => \N__53146\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_3_LC_3_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20786\,
            in1 => \N__20840\,
            in2 => \_gnd_net_\,
            in3 => \N__20823\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3\,
            clk => \N__53260\,
            ce => 'H',
            sr => \N__53146\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_4_LC_3_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20792\,
            in1 => \N__21086\,
            in2 => \_gnd_net_\,
            in3 => \N__20820\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4\,
            clk => \N__53260\,
            ce => 'H',
            sr => \N__53146\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_5_LC_3_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20787\,
            in1 => \N__21110\,
            in2 => \_gnd_net_\,
            in3 => \N__20817\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5\,
            clk => \N__53260\,
            ce => 'H',
            sr => \N__53146\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_6_LC_3_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20793\,
            in1 => \N__20814\,
            in2 => \_gnd_net_\,
            in3 => \N__20796\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5\,
            carryout => \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6\,
            clk => \N__53260\,
            ce => 'H',
            sr => \N__53146\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_i_7_LC_3_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20788\,
            in1 => \N__20756\,
            in2 => \_gnd_net_\,
            in3 => \N__20760\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53260\,
            ce => 'H',
            sr => \N__53146\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_c_LC_3_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20735\,
            in2 => \N__21176\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_4_0_\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_LUT4_0_LC_3_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21409\,
            in2 => \_gnd_net_\,
            in3 => \N__20937\,
            lcout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_LUT4_0_LC_3_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21701\,
            in2 => \_gnd_net_\,
            in3 => \N__20934\,
            lcout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_LUT4_0_LC_3_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22639\,
            in2 => \_gnd_net_\,
            in3 => \N__20931\,
            lcout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_4_LC_3_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20986\,
            in1 => \N__20928\,
            in2 => \_gnd_net_\,
            in3 => \N__20916\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4\,
            clk => \N__53266\,
            ce => 'H',
            sr => \N__53145\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_0_LC_3_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37824\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_1_LC_3_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__37907\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_2_LC_3_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37828\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO\,
            carryout => \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_5_LC_3_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20909\,
            in2 => \_gnd_net_\,
            in3 => \N__20913\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53270\,
            ce => \N__20985\,
            sr => \N__53143\
        );

    \spi_master_inst.sclk_gen_u0.o_sclk_RNIH6AC_LC_3_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__22492\,
            in1 => \N__23688\,
            in2 => \_gnd_net_\,
            in3 => \N__21059\,
            lcout => \spi_master_inst.o_sclk_RNIH6AC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_ft_ibuf_RNI4OFN_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__23892\,
            in1 => \N__23964\,
            in2 => \_gnd_net_\,
            in3 => \N__24040\,
            lcout => un3_trig_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_ft_ibuf_RNI4OFN_0_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__23931\,
            in1 => \N__23907\,
            in2 => \_gnd_net_\,
            in3 => \N__24024\,
            lcout => un3_trig_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI70MD9_0_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__21297\,
            in1 => \N__21429\,
            in2 => \N__21387\,
            in3 => \N__21180\,
            lcout => \DAC_mosi_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.div_clk_i_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__21129\,
            in1 => \N__21117\,
            in2 => \_gnd_net_\,
            in3 => \N__21093\,
            lcout => \spi_master_inst.sclk_gen_u0.div_clk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53255\,
            ce => 'H',
            sr => \N__53142\
        );

    \spi_master_inst.sclk_gen_u0.o_sclk_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22483\,
            in2 => \_gnd_net_\,
            in3 => \N__23694\,
            lcout => \DAC_sclk_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53255\,
            ce => 'H',
            sr => \N__53142\
        );

    \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_i_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011011000"
        )
    port map (
            in0 => \N__20995\,
            in1 => \N__21028\,
            in2 => \N__27026\,
            in3 => \N__21296\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53255\,
            ce => 'H',
            sr => \N__53142\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_2_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001110001001100"
        )
    port map (
            in0 => \N__21030\,
            in1 => \N__21692\,
            in2 => \N__21000\,
            in3 => \N__21039\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53255\,
            ce => 'H',
            sr => \N__53142\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_3_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011010001110000"
        )
    port map (
            in0 => \N__21029\,
            in1 => \N__20999\,
            in2 => \N__22636\,
            in3 => \N__20952\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53255\,
            ce => 'H',
            sr => \N__53142\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_0_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101111101110"
        )
    port map (
            in0 => \N__21460\,
            in1 => \N__21570\,
            in2 => \_gnd_net_\,
            in3 => \N__21255\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_5_0_\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_0\,
            clk => \N__53261\,
            ce => 'H',
            sr => \N__53141\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_1_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21455\,
            in1 => \N__21624\,
            in2 => \_gnd_net_\,
            in3 => \N__21252\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_0\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_1\,
            clk => \N__53261\,
            ce => 'H',
            sr => \N__53141\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_2_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21461\,
            in1 => \N__21605\,
            in2 => \_gnd_net_\,
            in3 => \N__21249\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_1\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_2\,
            clk => \N__53261\,
            ce => 'H',
            sr => \N__53141\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_3_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21456\,
            in1 => \N__21642\,
            in2 => \_gnd_net_\,
            in3 => \N__21246\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_2\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_3\,
            clk => \N__53261\,
            ce => 'H',
            sr => \N__53141\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_4_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21462\,
            in1 => \N__21192\,
            in2 => \_gnd_net_\,
            in3 => \N__21243\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_3\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_4\,
            clk => \N__53261\,
            ce => 'H',
            sr => \N__53141\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_5_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21457\,
            in1 => \N__21219\,
            in2 => \_gnd_net_\,
            in3 => \N__21240\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_4\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_5\,
            clk => \N__53261\,
            ce => 'H',
            sr => \N__53141\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_6_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21458\,
            in1 => \N__21231\,
            in2 => \_gnd_net_\,
            in3 => \N__21237\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_5\,
            carryout => \spi_master_inst.sclk_gen_u0.delay_count_i_cry_6\,
            clk => \N__53261\,
            ce => 'H',
            sr => \N__53141\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_7_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21206\,
            in1 => \N__21459\,
            in2 => \_gnd_net_\,
            in3 => \N__21234\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53261\,
            ce => 'H',
            sr => \N__53141\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_RNIQU1N1_7_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21230\,
            in1 => \N__21218\,
            in2 => \N__21207\,
            in3 => \N__21191\,
            lcout => \spi_master_inst.sclk_gen_u0.N_1666\,
            ltout => \spi_master_inst.sclk_gen_u0.N_1666_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_0_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__21321\,
            in1 => \N__21315\,
            in2 => \N__21324\,
            in3 => \N__21471\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53267\,
            ce => 'H',
            sr => \N__53136\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_RNIAE1N1_0_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__21569\,
            in1 => \N__21623\,
            in2 => \N__21606\,
            in3 => \N__21641\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4\,
            ltout => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0IPL3_0_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21314\,
            in2 => \N__21306\,
            in3 => \N__21585\,
            lcout => \spi_master_inst.sclk_gen_u0.N_48\,
            ltout => \spi_master_inst.sclk_gen_u0.N_48_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_4_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__23727\,
            in1 => \_gnd_net_\,
            in2 => \N__21303\,
            in3 => \N__27003\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53267\,
            ce => 'H',
            sr => \N__53136\
        );

    \spi_master_inst.sclk_gen_u0.o_ss_start_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101110100"
        )
    port map (
            in0 => \N__27002\,
            in1 => \N__23726\,
            in2 => \N__21298\,
            in3 => \N__21470\,
            lcout => \spi_master_inst.ss_start_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53267\,
            ce => 'H',
            sr => \N__53136\
        );

    \trig_ft_ibuf_RNI4OFN_2_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__23901\,
            in1 => \N__23965\,
            in2 => \_gnd_net_\,
            in3 => \N__24041\,
            lcout => un3_trig_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_ft_ibuf_RNI4OFN_3_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__23966\,
            in1 => \_gnd_net_\,
            in2 => \N__24056\,
            in3 => \N__23902\,
            lcout => un3_trig_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sSingleCont_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22215\,
            in2 => \_gnd_net_\,
            in3 => \N__21978\,
            lcout => \LED_MODE_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53273\,
            ce => 'H',
            sr => \N__53119\
        );

    \sSPI_MSB0LSB1_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101001001011010"
        )
    port map (
            in0 => \N__27911\,
            in1 => \N__32215\,
            in2 => \N__27956\,
            in3 => \N__31977\,
            lcout => \sSPI_MSB0LSBZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47842\,
            ce => 'H',
            sr => \N__53106\
        );

    \un4_spoff_cry_0_c_inv_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21378\,
            in2 => \N__34245\,
            in3 => \N__21717\,
            lcout => \sEEPonPoff_i_0\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => un4_spoff_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_1_c_inv_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21372\,
            in2 => \N__35064\,
            in3 => \N__21783\,
            lcout => \sEEPonPoff_i_1\,
            ltout => OPEN,
            carryin => un4_spoff_cry_0,
            carryout => un4_spoff_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_2_c_inv_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21777\,
            in1 => \N__21366\,
            in2 => \N__34968\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoff_i_2\,
            ltout => OPEN,
            carryin => un4_spoff_cry_1,
            carryout => un4_spoff_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_3_c_inv_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34857\,
            in2 => \N__21360\,
            in3 => \N__21771\,
            lcout => \sEEPonPoff_i_3\,
            ltout => OPEN,
            carryin => un4_spoff_cry_2,
            carryout => un4_spoff_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_4_c_inv_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21351\,
            in2 => \N__36883\,
            in3 => \N__21765\,
            lcout => \sEEPonPoff_i_4\,
            ltout => OPEN,
            carryin => un4_spoff_cry_3,
            carryout => un4_spoff_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_5_c_inv_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34728\,
            in2 => \N__21345\,
            in3 => \N__21759\,
            lcout => \sEEPonPoff_i_5\,
            ltout => OPEN,
            carryin => un4_spoff_cry_4,
            carryout => un4_spoff_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_6_c_inv_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21753\,
            in1 => \N__21336\,
            in2 => \N__34620\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoff_i_6\,
            ltout => OPEN,
            carryin => un4_spoff_cry_5,
            carryout => un4_spoff_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_7_c_inv_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21330\,
            in2 => \N__34494\,
            in3 => \N__21747\,
            lcout => \sEEPonPoff_i_7\,
            ltout => OPEN,
            carryin => un4_spoff_cry_6,
            carryout => un4_spoff_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_8_c_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37841\,
            in2 => \N__35889\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => un4_spoff_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_9_c_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35763\,
            in2 => \N__37911\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_8,
            carryout => un4_spoff_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_10_c_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37829\,
            in2 => \N__35654\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_9,
            carryout => un4_spoff_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_11_c_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35541\,
            in2 => \N__37908\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_10,
            carryout => un4_spoff_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_12_c_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37833\,
            in2 => \N__35418\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_11,
            carryout => un4_spoff_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_13_c_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35311\,
            in2 => \N__37909\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_12,
            carryout => un4_spoff_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_14_c_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37837\,
            in2 => \N__35208\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_13,
            carryout => un4_spoff_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_15_c_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36659\,
            in2 => \N__37910\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_14,
            carryout => un4_spoff_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_16_c_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37865\,
            in2 => \N__36546\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => un4_spoff_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_17_c_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36444\,
            in2 => \N__37929\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_16,
            carryout => un4_spoff_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_18_c_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37869\,
            in2 => \N__36346\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_17,
            carryout => un4_spoff_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_19_c_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36254\,
            in2 => \N__37930\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_18,
            carryout => un4_spoff_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_20_c_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37873\,
            in2 => \N__36169\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_19,
            carryout => un4_spoff_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIR3KA_20_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36072\,
            in2 => \N__37928\,
            in3 => \N__36158\,
            lcout => un1_reset_rpi_inv_2_i_o3_8,
            ltout => OPEN,
            carryin => un4_spoff_cry_20,
            carryout => un4_spoff_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_22_c_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37874\,
            in2 => \N__36000\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_21,
            carryout => un4_spoff_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_23_c_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37088\,
            in2 => \N__37931\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_spoff_cry_22,
            carryout => un4_spoff_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_spoff_cry_23_THRU_LUT4_0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21432\,
            lcout => \un4_spoff_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIUNHB4_1_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21486\,
            in1 => \N__21477\,
            in2 => \_gnd_net_\,
            in3 => \N__21423\,
            lcout => \spi_master_inst.spi_data_path_u1.N_1423\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI60IB4_1_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21651\,
            in1 => \N__21507\,
            in2 => \_gnd_net_\,
            in3 => \N__21422\,
            lcout => \spi_master_inst.spi_data_path_u1.N_1416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI73G42_2_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21694\,
            in1 => \N__21990\,
            in2 => \_gnd_net_\,
            in3 => \N__21984\,
            lcout => \spi_master_inst.spi_data_path_u1.N_1415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4Q_14_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22458\,
            in1 => \N__21501\,
            in2 => \_gnd_net_\,
            in3 => \N__22628\,
            lcout => OPEN,
            ltout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIICLT1_2_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__21695\,
            in1 => \_gnd_net_\,
            in2 => \N__21489\,
            in3 => \N__22398\,
            lcout => \spi_master_inst.spi_data_path_u1.N_1419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01_0_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22627\,
            in1 => \N__22437\,
            in2 => \_gnd_net_\,
            in3 => \N__22446\,
            lcout => OPEN,
            ltout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI3VF42_2_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22569\,
            in1 => \_gnd_net_\,
            in2 => \N__21480\,
            in3 => \N__21693\,
            lcout => \spi_master_inst.spi_data_path_u1.N_1422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI1JPL3_1_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21524\,
            in2 => \_gnd_net_\,
            in3 => \N__21948\,
            lcout => \spi_master_inst.sclk_gen_u0.N_1520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4Q_11_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23772\,
            in1 => \N__23580\,
            in2 => \_gnd_net_\,
            in3 => \N__22617\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNI6TQC_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21536\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_start_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4Q_15_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22618\,
            in1 => \N__22422\,
            in2 => \_gnd_net_\,
            in3 => \N__23781\,
            lcout => OPEN,
            ltout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIMGLT1_2_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__21711\,
            in1 => \_gnd_net_\,
            in2 => \N__21705\,
            in3 => \N__21696\,
            lcout => \spi_master_inst.spi_data_path_u1.N_1412\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_RNI6OGR_1_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21640\,
            in2 => \_gnd_net_\,
            in3 => \N__21622\,
            lcout => OPEN,
            ltout => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4D3E3_0_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__21601\,
            in1 => \N__21584\,
            in2 => \N__21573\,
            in3 => \N__21568\,
            lcout => \spi_master_inst.sclk_gen_u0.N_1515\,
            ltout => \spi_master_inst.sclk_gen_u0.N_1515_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0RFT3_1_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21964\,
            in2 => \N__21552\,
            in3 => \N__21520\,
            lcout => \spi_master_inst.sclk_gen_u0.N_36\,
            ltout => \spi_master_inst.sclk_gen_u0.N_36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNO_0_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__23717\,
            in1 => \N__27000\,
            in2 => \N__21549\,
            in3 => \N__21546\,
            lcout => OPEN,
            ltout => \spi_master_inst.sclk_gen_u0.N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.delay_count_start_i_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111110001101"
        )
    port map (
            in0 => \N__23692\,
            in1 => \N__21537\,
            in2 => \N__21540\,
            in3 => \N__23756\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_count_start_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53256\,
            ce => 'H',
            sr => \N__53120\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_1_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23757\,
            in1 => \N__23693\,
            in2 => \N__21525\,
            in3 => \N__21950\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53256\,
            ce => 'H',
            sr => \N__53120\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_3_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__21965\,
            in1 => \N__27001\,
            in2 => \N__23728\,
            in3 => \N__21951\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53256\,
            ce => 'H',
            sr => \N__53120\
        );

    \sTrigCounter_RNO_2_0_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100011111100"
        )
    port map (
            in0 => \N__24927\,
            in1 => \N__24488\,
            in2 => \N__22091\,
            in3 => \N__29094\,
            lcout => g1_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_ft_ibuf_RNI4OFN_5_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__24057\,
            in1 => \N__23900\,
            in2 => \_gnd_net_\,
            in3 => \N__23970\,
            lcout => un3_trig_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPon_0_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51258\,
            lcout => \sEEPonZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47836\,
            ce => \N__30896\,
            sr => \N__53091\
        );

    \sEEPon_1_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50675\,
            lcout => \sEEPonZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47836\,
            ce => \N__30896\,
            sr => \N__53091\
        );

    \sEEPon_7_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48798\,
            lcout => \sEEPonZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47836\,
            ce => \N__30896\,
            sr => \N__53091\
        );

    \sEEPon_3_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49821\,
            lcout => \sEEPonZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47836\,
            ce => \N__30896\,
            sr => \N__53091\
        );

    \sEEPon_4_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49345\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47836\,
            ce => \N__30896\,
            sr => \N__53091\
        );

    \sEEPon_6_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48306\,
            lcout => \sEEPonZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47836\,
            ce => \N__30896\,
            sr => \N__53091\
        );

    \sEEPon_5_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47118\,
            lcout => \sEEPonZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47827\,
            ce => \N__30900\,
            sr => \N__53080\
        );

    \sEEPon_2_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50283\,
            lcout => \sEEPonZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47827\,
            ce => \N__30900\,
            sr => \N__53080\
        );

    \sEEPonPoff_0_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51232\,
            lcout => \sEEPonPoffZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47819\,
            ce => \N__30810\,
            sr => \N__53068\
        );

    \sEEPonPoff_1_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50676\,
            lcout => \sEEPonPoffZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47819\,
            ce => \N__30810\,
            sr => \N__53068\
        );

    \sEEPonPoff_2_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50285\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoffZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47819\,
            ce => \N__30810\,
            sr => \N__53068\
        );

    \sEEPonPoff_3_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49823\,
            lcout => \sEEPonPoffZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47819\,
            ce => \N__30810\,
            sr => \N__53068\
        );

    \sEEPonPoff_4_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49347\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoffZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47819\,
            ce => \N__30810\,
            sr => \N__53068\
        );

    \sEEPonPoff_5_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47072\,
            lcout => \sEEPonPoffZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47819\,
            ce => \N__30810\,
            sr => \N__53068\
        );

    \sEEPonPoff_6_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48336\,
            lcout => \sEEPonPoffZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47819\,
            ce => \N__30810\,
            sr => \N__53068\
        );

    \sEEPonPoff_7_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48593\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPonPoffZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47819\,
            ce => \N__30810\,
            sr => \N__53068\
        );

    \un7_spon_cry_0_c_inv_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21741\,
            in1 => \N__21732\,
            in2 => \N__34243\,
            in3 => \_gnd_net_\,
            lcout => \sEEPon_i_0\,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => un7_spon_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_1_c_inv_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21885\,
            in2 => \N__35063\,
            in3 => \N__21726\,
            lcout => \sEEPon_i_1\,
            ltout => OPEN,
            carryin => un7_spon_cry_0,
            carryout => un7_spon_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_2_c_inv_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21879\,
            in1 => \N__21870\,
            in2 => \N__34964\,
            in3 => \_gnd_net_\,
            lcout => \sEEPon_i_2\,
            ltout => OPEN,
            carryin => un7_spon_cry_1,
            carryout => un7_spon_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_3_c_inv_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34851\,
            in2 => \N__21855\,
            in3 => \N__21864\,
            lcout => \sEEPon_i_3\,
            ltout => OPEN,
            carryin => un7_spon_cry_2,
            carryout => un7_spon_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_4_c_inv_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21837\,
            in2 => \N__36882\,
            in3 => \N__21846\,
            lcout => \sEEPon_i_4\,
            ltout => OPEN,
            carryin => un7_spon_cry_3,
            carryout => un7_spon_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_5_c_inv_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21822\,
            in2 => \N__34727\,
            in3 => \N__21831\,
            lcout => \sEEPon_i_5\,
            ltout => OPEN,
            carryin => un7_spon_cry_4,
            carryout => un7_spon_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_6_c_inv_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21804\,
            in2 => \N__34619\,
            in3 => \N__21816\,
            lcout => \sEEPon_i_6\,
            ltout => OPEN,
            carryin => un7_spon_cry_5,
            carryout => un7_spon_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_7_c_inv_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21798\,
            in1 => \N__21789\,
            in2 => \N__34489\,
            in3 => \_gnd_net_\,
            lcout => \sEEPon_i_7\,
            ltout => OPEN,
            carryin => un7_spon_cry_6,
            carryout => un7_spon_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_8_c_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37944\,
            in2 => \N__35881\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_12_0_\,
            carryout => un7_spon_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_9_c_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35767\,
            in2 => \N__37971\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_8,
            carryout => un7_spon_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_10_c_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37932\,
            in2 => \N__35655\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_9,
            carryout => un7_spon_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_11_c_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35536\,
            in2 => \N__37968\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_10,
            carryout => un7_spon_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_12_c_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37936\,
            in2 => \N__35414\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_11,
            carryout => un7_spon_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_13_c_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35315\,
            in2 => \N__37969\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_12,
            carryout => un7_spon_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_14_c_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37940\,
            in2 => \N__35204\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_13,
            carryout => un7_spon_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_15_c_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36655\,
            in2 => \N__37970\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_14,
            carryout => un7_spon_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_16_c_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37912\,
            in2 => \N__36545\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_13_0_\,
            carryout => un7_spon_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_17_c_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36441\,
            in2 => \N__37964\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_16,
            carryout => un7_spon_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_18_c_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37916\,
            in2 => \N__36348\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_17,
            carryout => un7_spon_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_19_c_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36251\,
            in2 => \N__37965\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_18,
            carryout => un7_spon_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_20_c_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37920\,
            in2 => \N__36171\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_19,
            carryout => un7_spon_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_21_c_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36079\,
            in2 => \N__37966\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_20,
            carryout => un7_spon_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_22_c_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37924\,
            in2 => \N__35996\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_21,
            carryout => un7_spon_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un7_spon_cry_23_c_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37079\,
            in2 => \N__37967\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un7_spon_cry_22,
            carryout => un7_spon_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pon_obuf_RNO_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__36956\,
            in1 => \N__36840\,
            in2 => \_gnd_net_\,
            in3 => \N__21921\,
            lcout => \pon_obuf_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_0_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010011100"
        )
    port map (
            in0 => \N__22167\,
            in1 => \N__31350\,
            in2 => \N__32590\,
            in3 => \N__21891\,
            lcout => \sTrigCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47844\,
            ce => 'H',
            sr => \N__27541\
        );

    \sTrigCounter_RNO_0_0_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__24384\,
            in1 => \N__21900\,
            in2 => \N__24310\,
            in3 => \N__24720\,
            lcout => g1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sSPI_MSB0LSB1_RNIFIB13_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__32175\,
            in1 => \N__27981\,
            in2 => \N__27912\,
            in3 => \N__22347\,
            lcout => \un1_spi_data_miso_0_sqmuxa_1_i_0_N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4Q_13_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22630\,
            in1 => \N__23565\,
            in2 => \_gnd_net_\,
            in3 => \N__22404\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01_1_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22410\,
            in1 => \N__22428\,
            in2 => \_gnd_net_\,
            in3 => \N__22629\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEESingleCont_er_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51203\,
            lcout => \sEESingleContZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47849\,
            ce => \N__21930\,
            sr => \N__53121\
        );

    \sTrigCounter_RNO_5_5_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110001010100"
        )
    port map (
            in0 => \N__29106\,
            in1 => \N__24507\,
            in2 => \N__23628\,
            in3 => \N__24942\,
            lcout => g0_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI3LPL3_3_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21966\,
            in2 => \_gnd_net_\,
            in3 => \N__21949\,
            lcout => \spi_master_inst.sclk_gen_u0.N_150_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEESingleCont_er_RNO_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__43287\,
            in1 => \N__31107\,
            in2 => \N__44469\,
            in3 => \N__44751\,
            lcout => \sEESingleCont_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_4_2_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111000100"
        )
    port map (
            in0 => \N__29101\,
            in1 => \N__24429\,
            in2 => \N__24938\,
            in3 => \N__24467\,
            lcout => g0_2_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_prev_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__23972\,
            in1 => \N__23899\,
            in2 => \_gnd_net_\,
            in3 => \N__24059\,
            lcout => \trig_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47837\,
            ce => 'H',
            sr => \N__53092\
        );

    \trig_ft_ibuf_RNIM2UO_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__24058\,
            in1 => \N__23971\,
            in2 => \N__23906\,
            in3 => \N__24464\,
            lcout => \N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_3_3_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111010"
        )
    port map (
            in0 => \N__24465\,
            in1 => \N__24910\,
            in2 => \N__22023\,
            in3 => \N__29099\,
            lcout => g1_0_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_4_3_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111000100"
        )
    port map (
            in0 => \N__29102\,
            in1 => \N__22022\,
            in2 => \N__24939\,
            in3 => \N__24468\,
            lcout => g0_2_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_3_4_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111010"
        )
    port map (
            in0 => \N__24466\,
            in1 => \N__24911\,
            in2 => \N__22008\,
            in3 => \N__29100\,
            lcout => g1_0_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_5_4_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111000100"
        )
    port map (
            in0 => \N__29103\,
            in1 => \N__22007\,
            in2 => \N__24940\,
            in3 => \N__24469\,
            lcout => g0_2_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_4_5_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24229\,
            in1 => \N__24203\,
            in2 => \N__32623\,
            in3 => \N__24602\,
            lcout => OPEN,
            ltout => \g1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_1_5_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31299\,
            in2 => \N__21993\,
            in3 => \N__31387\,
            lcout => g1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPointerReset_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__51257\,
            in1 => \N__43855\,
            in2 => \N__33391\,
            in3 => \N__28959\,
            lcout => \sEEPointerResetZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47828\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sPeriod_prev_RNIRSLG_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24257\,
            in2 => \_gnd_net_\,
            in3 => \N__24361\,
            lcout => un1_reset_rpi_inv_2_i_o3_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPeriod_0_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51259\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47820\,
            ce => \N__24519\,
            sr => \N__53069\
        );

    \sEEPeriod_1_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50592\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47820\,
            ce => \N__24519\,
            sr => \N__53069\
        );

    \sEEPeriod_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50282\,
            lcout => \sEEPeriodZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47820\,
            ce => \N__24519\,
            sr => \N__53069\
        );

    \sEEPeriod_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49820\,
            lcout => \sEEPeriodZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47820\,
            ce => \N__24519\,
            sr => \N__53069\
        );

    \sEEPeriod_4_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49354\,
            lcout => \sEEPeriodZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47820\,
            ce => \N__24519\,
            sr => \N__53069\
        );

    \sEEPeriod_5_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47063\,
            lcout => \sEEPeriodZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47820\,
            ce => \N__24519\,
            sr => \N__53069\
        );

    \sEEPeriod_6_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48153\,
            lcout => \sEEPeriodZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47820\,
            ce => \N__24519\,
            sr => \N__53069\
        );

    \sEEPeriod_7_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48776\,
            lcout => \sEEPeriodZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47820\,
            ce => \N__24519\,
            sr => \N__53069\
        );

    \sTrigCounter_RNO_3_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111010"
        )
    port map (
            in0 => \N__24490\,
            in1 => \N__24878\,
            in2 => \N__22133\,
            in3 => \N__29097\,
            lcout => g1_0_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigInternal_prev_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29098\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEETrigInternal_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47812\,
            ce => 'H',
            sr => \N__53058\
        );

    \sEETrigInternal_prev_RNISEUG_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24874\,
            in2 => \_gnd_net_\,
            in3 => \N__29095\,
            lcout => OPEN,
            ltout => \sEETrigInternal_prev_RNISEUGZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigInternal_RNIOMLD1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__22040\,
            in1 => \N__22280\,
            in2 => \N__22026\,
            in3 => \N__24491\,
            lcout => \sTrigInternal_RNIOMLDZ0Z1\,
            ltout => \sTrigInternal_RNIOMLDZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigInternal_RNO_0_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__36958\,
            in1 => \N__36859\,
            in2 => \N__22053\,
            in3 => \N__24816\,
            lcout => OPEN,
            ltout => \sTrigInternal_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigInternal_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100000011"
        )
    port map (
            in0 => \N__24740\,
            in1 => \N__22050\,
            in2 => \N__22044\,
            in3 => \N__24718\,
            lcout => \sTrigInternalZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47812\,
            ce => 'H',
            sr => \N__53058\
        );

    \trig_prev_RNIIHS91_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111000100"
        )
    port map (
            in0 => \N__29096\,
            in1 => \N__22041\,
            in2 => \N__24909\,
            in3 => \N__24489\,
            lcout => \N_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPeriod_16_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51260\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47803\,
            ce => \N__28923\,
            sr => \N__53048\
        );

    \sEEPeriod_17_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50599\,
            lcout => \sEEPeriodZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47803\,
            ce => \N__28923\,
            sr => \N__53048\
        );

    \sEEPeriod_18_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50284\,
            lcout => \sEEPeriodZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47803\,
            ce => \N__28923\,
            sr => \N__53048\
        );

    \sEEPeriod_19_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49822\,
            lcout => \sEEPeriodZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47803\,
            ce => \N__28923\,
            sr => \N__53048\
        );

    \sEEPeriod_20_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49346\,
            lcout => \sEEPeriodZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47803\,
            ce => \N__28923\,
            sr => \N__53048\
        );

    \sEEPeriod_21_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47064\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47803\,
            ce => \N__28923\,
            sr => \N__53048\
        );

    \sEEPeriod_22_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48305\,
            lcout => \sEEPeriodZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47803\,
            ce => \N__28923\,
            sr => \N__53048\
        );

    \sEEPeriod_23_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48769\,
            lcout => \sEEPeriodZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47803\,
            ce => \N__28923\,
            sr => \N__53048\
        );

    \sTrigCounter_RNO_4_1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111000100"
        )
    port map (
            in0 => \N__29105\,
            in1 => \N__22134\,
            in2 => \N__24945\,
            in3 => \N__24509\,
            lcout => g0_2_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNI743O1_18_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22110\,
            in1 => \N__36253\,
            in2 => \N__23031\,
            in3 => \N__36332\,
            lcout => OPEN,
            ltout => \un1_reset_rpi_inv_2_i_o3_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIRQR25_10_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22068\,
            in1 => \N__24972\,
            in2 => \N__22101\,
            in3 => \N__22185\,
            lcout => \N_1479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_3_0_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111010"
        )
    port map (
            in0 => \N__24508\,
            in1 => \N__24934\,
            in2 => \N__22098\,
            in3 => \N__29104\,
            lcout => g0_2_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_1_2_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__31280\,
            in1 => \N__32595\,
            in2 => \_gnd_net_\,
            in3 => \N__31363\,
            lcout => g1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNI6K4L_16_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36529\,
            in1 => \N__36654\,
            in2 => \N__35202\,
            in3 => \N__36430\,
            lcout => un1_reset_rpi_inv_2_i_o3_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_2_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__36934\,
            in1 => \N__36813\,
            in2 => \N__22062\,
            in3 => \N__24798\,
            lcout => g2_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_2_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22311\,
            in1 => \N__22323\,
            in2 => \N__22341\,
            in3 => \N__25185\,
            lcout => OPEN,
            ltout => \sbuttonModeStatus_0_sqmuxa_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__23013\,
            in1 => \N__22205\,
            in2 => \N__22218\,
            in3 => \N__25248\,
            lcout => \sbuttonModeStatusZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_1_1_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__24380\,
            in1 => \N__22194\,
            in2 => \N__24309\,
            in3 => \N__24719\,
            lcout => g1_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIOUF02_23_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37075\,
            in1 => \N__34452\,
            in2 => \N__23022\,
            in3 => \N__34574\,
            lcout => un1_reset_rpi_inv_2_i_o3_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIJ0NP_17_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36629\,
            in1 => \N__35163\,
            in2 => \N__36443\,
            in3 => \N__36805\,
            lcout => op_gt_op_gt_un13_striginternallto23_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_1_0_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__36806\,
            in1 => \N__36955\,
            in2 => \N__22179\,
            in3 => \N__24797\,
            lcout => g2_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_0_1_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32631\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31349\,
            lcout => OPEN,
            ltout => \g1_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_1_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010011010"
        )
    port map (
            in0 => \N__31262\,
            in1 => \N__22161\,
            in2 => \N__22155\,
            in3 => \N__22152\,
            lcout => \sTrigCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47829\,
            ce => 'H',
            sr => \N__27543\
        );

    \sCounter_RNIVUR25_10_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24987\,
            in1 => \N__22239\,
            in2 => \N__22146\,
            in3 => \N__22296\,
            lcout => op_gt_op_gt_un13_striginternal_0,
            ltout => \op_gt_op_gt_un13_striginternal_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigInternal_RNIMEFL5_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110101"
        )
    port map (
            in0 => \N__32633\,
            in1 => \N__22289\,
            in2 => \N__22137\,
            in3 => \N__24799\,
            lcout => \LED_ACQ_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIAME71_8_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35738\,
            in1 => \N__34454\,
            in2 => \N__34594\,
            in3 => \N__35849\,
            lcout => OPEN,
            ltout => \op_gt_op_gt_un13_striginternallto23_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIQVE02_16_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__36525\,
            in1 => \N__34700\,
            in2 => \N__22299\,
            in3 => \N__34834\,
            lcout => op_gt_op_gt_un13_striginternallto23_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LED_ACQ_obuf_RNO_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001100"
        )
    port map (
            in0 => \N__22290\,
            in1 => \N__32632\,
            in2 => \N__22269\,
            in3 => \N__24822\,
            lcout => \LED_ACQ_obuf_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNISQHJ1_18_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__25488\,
            in1 => \N__36228\,
            in2 => \N__24960\,
            in3 => \N__36309\,
            lcout => op_gt_op_gt_un13_striginternallto23_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterRAM_0_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22373\,
            in1 => \N__27392\,
            in2 => \_gnd_net_\,
            in3 => \N__22233\,
            lcout => \sCounterRAMZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \sCounterRAM_cry_0\,
            clk => \N__47845\,
            ce => 'H',
            sr => \N__53007\
        );

    \sCounterRAM_1_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22377\,
            in1 => \N__28013\,
            in2 => \_gnd_net_\,
            in3 => \N__22230\,
            lcout => \sCounterRAMZ0Z_1\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_0\,
            carryout => \sCounterRAM_cry_1\,
            clk => \N__47845\,
            ce => 'H',
            sr => \N__53007\
        );

    \sCounterRAM_2_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22374\,
            in1 => \N__28034\,
            in2 => \_gnd_net_\,
            in3 => \N__22227\,
            lcout => \sCounterRAMZ0Z_2\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_1\,
            carryout => \sCounterRAM_cry_2\,
            clk => \N__47845\,
            ce => 'H',
            sr => \N__53007\
        );

    \sCounterRAM_3_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22378\,
            in1 => \N__25307\,
            in2 => \_gnd_net_\,
            in3 => \N__22224\,
            lcout => \sCounterRAMZ0Z_3\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_2\,
            carryout => \sCounterRAM_cry_3\,
            clk => \N__47845\,
            ce => 'H',
            sr => \N__53007\
        );

    \sCounterRAM_4_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__22375\,
            in1 => \_gnd_net_\,
            in2 => \N__27437\,
            in3 => \N__22221\,
            lcout => \sCounterRAMZ0Z_4\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_3\,
            carryout => \sCounterRAM_cry_4\,
            clk => \N__47845\,
            ce => 'H',
            sr => \N__53007\
        );

    \sCounterRAM_5_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22379\,
            in1 => \N__27452\,
            in2 => \_gnd_net_\,
            in3 => \N__22386\,
            lcout => \sCounterRAMZ0Z_5\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_4\,
            carryout => \sCounterRAM_cry_5\,
            clk => \N__47845\,
            ce => 'H',
            sr => \N__53007\
        );

    \sCounterRAM_6_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22376\,
            in1 => \N__25323\,
            in2 => \_gnd_net_\,
            in3 => \N__22383\,
            lcout => \sCounterRAMZ0Z_6\,
            ltout => OPEN,
            carryin => \sCounterRAM_cry_5\,
            carryout => \sCounterRAM_cry_6\,
            clk => \N__47845\,
            ce => 'H',
            sr => \N__53007\
        );

    \sCounterRAM_7_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22380\,
            in1 => \N__27410\,
            in2 => \_gnd_net_\,
            in3 => \N__22350\,
            lcout => \sCounterRAMZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47845\,
            ce => 'H',
            sr => \N__53007\
        );

    \RAM_DATA_cl_10_15_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__31944\,
            in1 => \N__26610\,
            in2 => \N__32676\,
            in3 => \N__32177\,
            lcout => \RAM_DATA_cl_10Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47850\,
            ce => 'H',
            sr => \N__52999\
        );

    \sADC_clk_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__31943\,
            in1 => \N__27602\,
            in2 => \N__38229\,
            in3 => \N__32176\,
            lcout => \ADC_clk_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47850\,
            ce => 'H',
            sr => \N__52999\
        );

    \sSPI_MSB0LSB1_RNIO3VP1_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001100"
        )
    port map (
            in0 => \N__31693\,
            in1 => \N__27907\,
            in2 => \N__27980\,
            in3 => \N__31942\,
            lcout => \sSPI_MSB0LSB1_RNIO3VPZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_7_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23468\,
            in1 => \N__23483\,
            in2 => \N__23547\,
            in3 => \N__23498\,
            lcout => \sbuttonModeStatus_0_sqmuxa_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_5_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23336\,
            in1 => \N__23351\,
            in2 => \N__23322\,
            in3 => \N__23366\,
            lcout => \sbuttonModeStatus_0_sqmuxa_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_6_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23273\,
            in1 => \N__23288\,
            in2 => \N__23517\,
            in3 => \N__23303\,
            lcout => \sbuttonModeStatus_0_sqmuxa_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_14_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25704\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53246\,
            ce => 'H',
            sr => \N__53131\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_0_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28890\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53249\,
            ce => 'H',
            sr => \N__53122\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_8_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28866\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53249\,
            ce => 'H',
            sr => \N__53122\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_9_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28854\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53249\,
            ce => 'H',
            sr => \N__53122\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_7_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28878\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53249\,
            ce => 'H',
            sr => \N__53122\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_1_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25740\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53249\,
            ce => 'H',
            sr => \N__53122\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_13_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28752\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53249\,
            ce => 'H',
            sr => \N__53122\
        );

    \sPeriod_prev_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__36972\,
            in1 => \N__36877\,
            in2 => \_gnd_net_\,
            in3 => \N__24825\,
            lcout => \sPeriod_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47846\,
            ce => 'H',
            sr => \N__53107\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4Q_10_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23763\,
            in1 => \N__23586\,
            in2 => \_gnd_net_\,
            in3 => \N__22640\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4Q_12_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__22641\,
            in1 => \N__23571\,
            in2 => \_gnd_net_\,
            in3 => \N__23592\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_done_reg2_i_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28812\,
            lcout => \spi_slave_inst.rx_done_reg2_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47846\,
            ce => 'H',
            sr => \N__53107\
        );

    \spi_master_inst.sclk_gen_u0.falling_count_start_i_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__23643\,
            in1 => \N__23649\,
            in2 => \_gnd_net_\,
            in3 => \N__22555\,
            lcout => \spi_master_inst.sclk_gen_u0.falling_count_start_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53253\,
            ce => 'H',
            sr => \N__53093\
        );

    \spi_master_inst.sclk_gen_u0.spim_clk_state_i_2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__22556\,
            in1 => \N__23682\,
            in2 => \_gnd_net_\,
            in3 => \N__23750\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53253\,
            ce => 'H',
            sr => \N__53093\
        );

    \spi_master_inst.sclk_gen_u0.sclk_count_start_i_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__22557\,
            in1 => \N__22513\,
            in2 => \N__23739\,
            in3 => \N__22545\,
            lcout => \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53253\,
            ce => 'H',
            sr => \N__53093\
        );

    \spi_master_inst.sclk_gen_u0.delay_clk_i_RNISHDJ_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__22464\,
            in1 => \N__22493\,
            in2 => \_gnd_net_\,
            in3 => \N__23642\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.delay_clk_i_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22494\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_master_inst.sclk_gen_u0.delay_clk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53253\,
            ce => 'H',
            sr => \N__53093\
        );

    \sEETrigCounter_4_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49361\,
            lcout => \sEETrigCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47830\,
            ce => \N__31020\,
            sr => \N__53081\
        );

    \sEETrigCounter_5_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46970\,
            lcout => \sEETrigCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47830\,
            ce => \N__31020\,
            sr => \N__53081\
        );

    \sEETrigCounter_6_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48146\,
            lcout => \sEETrigCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47830\,
            ce => \N__31020\,
            sr => \N__53081\
        );

    \sEETrigCounter_7_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48736\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEETrigCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47830\,
            ce => \N__31020\,
            sr => \N__53081\
        );

    \sTrigCounter_RNO_2_2_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__36973\,
            in1 => \N__36848\,
            in2 => \N__22713\,
            in3 => \N__24818\,
            lcout => OPEN,
            ltout => \g2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_2_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100110"
        )
    port map (
            in0 => \N__24611\,
            in1 => \N__22704\,
            in2 => \N__22692\,
            in3 => \N__22689\,
            lcout => \sTrigCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47821\,
            ce => 'H',
            sr => \N__27542\
        );

    \sTrigCounter_RNO_0_2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__24357\,
            in1 => \N__24259\,
            in2 => \N__24714\,
            in3 => \N__24405\,
            lcout => g1_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_2_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__24817\,
            in1 => \N__22683\,
            in2 => \N__36873\,
            in3 => \N__36974\,
            lcout => OPEN,
            ltout => \g2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_3_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000110"
        )
    port map (
            in0 => \N__22674\,
            in1 => \N__24204\,
            in2 => \N__22677\,
            in3 => \N__22659\,
            lcout => \sTrigCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47821\,
            ce => 'H',
            sr => \N__27542\
        );

    \sTrigCounter_RNO_1_3_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24610\,
            in1 => \N__31300\,
            in2 => \N__32594\,
            in3 => \N__31388\,
            lcout => g1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_0_3_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__22665\,
            in1 => \N__24258\,
            in2 => \N__24376\,
            in3 => \N__24703\,
            lcout => g1_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_2_4_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__36959\,
            in1 => \N__36860\,
            in2 => \N__22653\,
            in3 => \N__24824\,
            lcout => OPEN,
            ltout => \g2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_4_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100110"
        )
    port map (
            in0 => \N__24230\,
            in1 => \N__24567\,
            in2 => \N__22812\,
            in3 => \N__22800\,
            lcout => \sTrigCounterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47813\,
            ce => 'H',
            sr => \N__27540\
        );

    \sTrigCounter_RNO_0_4_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__24377\,
            in1 => \N__22809\,
            in2 => \N__24314\,
            in3 => \N__24699\,
            lcout => g1_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_2_5_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__24823\,
            in1 => \N__22794\,
            in2 => \N__36878\,
            in3 => \N__36960\,
            lcout => OPEN,
            ltout => \g2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_5_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100110"
        )
    port map (
            in0 => \N__24651\,
            in1 => \N__22782\,
            in2 => \N__22776\,
            in3 => \N__24390\,
            lcout => \sTrigCounterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47813\,
            ce => 'H',
            sr => \N__27540\
        );

    \un4_speriod_cry_0_c_inv_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34230\,
            in2 => \N__22767\,
            in3 => \N__22773\,
            lcout => \sEEPeriod_i_0\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => un4_speriod_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_1_c_inv_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35058\,
            in2 => \N__22752\,
            in3 => \N__22758\,
            lcout => \sEEPeriod_i_1\,
            ltout => OPEN,
            carryin => un4_speriod_cry_0,
            carryout => un4_speriod_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_2_c_inv_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34957\,
            in2 => \N__22737\,
            in3 => \N__22743\,
            lcout => \sEEPeriod_i_2\,
            ltout => OPEN,
            carryin => un4_speriod_cry_1,
            carryout => un4_speriod_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_3_c_inv_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34852\,
            in2 => \N__22722\,
            in3 => \N__22728\,
            lcout => \sEEPeriod_i_3\,
            ltout => OPEN,
            carryin => un4_speriod_cry_2,
            carryout => un4_speriod_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_4_c_inv_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36855\,
            in2 => \N__22902\,
            in3 => \N__22908\,
            lcout => \sEEPeriod_i_4\,
            ltout => OPEN,
            carryin => un4_speriod_cry_3,
            carryout => un4_speriod_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_5_c_inv_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34710\,
            in2 => \N__22887\,
            in3 => \N__22893\,
            lcout => \sEEPeriod_i_5\,
            ltout => OPEN,
            carryin => un4_speriod_cry_4,
            carryout => un4_speriod_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_6_c_inv_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34605\,
            in2 => \N__22872\,
            in3 => \N__22878\,
            lcout => \sEEPeriod_i_6\,
            ltout => OPEN,
            carryin => un4_speriod_cry_5,
            carryout => un4_speriod_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_7_c_inv_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34479\,
            in2 => \N__22857\,
            in3 => \N__22863\,
            lcout => \sEEPeriod_i_7\,
            ltout => OPEN,
            carryin => un4_speriod_cry_6,
            carryout => un4_speriod_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_8_c_inv_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35877\,
            in2 => \N__22848\,
            in3 => \N__24999\,
            lcout => \sEEPeriod_i_8\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => un4_speriod_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_9_c_inv_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35762\,
            in2 => \N__22839\,
            in3 => \N__24993\,
            lcout => \sEEPeriod_i_9\,
            ltout => OPEN,
            carryin => un4_speriod_cry_8,
            carryout => un4_speriod_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_10_c_inv_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35647\,
            in2 => \N__22830\,
            in3 => \N__24561\,
            lcout => \sEEPeriod_i_10\,
            ltout => OPEN,
            carryin => un4_speriod_cry_9,
            carryout => un4_speriod_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_11_c_inv_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35532\,
            in2 => \N__22821\,
            in3 => \N__24555\,
            lcout => \sEEPeriod_i_11\,
            ltout => OPEN,
            carryin => un4_speriod_cry_10,
            carryout => un4_speriod_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_12_c_inv_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35410\,
            in2 => \N__23004\,
            in3 => \N__24549\,
            lcout => \sEEPeriod_i_12\,
            ltout => OPEN,
            carryin => un4_speriod_cry_11,
            carryout => un4_speriod_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_13_c_inv_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35306\,
            in2 => \N__22995\,
            in3 => \N__24543\,
            lcout => \sEEPeriod_i_13\,
            ltout => OPEN,
            carryin => un4_speriod_cry_12,
            carryout => un4_speriod_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_14_c_inv_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35195\,
            in2 => \N__22986\,
            in3 => \N__25011\,
            lcout => \sEEPeriod_i_14\,
            ltout => OPEN,
            carryin => un4_speriod_cry_13,
            carryout => un4_speriod_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_15_c_inv_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36637\,
            in2 => \N__22977\,
            in3 => \N__25005\,
            lcout => \sEEPeriod_i_15\,
            ltout => OPEN,
            carryin => un4_speriod_cry_14,
            carryout => un4_speriod_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_16_c_inv_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36531\,
            in2 => \N__22962\,
            in3 => \N__22968\,
            lcout => \sEEPeriod_i_16\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => un4_speriod_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_17_c_inv_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36426\,
            in2 => \N__22947\,
            in3 => \N__22953\,
            lcout => \sEEPeriod_i_17\,
            ltout => OPEN,
            carryin => un4_speriod_cry_16,
            carryout => un4_speriod_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_18_c_inv_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36345\,
            in2 => \N__22932\,
            in3 => \N__22938\,
            lcout => \sEEPeriod_i_18\,
            ltout => OPEN,
            carryin => un4_speriod_cry_17,
            carryout => un4_speriod_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_19_c_inv_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36252\,
            in2 => \N__22917\,
            in3 => \N__22923\,
            lcout => \sEEPeriod_i_19\,
            ltout => OPEN,
            carryin => un4_speriod_cry_18,
            carryout => un4_speriod_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_20_c_inv_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36162\,
            in2 => \N__23082\,
            in3 => \N__23088\,
            lcout => \sEEPeriod_i_20\,
            ltout => OPEN,
            carryin => un4_speriod_cry_19,
            carryout => un4_speriod_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_21_c_inv_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23067\,
            in2 => \N__36080\,
            in3 => \N__23073\,
            lcout => \sEEPeriod_i_21\,
            ltout => OPEN,
            carryin => un4_speriod_cry_20,
            carryout => un4_speriod_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_22_c_inv_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23055\,
            in2 => \N__35995\,
            in3 => \N__23061\,
            lcout => \sEEPeriod_i_22\,
            ltout => OPEN,
            carryin => un4_speriod_cry_21,
            carryout => un4_speriod_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_23_c_inv_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37074\,
            in2 => \N__23043\,
            in3 => \N__23049\,
            lcout => \sEEPeriod_i_23\,
            ltout => OPEN,
            carryin => un4_speriod_cry_22,
            carryout => un4_speriod_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_23_THRU_LUT4_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23034\,
            lcout => \un4_speriod_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNI3GS21_22_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34929\,
            in1 => \N__34201\,
            in2 => \N__35979\,
            in3 => \N__35024\,
            lcout => un1_reset_rpi_inv_2_i_o3_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNI5HE71_8_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35857\,
            in1 => \N__34695\,
            in2 => \N__35761\,
            in3 => \N__34827\,
            lcout => un1_reset_rpi_inv_2_i_o3_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23415\,
            in1 => \N__23436\,
            in2 => \N__23397\,
            in3 => \N__23454\,
            lcout => \sbuttonModeStatus_0_sqmuxa_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23244\,
            in1 => \N__34207\,
            in2 => \_gnd_net_\,
            in3 => \N__23007\,
            lcout => un7_spon_0,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \sCounter_cry_0\,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__53016\
        );

    \sCounter_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23223\,
            in1 => \N__35034\,
            in2 => \_gnd_net_\,
            in3 => \N__23115\,
            lcout => un7_spon_1,
            ltout => OPEN,
            carryin => \sCounter_cry_0\,
            carryout => \sCounter_cry_1\,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__53016\
        );

    \sCounter_2_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23245\,
            in1 => \N__34941\,
            in2 => \_gnd_net_\,
            in3 => \N__23112\,
            lcout => un7_spon_2,
            ltout => OPEN,
            carryin => \sCounter_cry_1\,
            carryout => \sCounter_cry_2\,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__53016\
        );

    \sCounter_3_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23224\,
            in1 => \N__34833\,
            in2 => \_gnd_net_\,
            in3 => \N__23109\,
            lcout => un7_spon_3,
            ltout => OPEN,
            carryin => \sCounter_cry_2\,
            carryout => \sCounter_cry_3\,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__53016\
        );

    \sCounter_4_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23246\,
            in1 => \N__36804\,
            in2 => \_gnd_net_\,
            in3 => \N__23106\,
            lcout => un7_spon_4,
            ltout => OPEN,
            carryin => \sCounter_cry_3\,
            carryout => \sCounter_cry_4\,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__53016\
        );

    \sCounter_5_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23225\,
            in1 => \N__34699\,
            in2 => \_gnd_net_\,
            in3 => \N__23103\,
            lcout => un7_spon_5,
            ltout => OPEN,
            carryin => \sCounter_cry_4\,
            carryout => \sCounter_cry_5\,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__53016\
        );

    \sCounter_6_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23247\,
            in1 => \N__34575\,
            in2 => \_gnd_net_\,
            in3 => \N__23100\,
            lcout => un7_spon_6,
            ltout => OPEN,
            carryin => \sCounter_cry_5\,
            carryout => \sCounter_cry_6\,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__53016\
        );

    \sCounter_7_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23226\,
            in1 => \N__34453\,
            in2 => \_gnd_net_\,
            in3 => \N__23097\,
            lcout => un7_spon_7,
            ltout => OPEN,
            carryin => \sCounter_cry_6\,
            carryout => \sCounter_cry_7\,
            clk => \N__47822\,
            ce => 'H',
            sr => \N__53016\
        );

    \sCounter_8_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23218\,
            in1 => \N__35850\,
            in2 => \_gnd_net_\,
            in3 => \N__23094\,
            lcout => un7_spon_8,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \sCounter_cry_8\,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__53008\
        );

    \sCounter_9_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23230\,
            in1 => \N__35739\,
            in2 => \_gnd_net_\,
            in3 => \N__23091\,
            lcout => un7_spon_9,
            ltout => OPEN,
            carryin => \sCounter_cry_8\,
            carryout => \sCounter_cry_9\,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__53008\
        );

    \sCounter_10_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23215\,
            in1 => \N__35627\,
            in2 => \_gnd_net_\,
            in3 => \N__23142\,
            lcout => un7_spon_10,
            ltout => OPEN,
            carryin => \sCounter_cry_9\,
            carryout => \sCounter_cry_10\,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__53008\
        );

    \sCounter_11_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23227\,
            in1 => \N__35516\,
            in2 => \_gnd_net_\,
            in3 => \N__23139\,
            lcout => un7_spon_11,
            ltout => OPEN,
            carryin => \sCounter_cry_10\,
            carryout => \sCounter_cry_11\,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__53008\
        );

    \sCounter_12_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23216\,
            in1 => \N__35379\,
            in2 => \_gnd_net_\,
            in3 => \N__23136\,
            lcout => un7_spon_12,
            ltout => OPEN,
            carryin => \sCounter_cry_11\,
            carryout => \sCounter_cry_12\,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__53008\
        );

    \sCounter_13_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23228\,
            in1 => \N__35291\,
            in2 => \_gnd_net_\,
            in3 => \N__23133\,
            lcout => un7_spon_13,
            ltout => OPEN,
            carryin => \sCounter_cry_12\,
            carryout => \sCounter_cry_13\,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__53008\
        );

    \sCounter_14_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23217\,
            in1 => \N__35164\,
            in2 => \_gnd_net_\,
            in3 => \N__23130\,
            lcout => un7_spon_14,
            ltout => OPEN,
            carryin => \sCounter_cry_13\,
            carryout => \sCounter_cry_14\,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__53008\
        );

    \sCounter_15_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23229\,
            in1 => \N__36633\,
            in2 => \_gnd_net_\,
            in3 => \N__23127\,
            lcout => un7_spon_15,
            ltout => OPEN,
            carryin => \sCounter_cry_14\,
            carryout => \sCounter_cry_15\,
            clk => \N__47831\,
            ce => 'H',
            sr => \N__53008\
        );

    \sCounter_16_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23240\,
            in1 => \N__36521\,
            in2 => \_gnd_net_\,
            in3 => \N__23124\,
            lcout => un7_spon_16,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \sCounter_cry_16\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__53000\
        );

    \sCounter_17_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23219\,
            in1 => \N__36405\,
            in2 => \_gnd_net_\,
            in3 => \N__23121\,
            lcout => un7_spon_17,
            ltout => OPEN,
            carryin => \sCounter_cry_16\,
            carryout => \sCounter_cry_17\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__53000\
        );

    \sCounter_18_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23241\,
            in1 => \N__36327\,
            in2 => \_gnd_net_\,
            in3 => \N__23118\,
            lcout => un7_spon_18,
            ltout => OPEN,
            carryin => \sCounter_cry_17\,
            carryout => \sCounter_cry_18\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__53000\
        );

    \sCounter_19_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23220\,
            in1 => \N__36229\,
            in2 => \_gnd_net_\,
            in3 => \N__23259\,
            lcout => un7_spon_19,
            ltout => OPEN,
            carryin => \sCounter_cry_18\,
            carryout => \sCounter_cry_19\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__53000\
        );

    \sCounter_20_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23242\,
            in1 => \N__36136\,
            in2 => \_gnd_net_\,
            in3 => \N__23256\,
            lcout => un7_spon_20,
            ltout => OPEN,
            carryin => \sCounter_cry_19\,
            carryout => \sCounter_cry_20\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__53000\
        );

    \sCounter_21_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23221\,
            in1 => \N__36064\,
            in2 => \_gnd_net_\,
            in3 => \N__23253\,
            lcout => un7_spon_21,
            ltout => OPEN,
            carryin => \sCounter_cry_20\,
            carryout => \sCounter_cry_21\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__53000\
        );

    \sCounter_22_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23243\,
            in1 => \N__35950\,
            in2 => \_gnd_net_\,
            in3 => \N__23250\,
            lcout => un7_spon_22,
            ltout => OPEN,
            carryin => \sCounter_cry_21\,
            carryout => \sCounter_cry_22\,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__53000\
        );

    \sCounter_23_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__23222\,
            in1 => \N__37053\,
            in2 => \_gnd_net_\,
            in3 => \N__23154\,
            lcout => un7_spon_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47838\,
            ce => 'H',
            sr => \N__53000\
        );

    \sbuttonModeStatus_RNO_3_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26274\,
            in2 => \N__26313\,
            in3 => \N__32500\,
            lcout => \sbuttonModeStatus_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => un1_button_debounce_counter_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \button_debounce_counter_2_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32496\,
            in1 => \N__25197\,
            in2 => \_gnd_net_\,
            in3 => \N__23151\,
            lcout => \button_debounce_counterZ0Z_2\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_1,
            carryout => un1_button_debounce_counter_cry_2,
            clk => \N__53280\,
            ce => 'H',
            sr => \N__26240\
        );

    \button_debounce_counter_3_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32634\,
            in1 => \N__25224\,
            in2 => \_gnd_net_\,
            in3 => \N__23148\,
            lcout => \button_debounce_counterZ0Z_3\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_2,
            carryout => un1_button_debounce_counter_cry_3,
            clk => \N__53280\,
            ce => 'H',
            sr => \N__26240\
        );

    \button_debounce_counter_4_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32497\,
            in1 => \N__25236\,
            in2 => \_gnd_net_\,
            in3 => \N__23145\,
            lcout => \button_debounce_counterZ0Z_4\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_3,
            carryout => un1_button_debounce_counter_cry_4,
            clk => \N__53280\,
            ce => 'H',
            sr => \N__26240\
        );

    \button_debounce_counter_5_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32635\,
            in1 => \N__25211\,
            in2 => \_gnd_net_\,
            in3 => \N__23370\,
            lcout => \button_debounce_counterZ0Z_5\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_4,
            carryout => un1_button_debounce_counter_cry_5,
            clk => \N__53280\,
            ce => 'H',
            sr => \N__26240\
        );

    \button_debounce_counter_6_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32498\,
            in1 => \N__23367\,
            in2 => \_gnd_net_\,
            in3 => \N__23355\,
            lcout => \button_debounce_counterZ0Z_6\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_5,
            carryout => un1_button_debounce_counter_cry_6,
            clk => \N__53280\,
            ce => 'H',
            sr => \N__26240\
        );

    \button_debounce_counter_7_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32636\,
            in1 => \N__23352\,
            in2 => \_gnd_net_\,
            in3 => \N__23340\,
            lcout => \button_debounce_counterZ0Z_7\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_6,
            carryout => un1_button_debounce_counter_cry_7,
            clk => \N__53280\,
            ce => 'H',
            sr => \N__26240\
        );

    \button_debounce_counter_8_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32499\,
            in1 => \N__23337\,
            in2 => \_gnd_net_\,
            in3 => \N__23325\,
            lcout => \button_debounce_counterZ0Z_8\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_7,
            carryout => un1_button_debounce_counter_cry_8,
            clk => \N__53280\,
            ce => 'H',
            sr => \N__26240\
        );

    \button_debounce_counter_9_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32684\,
            in1 => \N__23321\,
            in2 => \_gnd_net_\,
            in3 => \N__23307\,
            lcout => \button_debounce_counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => un1_button_debounce_counter_cry_9,
            clk => \N__53281\,
            ce => 'H',
            sr => \N__26241\
        );

    \button_debounce_counter_10_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32677\,
            in1 => \N__23304\,
            in2 => \_gnd_net_\,
            in3 => \N__23292\,
            lcout => \button_debounce_counterZ0Z_10\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_9,
            carryout => un1_button_debounce_counter_cry_10,
            clk => \N__53281\,
            ce => 'H',
            sr => \N__26241\
        );

    \button_debounce_counter_11_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32681\,
            in1 => \N__23289\,
            in2 => \_gnd_net_\,
            in3 => \N__23277\,
            lcout => \button_debounce_counterZ0Z_11\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_10,
            carryout => un1_button_debounce_counter_cry_11,
            clk => \N__53281\,
            ce => 'H',
            sr => \N__26241\
        );

    \button_debounce_counter_12_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32678\,
            in1 => \N__23274\,
            in2 => \_gnd_net_\,
            in3 => \N__23262\,
            lcout => \button_debounce_counterZ0Z_12\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_11,
            carryout => un1_button_debounce_counter_cry_12,
            clk => \N__53281\,
            ce => 'H',
            sr => \N__26241\
        );

    \button_debounce_counter_13_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32682\,
            in1 => \N__23516\,
            in2 => \_gnd_net_\,
            in3 => \N__23502\,
            lcout => \button_debounce_counterZ0Z_13\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_12,
            carryout => un1_button_debounce_counter_cry_13,
            clk => \N__53281\,
            ce => 'H',
            sr => \N__26241\
        );

    \button_debounce_counter_14_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32679\,
            in1 => \N__23499\,
            in2 => \_gnd_net_\,
            in3 => \N__23487\,
            lcout => \button_debounce_counterZ0Z_14\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_13,
            carryout => un1_button_debounce_counter_cry_14,
            clk => \N__53281\,
            ce => 'H',
            sr => \N__26241\
        );

    \button_debounce_counter_15_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32683\,
            in1 => \N__23484\,
            in2 => \_gnd_net_\,
            in3 => \N__23472\,
            lcout => \button_debounce_counterZ0Z_15\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_14,
            carryout => un1_button_debounce_counter_cry_15,
            clk => \N__53281\,
            ce => 'H',
            sr => \N__26241\
        );

    \button_debounce_counter_16_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32680\,
            in1 => \N__23469\,
            in2 => \_gnd_net_\,
            in3 => \N__23457\,
            lcout => \button_debounce_counterZ0Z_16\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_15,
            carryout => un1_button_debounce_counter_cry_16,
            clk => \N__53281\,
            ce => 'H',
            sr => \N__26241\
        );

    \button_debounce_counter_17_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32685\,
            in1 => \N__23450\,
            in2 => \_gnd_net_\,
            in3 => \N__23439\,
            lcout => \button_debounce_counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => un1_button_debounce_counter_cry_17,
            clk => \N__53282\,
            ce => 'H',
            sr => \N__26242\
        );

    \button_debounce_counter_18_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32688\,
            in1 => \N__23429\,
            in2 => \_gnd_net_\,
            in3 => \N__23418\,
            lcout => \button_debounce_counterZ0Z_18\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_17,
            carryout => un1_button_debounce_counter_cry_18,
            clk => \N__53282\,
            ce => 'H',
            sr => \N__26242\
        );

    \button_debounce_counter_19_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32686\,
            in1 => \N__23411\,
            in2 => \_gnd_net_\,
            in3 => \N__23400\,
            lcout => \button_debounce_counterZ0Z_19\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_18,
            carryout => un1_button_debounce_counter_cry_19,
            clk => \N__53282\,
            ce => 'H',
            sr => \N__26242\
        );

    \button_debounce_counter_20_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32689\,
            in1 => \N__23387\,
            in2 => \_gnd_net_\,
            in3 => \N__23376\,
            lcout => \button_debounce_counterZ0Z_20\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_19,
            carryout => un1_button_debounce_counter_cry_20,
            clk => \N__53282\,
            ce => 'H',
            sr => \N__26242\
        );

    \button_debounce_counter_21_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32687\,
            in1 => \N__25286\,
            in2 => \_gnd_net_\,
            in3 => \N__23373\,
            lcout => \button_debounce_counterZ0Z_21\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_20,
            carryout => un1_button_debounce_counter_cry_21,
            clk => \N__53282\,
            ce => 'H',
            sr => \N__26242\
        );

    \button_debounce_counter_22_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32690\,
            in1 => \N__25265\,
            in2 => \_gnd_net_\,
            in3 => \N__23553\,
            lcout => \button_debounce_counterZ0Z_22\,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_21,
            carryout => un1_button_debounce_counter_cry_22,
            clk => \N__53282\,
            ce => 'H',
            sr => \N__26242\
        );

    \un1_button_debounce_counter_cry_22_c_THRU_CRY_0_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38020\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_button_debounce_counter_cry_22,
            carryout => \un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_button_debounce_counter_cry_22_c_THRU_CRY_1_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__38068\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO\,
            carryout => \un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \button_debounce_counter_esr_23_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23543\,
            in2 => \_gnd_net_\,
            in3 => \N__23550\,
            lcout => \button_debounce_counterZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53283\,
            ce => \N__25470\,
            sr => \N__26243\
        );

    \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_c_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25552\,
            in2 => \N__25503\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_3_0_\,
            carryout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_LUT4_0_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25574\,
            in2 => \_gnd_net_\,
            in3 => \N__23529\,
            lcout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0\,
            carryout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_LUT4_0_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25774\,
            in2 => \_gnd_net_\,
            in3 => \N__23526\,
            lcout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1\,
            carryout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_3_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25590\,
            in2 => \_gnd_net_\,
            in3 => \N__23523\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2\,
            carryout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3\,
            clk => \N__30703\,
            ce => 'H',
            sr => \N__53123\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_4_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25533\,
            in2 => \_gnd_net_\,
            in3 => \N__23520\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3\,
            carryout => \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4\,
            clk => \N__30703\,
            ce => 'H',
            sr => \N__53123\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_5_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25796\,
            in2 => \_gnd_net_\,
            in3 => \N__23607\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30703\,
            ce => 'H',
            sr => \N__53123\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_1_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010100000111100"
        )
    port map (
            in0 => \N__33222\,
            in1 => \N__23604\,
            in2 => \N__25578\,
            in3 => \N__25517\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30705\,
            ce => 'H',
            sr => \N__53108\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_2_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101110110000"
        )
    port map (
            in0 => \N__33223\,
            in1 => \N__25518\,
            in2 => \N__25779\,
            in3 => \N__23598\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30705\,
            ce => 'H',
            sr => \N__53108\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_0_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000010100"
        )
    port map (
            in0 => \N__25516\,
            in1 => \N__25502\,
            in2 => \N__25557\,
            in3 => \N__33221\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30705\,
            ce => 'H',
            sr => \N__53108\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_12_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25716\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53250\,
            ce => 'H',
            sr => \N__53094\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_2_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25728\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53250\,
            ce => 'H',
            sr => \N__53094\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_3_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25710\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53250\,
            ce => 'H',
            sr => \N__53094\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_4_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28737\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53250\,
            ce => 'H',
            sr => \N__53094\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_5_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28728\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53250\,
            ce => 'H',
            sr => \N__53094\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_15_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25986\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53250\,
            ce => 'H',
            sr => \N__53094\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_11_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25722\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53250\,
            ce => 'H',
            sr => \N__53094\
        );

    \spi_master_inst.spi_data_path_u1.txdata_reg_i_10_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28761\,
            lcout => \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53250\,
            ce => 'H',
            sr => \N__53094\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNISEQE3_1_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__25964\,
            in1 => \N__24072\,
            in2 => \N__25947\,
            in3 => \N__23613\,
            lcout => \spi_master_inst.sclk_gen_u0.N_158_7\,
            ltout => \spi_master_inst.sclk_gen_u0.N_158_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNO_0_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__23735\,
            in1 => \N__26994\,
            in2 => \N__23697\,
            in3 => \N__23678\,
            lcout => \spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNIK09A_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23641\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_master_inst.sclk_gen_u0.falling_count_start_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_ft_ibuf_RNI4OFN_1_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__24065\,
            in1 => \N__23978\,
            in2 => \_gnd_net_\,
            in3 => \N__23877\,
            lcout => un3_trig_0_0,
            ltout => \un3_trig_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_3_5_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111010"
        )
    port map (
            in0 => \N__24506\,
            in1 => \N__24941\,
            in2 => \N__23616\,
            in3 => \N__29093\,
            lcout => g1_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNIKGMR_0_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25913\,
            in2 => \_gnd_net_\,
            in3 => \N__25979\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNILEDN1_7_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25898\,
            in1 => \N__25829\,
            in2 => \N__25884\,
            in3 => \N__25928\,
            lcout => \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_ft_ibuf_RNI4OFN_4_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__24066\,
            in1 => \N__23979\,
            in2 => \_gnd_net_\,
            in3 => \N__23878\,
            lcout => un3_trig_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNINQ4B1_2_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__26013\,
            in1 => \_gnd_net_\,
            in2 => \N__26082\,
            in3 => \N__26111\,
            lcout => OPEN,
            ltout => \un8_trig_prev_0_c5_a0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNII5M43_6_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001101100"
        )
    port map (
            in0 => \N__24163\,
            in1 => \N__23808\,
            in2 => \N__23826\,
            in3 => \N__23820\,
            lcout => un10_trig_prev_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIHO9M2_5_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101010101010"
        )
    port map (
            in0 => \N__23819\,
            in1 => \N__26116\,
            in2 => \N__24165\,
            in3 => \N__23789\,
            lcout => un10_trig_prev_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIPGOS_2_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26012\,
            in2 => \_gnd_net_\,
            in3 => \N__26076\,
            lcout => un8_trig_prev_0_c4_a0_1,
            ltout => \un8_trig_prev_0_c4_a0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIHCT72_4_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100010000"
        )
    port map (
            in0 => \N__26036\,
            in1 => \N__26115\,
            in2 => \N__23823\,
            in3 => \N__24176\,
            lcout => un10_trig_prev_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIV25B1_6_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23818\,
            in2 => \N__26120\,
            in3 => \N__23807\,
            lcout => OPEN,
            ltout => \un8_trig_prev_0_c7_a0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIKJ2J3_7_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__23799\,
            in1 => \N__24164\,
            in2 => \N__23793\,
            in3 => \N__23790\,
            lcout => un10_trig_prev_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIQHOS_4_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24177\,
            in3 => \N__26035\,
            lcout => un8_trig_prev_0_c5_a0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_0_c_inv_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24147\,
            in2 => \N__26055\,
            in3 => \N__31379\,
            lcout => \sTrigCounter_i_0\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => un10_trig_prev_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_1_c_inv_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24141\,
            in2 => \N__25995\,
            in3 => \N__31298\,
            lcout => \sTrigCounter_i_1\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_0,
            carryout => un10_trig_prev_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_2_c_inv_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26061\,
            in2 => \N__24135\,
            in3 => \N__24612\,
            lcout => \sTrigCounter_i_2\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_1,
            carryout => un10_trig_prev_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_3_c_inv_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24200\,
            in1 => \N__24126\,
            in2 => \N__26094\,
            in3 => \_gnd_net_\,
            lcout => \sTrigCounter_i_3\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_2,
            carryout => un10_trig_prev_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_4_c_inv_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24231\,
            in1 => \N__24111\,
            in2 => \N__24120\,
            in3 => \_gnd_net_\,
            lcout => \sTrigCounter_i_4\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_3,
            carryout => un10_trig_prev_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_5_c_inv_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24096\,
            in2 => \N__24105\,
            in3 => \N__24645\,
            lcout => \sTrigCounter_i_5\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_4,
            carryout => un10_trig_prev_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_6_c_inv_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25076\,
            in1 => \N__24081\,
            in2 => \N__24090\,
            in3 => \_gnd_net_\,
            lcout => \sTrigCounter_i_6\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_5,
            carryout => un10_trig_prev_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_7_c_inv_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24528\,
            in2 => \N__24537\,
            in3 => \N__25032\,
            lcout => \sTrigCounter_i_7\,
            ltout => OPEN,
            carryin => un10_trig_prev_cry_6,
            carryout => un10_trig_prev_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un10_trig_prev_cry_7_THRU_LUT4_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24522\,
            lcout => \un10_trig_prev_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_1_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__46451\,
            in1 => \N__31106\,
            in2 => \N__44478\,
            in3 => \N__44745\,
            lcout => \sAddress_RNI9IH12_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_3_2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111010"
        )
    port map (
            in0 => \N__24510\,
            in1 => \N__24943\,
            in2 => \N__24428\,
            in3 => \N__29084\,
            lcout => g1_0_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_0_5_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__24273\,
            in1 => \N__24378\,
            in2 => \N__24713\,
            in3 => \N__24399\,
            lcout => g1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_0_7_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__24379\,
            in1 => \N__24272\,
            in2 => \N__27576\,
            in3 => \N__24694\,
            lcout => \N_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNI9UM4_4_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24228\,
            in2 => \_gnd_net_\,
            in3 => \N__24201\,
            lcout => \un1_sTrigCounter_ac0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_4_4_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32562\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24202\,
            lcout => g1_0_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_2_6_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31293\,
            in2 => \_gnd_net_\,
            in3 => \N__31390\,
            lcout => OPEN,
            ltout => \un1_sTrigCounter_ac0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_1_6_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24626\,
            in1 => \N__24646\,
            in2 => \N__24744\,
            in3 => \N__24613\,
            lcout => OPEN,
            ltout => \un1_sTrigCounter_ac0_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_0_6_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001010000"
        )
    port map (
            in0 => \N__27568\,
            in1 => \N__24741\,
            in2 => \N__24723\,
            in3 => \N__24698\,
            lcout => \un1_sTrigCounter_ac0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_2_7_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__31391\,
            in1 => \_gnd_net_\,
            in2 => \N__31302\,
            in3 => \N__24614\,
            lcout => OPEN,
            ltout => \un1_sTrigCounter_ac0_3_out_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_1_7_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24647\,
            in1 => \N__24627\,
            in2 => \N__24618\,
            in3 => \N__25077\,
            lcout => \un1_sTrigCounter_axbxc7_m7_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_RNO_1_4_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24615\,
            in1 => \N__31297\,
            in2 => \N__24576\,
            in3 => \N__31392\,
            lcout => g1_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPeriod_10_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50281\,
            lcout => \sEEPeriodZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47776\,
            ce => \N__28944\,
            sr => \N__53028\
        );

    \sEEPeriod_11_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49785\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47776\,
            ce => \N__28944\,
            sr => \N__53028\
        );

    \sEEPeriod_12_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49367\,
            lcout => \sEEPeriodZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47776\,
            ce => \N__28944\,
            sr => \N__53028\
        );

    \sEEPeriod_13_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47062\,
            lcout => \sEEPeriodZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47776\,
            ce => \N__28944\,
            sr => \N__53028\
        );

    \sEEPeriod_14_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48244\,
            lcout => \sEEPeriodZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47776\,
            ce => \N__28944\,
            sr => \N__53028\
        );

    \sEEPeriod_15_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48633\,
            lcout => \sEEPeriodZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47776\,
            ce => \N__28944\,
            sr => \N__53028\
        );

    \sEEPeriod_8_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51139\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPeriodZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47776\,
            ce => \N__28944\,
            sr => \N__53028\
        );

    \sEEPeriod_9_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50665\,
            lcout => \sEEPeriodZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47776\,
            ce => \N__28944\,
            sr => \N__53028\
        );

    \sCounter_RNIM34L_0_10_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35522\,
            in1 => \N__35298\,
            in2 => \N__35396\,
            in3 => \N__35632\,
            lcout => op_gt_op_gt_un13_striginternallto23_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIM34L_10_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35631\,
            in1 => \N__35380\,
            in2 => \N__35310\,
            in3 => \N__35521\,
            lcout => un1_reset_rpi_inv_2_i_o3_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIO6BU_23_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35981\,
            in1 => \N__34949\,
            in2 => \N__37089\,
            in3 => \N__35050\,
            lcout => op_gt_op_gt_un13_striginternallto23_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_speriod_cry_23_c_RNIHTOK1_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010110000"
        )
    port map (
            in0 => \N__24944\,
            in1 => \N__29060\,
            in2 => \N__24843\,
            in3 => \N__24790\,
            lcout => OPEN,
            ltout => \un1_reset_rpi_inv_2_i_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIT8E57_4_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111010101"
        )
    port map (
            in0 => \N__32547\,
            in1 => \N__36957\,
            in2 => \N__24747\,
            in3 => \N__36844\,
            lcout => un1_reset_rpi_inv_2_i_1,
            ltout => \un1_reset_rpi_inv_2_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sTrigCounter_6_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25075\,
            in2 => \N__25089\,
            in3 => \N__25086\,
            lcout => \sTrigCounterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47790\,
            ce => 'H',
            sr => \N__27536\
        );

    \sTrigCounter_7_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010010"
        )
    port map (
            in0 => \N__25056\,
            in1 => \N__25047\,
            in2 => \N__25031\,
            in3 => \N__25041\,
            lcout => \sTrigCounterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47790\,
            ce => 'H',
            sr => \N__27536\
        );

    \un1_spoff_cry_0_c_inv_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29316\,
            in2 => \N__26169\,
            in3 => \N__34200\,
            lcout => \sCounter_i_0\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => un1_spoff_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_1_c_inv_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26151\,
            in2 => \N__29307\,
            in3 => \N__35023\,
            lcout => \sCounter_i_1\,
            ltout => OPEN,
            carryin => un1_spoff_cry_0,
            carryout => un1_spoff_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_2_c_inv_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29292\,
            in2 => \N__26460\,
            in3 => \N__34925\,
            lcout => \sCounter_i_2\,
            ltout => OPEN,
            carryin => un1_spoff_cry_1,
            carryout => un1_spoff_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_3_c_inv_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29283\,
            in2 => \N__26442\,
            in3 => \N__34817\,
            lcout => \sCounter_i_3\,
            ltout => OPEN,
            carryin => un1_spoff_cry_2,
            carryout => un1_spoff_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_4_c_inv_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29274\,
            in2 => \N__26424\,
            in3 => \N__36782\,
            lcout => \sCounter_i_4\,
            ltout => OPEN,
            carryin => un1_spoff_cry_3,
            carryout => un1_spoff_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_5_c_inv_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29265\,
            in2 => \N__26406\,
            in3 => \N__34691\,
            lcout => \sCounter_i_5\,
            ltout => OPEN,
            carryin => un1_spoff_cry_4,
            carryout => un1_spoff_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_6_c_inv_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29256\,
            in2 => \N__26388\,
            in3 => \N__34567\,
            lcout => \sCounter_i_6\,
            ltout => OPEN,
            carryin => un1_spoff_cry_5,
            carryout => un1_spoff_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_7_c_inv_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34445\,
            in1 => \N__29247\,
            in2 => \N__26370\,
            in3 => \_gnd_net_\,
            lcout => \sCounter_i_7\,
            ltout => OPEN,
            carryin => un1_spoff_cry_6,
            carryout => un1_spoff_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_8_c_inv_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29355\,
            in2 => \N__26349\,
            in3 => \N__35842\,
            lcout => \sCounter_i_8\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => un1_spoff_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_9_c_inv_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29346\,
            in2 => \N__26331\,
            in3 => \N__35731\,
            lcout => \sCounter_i_9\,
            ltout => OPEN,
            carryin => un1_spoff_cry_8,
            carryout => un1_spoff_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_10_c_inv_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29238\,
            in2 => \N__26583\,
            in3 => \N__35617\,
            lcout => \sCounter_i_10\,
            ltout => OPEN,
            carryin => un1_spoff_cry_9,
            carryout => un1_spoff_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_11_c_inv_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29409\,
            in2 => \N__26565\,
            in3 => \N__35496\,
            lcout => \sCounter_i_11\,
            ltout => OPEN,
            carryin => un1_spoff_cry_10,
            carryout => un1_spoff_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_12_c_inv_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29397\,
            in2 => \N__26547\,
            in3 => \N__35369\,
            lcout => \sCounter_i_12\,
            ltout => OPEN,
            carryin => un1_spoff_cry_11,
            carryout => un1_spoff_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_13_c_inv_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29385\,
            in2 => \N__26529\,
            in3 => \N__35284\,
            lcout => \sCounter_i_13\,
            ltout => OPEN,
            carryin => un1_spoff_cry_12,
            carryout => un1_spoff_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_14_c_inv_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29376\,
            in2 => \N__26511\,
            in3 => \N__35156\,
            lcout => \sCounter_i_14\,
            ltout => OPEN,
            carryin => un1_spoff_cry_13,
            carryout => un1_spoff_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_15_c_inv_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26492\,
            in2 => \N__29367\,
            in3 => \N__36616\,
            lcout => \sCounter_i_15\,
            ltout => OPEN,
            carryin => un1_spoff_cry_14,
            carryout => un1_spoff_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_16_c_inv_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25137\,
            in2 => \_gnd_net_\,
            in3 => \N__36507\,
            lcout => \sCounter_i_16\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => un1_spoff_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_17_c_inv_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36406\,
            in1 => \N__25131\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sCounter_i_17\,
            ltout => OPEN,
            carryin => un1_spoff_cry_16,
            carryout => un1_spoff_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_18_c_inv_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36310\,
            in1 => \N__25125\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sCounter_i_18\,
            ltout => OPEN,
            carryin => un1_spoff_cry_17,
            carryout => un1_spoff_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_19_c_inv_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25119\,
            in2 => \_gnd_net_\,
            in3 => \N__36230\,
            lcout => \sCounter_i_19\,
            ltout => OPEN,
            carryin => un1_spoff_cry_18,
            carryout => un1_spoff_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_20_c_inv_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25113\,
            in2 => \_gnd_net_\,
            in3 => \N__36137\,
            lcout => \sCounter_i_20\,
            ltout => OPEN,
            carryin => un1_spoff_cry_19,
            carryout => un1_spoff_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_21_c_inv_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25107\,
            in2 => \_gnd_net_\,
            in3 => \N__36053\,
            lcout => \sCounter_i_21\,
            ltout => OPEN,
            carryin => un1_spoff_cry_20,
            carryout => un1_spoff_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_22_c_inv_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35951\,
            in1 => \N__25101\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sCounter_i_22\,
            ltout => OPEN,
            carryin => un1_spoff_cry_21,
            carryout => un1_spoff_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_spoff_cry_23_c_inv_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25095\,
            in2 => \_gnd_net_\,
            in3 => \N__37054\,
            lcout => \sCounter_i_23\,
            ltout => OPEN,
            carryin => un1_spoff_cry_22,
            carryout => un1_spoff_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \poff_obuf_RNO_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25350\,
            in2 => \_gnd_net_\,
            in3 => \N__25338\,
            lcout => \N_1612_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sRead_data_RNI74VQ_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__27474\,
            in1 => \N__25322\,
            in2 => \_gnd_net_\,
            in3 => \N__25308\,
            lcout => spi_data_miso_0_sqmuxa_2_i_o2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_1_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26309\,
            in1 => \N__25293\,
            in2 => \N__25275\,
            in3 => \N__25254\,
            lcout => \sbuttonModeStatus_0_sqmuxa_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sbuttonModeStatus_RNO_4_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25235\,
            in1 => \N__25223\,
            in2 => \N__25212\,
            in3 => \N__25196\,
            lcout => \sbuttonModeStatus_0_sqmuxa_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_0_c_inv_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34226\,
            in2 => \N__25173\,
            in3 => \N__26739\,
            lcout => \sEEDelayACQ_i_0\,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => un4_sacqtime_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_1_c_inv_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35051\,
            in2 => \N__25164\,
            in3 => \N__26733\,
            lcout => \sEEDelayACQ_i_1\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_0,
            carryout => un4_sacqtime_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_2_c_inv_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34942\,
            in2 => \N__25155\,
            in3 => \N__26727\,
            lcout => \sEEDelayACQ_i_2\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_1,
            carryout => un4_sacqtime_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_3_c_inv_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34835\,
            in2 => \N__25146\,
            in3 => \N__26721\,
            lcout => \sEEDelayACQ_i_3\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_2,
            carryout => un4_sacqtime_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_4_c_inv_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26715\,
            in1 => \N__36819\,
            in2 => \N__25419\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQ_i_4\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_3,
            carryout => un4_sacqtime_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_5_c_inv_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34706\,
            in2 => \N__25410\,
            in3 => \N__26709\,
            lcout => \sEEDelayACQ_i_5\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_4,
            carryout => un4_sacqtime_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_6_c_inv_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34601\,
            in2 => \N__25401\,
            in3 => \N__26808\,
            lcout => \sEEDelayACQ_i_6\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_5,
            carryout => un4_sacqtime_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_7_c_inv_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26802\,
            in1 => \N__25392\,
            in2 => \N__34475\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQ_i_7\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_6,
            carryout => un4_sacqtime_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_8_c_inv_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35870\,
            in2 => \N__25386\,
            in3 => \N__26760\,
            lcout => \sEEDelayACQ_i_8\,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => un4_sacqtime_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_9_c_inv_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35768\,
            in2 => \N__25377\,
            in3 => \N__26952\,
            lcout => \sEEDelayACQ_i_9\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_8,
            carryout => un4_sacqtime_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_10_c_inv_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35633\,
            in2 => \N__25368\,
            in3 => \N__26796\,
            lcout => \sEEDelayACQ_i_10\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_9,
            carryout => un4_sacqtime_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_11_c_inv_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35520\,
            in2 => \N__25359\,
            in3 => \N__26790\,
            lcout => \sEEDelayACQ_i_11\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_10,
            carryout => un4_sacqtime_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_12_c_inv_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35384\,
            in2 => \N__25452\,
            in3 => \N__26784\,
            lcout => \sEEDelayACQ_i_12\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_11,
            carryout => un4_sacqtime_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_13_c_inv_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35302\,
            in2 => \N__25443\,
            in3 => \N__26778\,
            lcout => \sEEDelayACQ_i_13\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_12,
            carryout => un4_sacqtime_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_14_c_inv_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35188\,
            in2 => \N__25434\,
            in3 => \N__26772\,
            lcout => \sEEDelayACQ_i_14\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_13,
            carryout => un4_sacqtime_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_15_c_inv_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25425\,
            in2 => \N__36653\,
            in3 => \N__26766\,
            lcout => \sEEDelayACQ_i_15\,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_14,
            carryout => un4_sacqtime_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_16_c_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36530\,
            in2 => \N__38072\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => un4_sacqtime_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_17_c_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36431\,
            in2 => \N__38070\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_16,
            carryout => un4_sacqtime_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_18_c_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36328\,
            in2 => \N__38073\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_17,
            carryout => un4_sacqtime_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_19_c_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36247\,
            in2 => \N__38071\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_18,
            carryout => un4_sacqtime_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_20_c_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36147\,
            in2 => \N__38074\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_19,
            carryout => un4_sacqtime_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounter_RNIR3KA_0_20_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__36148\,
            in1 => \N__36065\,
            in2 => \N__38069\,
            in3 => \_gnd_net_\,
            lcout => op_gt_op_gt_un13_striginternallto23_8,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_20,
            carryout => un4_sacqtime_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_22_c_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38033\,
            in2 => \N__35980\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_21,
            carryout => un4_sacqtime_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_23_c_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38043\,
            in2 => \N__37083\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un4_sacqtime_cry_22,
            carryout => un4_sacqtime_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_23_THRU_LUT4_0_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25473\,
            lcout => \un4_sacqtime_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \button_debounce_counter_esr_RNO_0_23_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__32624\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26250\,
            lcout => \LED3_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_0_LC_10_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26826\,
            in1 => \N__25661\,
            in2 => \N__25605\,
            in3 => \N__25604\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_2_0_\,
            carryout => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0\,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53124\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_1_LC_10_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26828\,
            in1 => \N__25674\,
            in2 => \_gnd_net_\,
            in3 => \N__25461\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0\,
            carryout => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1\,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53124\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_2_LC_10_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26827\,
            in1 => \N__25620\,
            in2 => \_gnd_net_\,
            in3 => \N__25458\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1\,
            carryout => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2\,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53124\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_3_LC_10_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25647\,
            in2 => \_gnd_net_\,
            in3 => \N__25455\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2\,
            carryout => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3\,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53124\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_4_LC_10_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25686\,
            in2 => \_gnd_net_\,
            in3 => \N__25692\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3\,
            carryout => \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4\,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53124\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_5_LC_10_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25635\,
            in2 => \_gnd_net_\,
            in3 => \N__25689\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53124\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_RNICMDR1_0_LC_10_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__25685\,
            in1 => \N__25673\,
            in2 => \N__25662\,
            in3 => \N__25646\,
            lcout => OPEN,
            ltout => \spi_slave_inst.rx_data_count_neg_sclk_i6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_RNILK4P2_5_LC_10_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__25634\,
            in1 => \_gnd_net_\,
            in2 => \N__25623\,
            in3 => \N__25619\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_i6\,
            ltout => \spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3_5_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000111"
        )
    port map (
            in0 => \N__52419\,
            in1 => \N__38525\,
            in2 => \N__25608\,
            in3 => \N__33286\,
            lcout => \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_RNICH5T1_0_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__25589\,
            in1 => \N__25573\,
            in2 => \N__25556\,
            in3 => \N__25532\,
            lcout => \spi_slave_inst.un23_i_ssn_3\,
            ltout => \spi_slave_inst.un23_i_ssn_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_RNI5DOR2_5_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25795\,
            in2 => \N__25521\,
            in3 => \N__25773\,
            lcout => \spi_slave_inst.un23_i_ssn\,
            ltout => \spi_slave_inst.un23_i_ssn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_data_count_pos_sclk_i_RNI4ODL3_5_LC_10_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000111"
        )
    port map (
            in0 => \N__52420\,
            in1 => \N__38526\,
            in2 => \N__25506\,
            in3 => \N__33287\,
            lcout => \spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.spi_cs_i_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__38527\,
            in1 => \_gnd_net_\,
            in2 => \N__33291\,
            in3 => \N__52421\,
            lcout => \spi_slave_inst.spi_cs_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_done_pos_sclk_i_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__25803\,
            in1 => \N__25797\,
            in2 => \_gnd_net_\,
            in3 => \N__25778\,
            lcout => \spi_slave_inst.rx_done_pos_sclk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30704\,
            ce => \N__30664\,
            sr => \N__53095\
        );

    \spi_master_inst.spi_data_path_u1.data_in_6_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42252\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53247\,
            ce => \N__28842\,
            sr => \N__53082\
        );

    \spi_master_inst.spi_data_path_u1.data_in_1_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37623\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53247\,
            ce => \N__28842\,
            sr => \N__53082\
        );

    \spi_master_inst.spi_data_path_u1.data_in_2_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26841\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53247\,
            ce => \N__28842\,
            sr => \N__53082\
        );

    \spi_master_inst.spi_data_path_u1.data_in_11_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37605\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53247\,
            ce => \N__28842\,
            sr => \N__53082\
        );

    \spi_master_inst.spi_data_path_u1.data_in_12_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37587\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53247\,
            ce => \N__28842\,
            sr => \N__53082\
        );

    \spi_master_inst.spi_data_path_u1.data_in_3_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41370\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53247\,
            ce => \N__28842\,
            sr => \N__53082\
        );

    \spi_master_inst.spi_data_path_u1.data_in_14_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37719\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53247\,
            ce => \N__28842\,
            sr => \N__53082\
        );

    \spi_master_inst.spi_data_path_u1.data_in_15_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37701\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53247\,
            ce => \N__28842\,
            sr => \N__53082\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_0_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25864\,
            in1 => \N__25980\,
            in2 => \_gnd_net_\,
            in3 => \N__25968\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_6_0_\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0\,
            clk => \N__53251\,
            ce => \N__25818\,
            sr => \N__53070\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_1_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25859\,
            in1 => \N__25965\,
            in2 => \_gnd_net_\,
            in3 => \N__25950\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1\,
            clk => \N__53251\,
            ce => \N__25818\,
            sr => \N__53070\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_2_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25865\,
            in1 => \N__25946\,
            in2 => \_gnd_net_\,
            in3 => \N__25932\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2\,
            clk => \N__53251\,
            ce => \N__25818\,
            sr => \N__53070\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_3_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25860\,
            in1 => \N__25929\,
            in2 => \_gnd_net_\,
            in3 => \N__25917\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3\,
            clk => \N__53251\,
            ce => \N__25818\,
            sr => \N__53070\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_4_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25866\,
            in1 => \N__25914\,
            in2 => \_gnd_net_\,
            in3 => \N__25902\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4\,
            clk => \N__53251\,
            ce => \N__25818\,
            sr => \N__53070\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_5_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25861\,
            in1 => \N__25899\,
            in2 => \_gnd_net_\,
            in3 => \N__25887\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5\,
            clk => \N__53251\,
            ce => \N__25818\,
            sr => \N__53070\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_6_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25862\,
            in1 => \N__25883\,
            in2 => \_gnd_net_\,
            in3 => \N__25869\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6\,
            ltout => OPEN,
            carryin => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5\,
            carryout => \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6\,
            clk => \N__53251\,
            ce => \N__25818\,
            sr => \N__53070\
        );

    \spi_master_inst.sclk_gen_u0.clk_falling_count_i_7_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__25830\,
            in1 => \N__25863\,
            in2 => \_gnd_net_\,
            in3 => \N__25833\,
            lcout => \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53251\,
            ce => \N__25818\,
            sr => \N__53070\
        );

    \sEETrigCounter_0_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51041\,
            lcout => \sEETrigCounterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47814\,
            ce => \N__31016\,
            sr => \N__53059\
        );

    \sEETrigCounter_1_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50692\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEETrigCounterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47814\,
            ce => \N__31016\,
            sr => \N__53059\
        );

    \sEETrigCounter_2_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50123\,
            lcout => \sEETrigCounterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47814\,
            ce => \N__31016\,
            sr => \N__53059\
        );

    \sEETrigCounter_3_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49651\,
            lcout => \sEETrigCounterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47814\,
            ce => \N__31016\,
            sr => \N__53059\
        );

    \sEETrigCounter_RNII1HP1_2_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100001"
        )
    port map (
            in0 => \N__26081\,
            in1 => \N__26042\,
            in2 => \N__26121\,
            in3 => \N__26014\,
            lcout => un10_trig_prev_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIKN4B1_2_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000101"
        )
    port map (
            in0 => \N__26016\,
            in1 => \_gnd_net_\,
            in2 => \N__26043\,
            in3 => \N__26080\,
            lcout => un10_trig_prev_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNIR6CE_0_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26037\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un10_trig_prev_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigCounter_RNINEOS_1_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26038\,
            in2 => \_gnd_net_\,
            in3 => \N__26015\,
            lcout => un10_trig_prev_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_22_0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51138\,
            lcout => \sDAC_mem_22Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47791\,
            ce => \N__39817\,
            sr => \N__53039\
        );

    \sDAC_mem_22_7_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48706\,
            lcout => \sDAC_mem_22Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47791\,
            ce => \N__39817\,
            sr => \N__53039\
        );

    \spi_slave_inst.rx_done_reg3_i_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28793\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_inst.rx_done_reg3_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47777\,
            ce => 'H',
            sr => \N__53029\
        );

    \spi_slave_inst.rx_ready_i_RNO_0_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26133\,
            in2 => \_gnd_net_\,
            in3 => \N__28792\,
            lcout => OPEN,
            ltout => \spi_slave_inst.rx_ready_i_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rx_ready_i_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__32466\,
            in1 => \N__33230\,
            in2 => \N__26127\,
            in3 => \N__27314\,
            lcout => spi_mosi_ready,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47777\,
            ce => 'H',
            sr => \N__53029\
        );

    \spi_mosi_ready_prev_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27315\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_mosi_ready_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47777\,
            ce => 'H',
            sr => \N__53029\
        );

    \spi_mosi_ready_prev2_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26208\,
            lcout => \spi_mosi_ready_prevZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47777\,
            ce => 'H',
            sr => \N__53029\
        );

    \spi_slave_inst.tx_ready_i_RNO_0_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27090\,
            in2 => \_gnd_net_\,
            in3 => \N__27105\,
            lcout => OPEN,
            ltout => \spi_slave_inst.un4_tx_done_reg2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_ready_i_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__32467\,
            in1 => \N__33231\,
            in2 => \N__26124\,
            in3 => \N__26183\,
            lcout => \spi_slave_inst.tx_ready_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47777\,
            ce => 'H',
            sr => \N__53029\
        );

    \spi_mosi_ready_prev3_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26220\,
            lcout => \spi_mosi_ready_prevZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47777\,
            ce => 'H',
            sr => \N__53029\
        );

    \button_debounce_counter_0_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__32468\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26298\,
            lcout => \button_debounce_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53262\,
            ce => 'H',
            sr => \N__26239\
        );

    \button_debounce_counter_1_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__26299\,
            in1 => \N__32469\,
            in2 => \_gnd_net_\,
            in3 => \N__26267\,
            lcout => \button_debounce_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53262\,
            ce => 'H',
            sr => \N__26239\
        );

    \spi_mosi_ready_prev3_RNILKER_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__26219\,
            in1 => \N__26207\,
            in2 => \N__26196\,
            in3 => \N__27313\,
            lcout => \spi_mosi_ready_prev3_RNILKERZ0\,
            ltout => \spi_mosi_ready_prev3_RNILKERZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_rpi_ibuf_RNI7JCV_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__32470\,
            in1 => \_gnd_net_\,
            in2 => \N__26187\,
            in3 => \_gnd_net_\,
            lcout => \reset_rpi_ibuf_RNI7JCVZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_0_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__31094\,
            in1 => \N__40395\,
            in2 => \N__27141\,
            in3 => \N__44749\,
            lcout => \sAddress_RNIA6242Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_ready_i_RNIBLID_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32398\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26184\,
            lcout => \spi_slave_inst.un4_i_wr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sRead_data_RNO_0_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27978\,
            in2 => \_gnd_net_\,
            in3 => \N__27882\,
            lcout => \N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sADC_clk_prev_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27621\,
            lcout => \sADC_clk_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47792\,
            ce => \N__26754\,
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_0_c_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34154\,
            in2 => \N__26168\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => un1_sacqtime_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_1_c_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35075\,
            in2 => \N__26150\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_0,
            carryout => un1_sacqtime_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_2_c_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34877\,
            in2 => \N__26459\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_1,
            carryout => un1_sacqtime_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_3_c_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34772\,
            in2 => \N__26441\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_2,
            carryout => un1_sacqtime_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_4_c_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34745\,
            in2 => \N__26423\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_3,
            carryout => un1_sacqtime_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_5_c_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34640\,
            in2 => \N__26405\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_4,
            carryout => un1_sacqtime_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_6_c_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34514\,
            in2 => \N__26387\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_5,
            carryout => un1_sacqtime_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_7_c_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34397\,
            in2 => \N__26366\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_6,
            carryout => un1_sacqtime_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_8_c_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35792\,
            in2 => \N__26348\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => un1_sacqtime_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_9_c_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35681\,
            in2 => \N__26330\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_8,
            carryout => un1_sacqtime_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_10_c_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35567\,
            in2 => \N__26582\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_9,
            carryout => un1_sacqtime_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_11_c_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35462\,
            in2 => \N__26564\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_10,
            carryout => un1_sacqtime_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_12_c_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35435\,
            in2 => \N__26546\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_11,
            carryout => un1_sacqtime_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_13_c_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35231\,
            in2 => \N__26528\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_12,
            carryout => un1_sacqtime_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_14_c_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35111\,
            in2 => \N__26510\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_13,
            carryout => un1_sacqtime_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_15_c_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36569\,
            in2 => \N__26493\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_14,
            carryout => un1_sacqtime_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_16_c_inv_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36517\,
            in1 => \_gnd_net_\,
            in2 => \N__26478\,
            in3 => \_gnd_net_\,
            lcout => un1_sacqtime_cry_16_sf,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => un1_sacqtime_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_17_c_inv_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36416\,
            in1 => \_gnd_net_\,
            in2 => \N__26469\,
            in3 => \_gnd_net_\,
            lcout => un1_sacqtime_cry_17_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_16,
            carryout => un1_sacqtime_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_18_c_inv_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26703\,
            in3 => \N__36323\,
            lcout => un1_sacqtime_cry_18_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_17,
            carryout => un1_sacqtime_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_19_c_inv_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26694\,
            in3 => \N__36231\,
            lcout => un1_sacqtime_cry_19_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_18,
            carryout => un1_sacqtime_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_20_c_inv_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26685\,
            in3 => \N__36146\,
            lcout => un1_sacqtime_cry_20_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_19,
            carryout => un1_sacqtime_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_21_c_inv_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36063\,
            in1 => \_gnd_net_\,
            in2 => \N__26676\,
            in3 => \_gnd_net_\,
            lcout => un1_sacqtime_cry_21_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_20,
            carryout => un1_sacqtime_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_22_c_inv_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26667\,
            in3 => \N__35960\,
            lcout => un1_sacqtime_cry_22_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_21,
            carryout => un1_sacqtime_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_23_c_inv_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__37058\,
            in1 => \_gnd_net_\,
            in2 => \N__26658\,
            in3 => \_gnd_net_\,
            lcout => un1_sacqtime_cry_23_sf,
            ltout => OPEN,
            carryin => un1_sacqtime_cry_22,
            carryout => un1_sacqtime_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_sacqtime_cry_23_THRU_LUT4_0_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26649\,
            lcout => \un1_sacqtime_cry_23_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_10_RNO_0_15_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__26627\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31670\,
            lcout => \N_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPointerReset_RNI2CQM_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__33475\,
            in1 => \N__31669\,
            in2 => \N__32178\,
            in3 => \N__31847\,
            lcout => \N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sADC_clk_prev_RNO_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__31848\,
            in1 => \N__32102\,
            in2 => \_gnd_net_\,
            in3 => \N__32413\,
            lcout => \N_76_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sADC_clk_prev_RNI4BVG_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__27636\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27606\,
            lcout => \N_71\,
            ltout => \N_71_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_15_RNO_0_15_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26742\,
            in3 => \N__28352\,
            lcout => \N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEDelayACQ_0_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51266\,
            lcout => \sEEDelayACQZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__27219\,
            sr => \N__52979\
        );

    \sEEDelayACQ_1_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50769\,
            lcout => \sEEDelayACQZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__27219\,
            sr => \N__52979\
        );

    \sEEDelayACQ_2_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50305\,
            lcout => \sEEDelayACQZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__27219\,
            sr => \N__52979\
        );

    \sEEDelayACQ_3_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49834\,
            lcout => \sEEDelayACQZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__27219\,
            sr => \N__52979\
        );

    \sEEDelayACQ_4_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49306\,
            lcout => \sEEDelayACQZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__27219\,
            sr => \N__52979\
        );

    \sEEDelayACQ_5_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47130\,
            lcout => \sEEDelayACQZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__27219\,
            sr => \N__52979\
        );

    \sEEDelayACQ_6_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48230\,
            lcout => \sEEDelayACQZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__27219\,
            sr => \N__52979\
        );

    \sEEDelayACQ_7_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48832\,
            lcout => \sEEDelayACQZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47839\,
            ce => \N__27219\,
            sr => \N__52979\
        );

    \sEEDelayACQ_10_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50306\,
            lcout => \sEEDelayACQZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => \N__26946\,
            sr => \N__52975\
        );

    \sEEDelayACQ_11_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49790\,
            lcout => \sEEDelayACQZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => \N__26946\,
            sr => \N__52975\
        );

    \sEEDelayACQ_12_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49189\,
            lcout => \sEEDelayACQZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => \N__26946\,
            sr => \N__52975\
        );

    \sEEDelayACQ_13_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47149\,
            lcout => \sEEDelayACQZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => \N__26946\,
            sr => \N__52975\
        );

    \sEEDelayACQ_14_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48231\,
            lcout => \sEEDelayACQZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => \N__26946\,
            sr => \N__52975\
        );

    \sEEDelayACQ_15_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48768\,
            lcout => \sEEDelayACQZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => \N__26946\,
            sr => \N__52975\
        );

    \sEEDelayACQ_8_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51267\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => \N__26946\,
            sr => \N__52975\
        );

    \sEEDelayACQ_9_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50770\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEDelayACQZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47847\,
            ce => \N__26946\,
            sr => \N__52975\
        );

    \RAM_DATA_cl_12_RNO_0_15_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26912\,
            in2 => \_gnd_net_\,
            in3 => \N__31708\,
            lcout => OPEN,
            ltout => \N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_12_15_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32502\,
            in1 => \N__32067\,
            in2 => \N__26934\,
            in3 => \N__31968\,
            lcout => \RAM_DATA_cl_12Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47851\,
            ce => 'H',
            sr => \N__52971\
        );

    \RAM_DATA_cl_11_RNO_0_15_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26879\,
            in2 => \_gnd_net_\,
            in3 => \N__31707\,
            lcout => OPEN,
            ltout => \N_94_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_11_15_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32501\,
            in1 => \N__32066\,
            in2 => \N__26901\,
            in3 => \N__31967\,
            lcout => \RAM_DATA_cl_11Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47851\,
            ce => 'H',
            sr => \N__52971\
        );

    \RAM_DATA_cl_14_RNO_0_15_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26852\,
            in2 => \_gnd_net_\,
            in3 => \N__31709\,
            lcout => OPEN,
            ltout => \N_104_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_14_15_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32503\,
            in1 => \N__32068\,
            in2 => \N__26868\,
            in3 => \N__31969\,
            lcout => \RAM_DATA_cl_14Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47851\,
            ce => 'H',
            sr => \N__52971\
        );

    \sDAC_data_2_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53243\,
            ce => \N__42234\,
            sr => \N__53109\
        );

    \spi_slave_inst.rx_done_neg_sclk_i_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__27065\,
            in1 => \N__33194\,
            in2 => \_gnd_net_\,
            in3 => \N__26829\,
            lcout => \spi_slave_inst.rx_done_neg_sclk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi_slave_inst.rx_done_neg_sclk_iC_net\,
            ce => 'H',
            sr => \N__53096\
        );

    \spi_slave_inst.rx_done_reg1_i_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27066\,
            in1 => \N__33214\,
            in2 => \_gnd_net_\,
            in3 => \N__27054\,
            lcout => \spi_slave_inst.rx_done_reg1_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47832\,
            ce => 'H',
            sr => \N__53083\
        );

    \spi_slave_inst.txdata_reg_i_5_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27378\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47832\,
            ce => 'H',
            sr => \N__53083\
        );

    \spi_slave_inst.txdata_reg_i_4_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27237\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47832\,
            ce => 'H',
            sr => \N__53083\
        );

    \spi_master_inst.spi_data_path_u1.tx_ready_i_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011110100"
        )
    port map (
            in0 => \N__27048\,
            in1 => \N__27041\,
            in2 => \N__28837\,
            in3 => \N__47306\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_ready_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53245\,
            ce => 'H',
            sr => \N__53071\
        );

    \spi_master_inst.spi_data_path_u1.tx_done_reg3_i_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27042\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53245\,
            ce => 'H',
            sr => \N__53071\
        );

    \spi_master_inst.spi_data_path_u1.tx_done_reg2_i_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27009\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53245\,
            ce => 'H',
            sr => \N__53071\
        );

    \spi_master_inst.spi_data_path_u1.tx_done_reg1_i_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27033\,
            lcout => \spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53245\,
            ce => 'H',
            sr => \N__53071\
        );

    \spi_master_inst.sclk_gen_u0.spi_start_i_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47307\,
            lcout => \spi_master_inst.sclk_gen_u0.spi_start_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53245\,
            ce => 'H',
            sr => \N__53071\
        );

    \spi_slave_inst.txdata_reg_i_RNI1IQC_0_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37153\,
            in1 => \N__26958\,
            in2 => \_gnd_net_\,
            in3 => \N__27078\,
            lcout => \spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.txdata_reg_i_RNI7OQC_3_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27204\,
            in1 => \N__27195\,
            in2 => \_gnd_net_\,
            in3 => \N__37162\,
            lcout => OPEN,
            ltout => \spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNIUCSS_1_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__27177\,
            in1 => \_gnd_net_\,
            in2 => \N__27129\,
            in3 => \N__37221\,
            lcout => \spi_slave_inst.N_1394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ8SS_1_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27162\,
            in1 => \N__27126\,
            in2 => \_gnd_net_\,
            in3 => \N__37220\,
            lcout => OPEN,
            ltout => \spi_slave_inst.N_1397_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNIA0LM2_0_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__33224\,
            in1 => \N__27120\,
            in2 => \N__27114\,
            in3 => \N__37251\,
            lcout => \spi_slave_inst.spi_miso\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_23_7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48599\,
            lcout => \sDAC_mem_23Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47804\,
            ce => \N__28989\,
            sr => \N__53049\
        );

    \sPointer_1_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011001000100"
        )
    port map (
            in0 => \N__29217\,
            in1 => \N__43832\,
            in2 => \_gnd_net_\,
            in3 => \N__29189\,
            lcout => \sPointerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47793\,
            ce => 'H',
            sr => \N__53040\
        );

    \spi_slave_inst.tx_done_reg1_i_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33159\,
            lcout => \spi_slave_inst.tx_done_reg1_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47793\,
            ce => 'H',
            sr => \N__53040\
        );

    \spi_slave_inst.tx_done_reg2_i_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27111\,
            lcout => \spi_slave_inst.tx_done_reg2_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47793\,
            ce => 'H',
            sr => \N__53040\
        );

    \spi_slave_inst.tx_done_reg3_i_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27104\,
            lcout => \spi_slave_inst.tx_done_reg3_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47793\,
            ce => 'H',
            sr => \N__53040\
        );

    \spi_slave_inst.txdata_reg_i_0_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27273\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47793\,
            ce => 'H',
            sr => \N__53040\
        );

    \spi_slave_inst.txdata_reg_i_3_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27246\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47793\,
            ce => 'H',
            sr => \N__53040\
        );

    \spi_slave_inst.txdata_reg_i_7_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27357\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47793\,
            ce => 'H',
            sr => \N__53040\
        );

    \spi_slave_inst.txdata_reg_i_RNI3KQC_1_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27168\,
            in1 => \N__27186\,
            in2 => \_gnd_net_\,
            in3 => \N__37163\,
            lcout => \spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.txdata_reg_i_1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27264\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47778\,
            ce => 'H',
            sr => \N__53030\
        );

    \spi_slave_inst.txdata_reg_i_RNI5MQC_2_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37164\,
            in1 => \N__27147\,
            in2 => \_gnd_net_\,
            in3 => \N__27153\,
            lcout => \spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.txdata_reg_i_2_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27255\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47778\,
            ce => 'H',
            sr => \N__53030\
        );

    \spi_slave_inst.txdata_reg_i_6_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27366\,
            lcout => \spi_slave_inst.txdata_reg_iZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47778\,
            ce => 'H',
            sr => \N__53030\
        );

    \sPointer_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000110101010"
        )
    port map (
            in0 => \N__29188\,
            in1 => \N__43833\,
            in2 => \_gnd_net_\,
            in3 => \N__29213\,
            lcout => \sPointerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47778\,
            ce => 'H',
            sr => \N__53030\
        );

    \sAddress_RNIAM2A_0_1_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000010"
        )
    port map (
            in0 => \N__44952\,
            in1 => \N__40326\,
            in2 => \N__40538\,
            in3 => \N__44869\,
            lcout => \N_206\,
            ltout => \N_206_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_1_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40327\,
            in1 => \N__31072\,
            in2 => \N__27222\,
            in3 => \N__44718\,
            lcout => \sAddress_RNIA6242_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIQ63A_6_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__30946\,
            in1 => \N__46485\,
            in2 => \N__30926\,
            in3 => \N__44613\,
            lcout => \N_141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_4_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49230\,
            in2 => \_gnd_net_\,
            in3 => \N__43843\,
            lcout => \sAddressZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47764\,
            ce => \N__43775\,
            sr => \N__53020\
        );

    \sAddress_6_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__43844\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48159\,
            lcout => \sAddressZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47764\,
            ce => \N__43775\,
            sr => \N__53020\
        );

    \sAddress_RNIFL15_6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30922\,
            in2 => \_gnd_net_\,
            in3 => \N__30947\,
            lcout => \sDAC_mem_30_1_sqmuxa_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_7_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__43845\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48592\,
            lcout => \sAddressZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47764\,
            ce => \N__43775\,
            sr => \N__53020\
        );

    \sEEPointerReset_RNO_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__43846\,
            in1 => \N__29191\,
            in2 => \N__32554\,
            in3 => \N__29128\,
            lcout => \N_269\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sPointer_RNIPU81_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29190\,
            in2 => \_gnd_net_\,
            in3 => \N__43847\,
            lcout => \N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_mosi_ready64_prev_e_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27312\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_mosi_ready64_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47754\,
            ce => \N__32515\,
            sr => \_gnd_net_\
        );

    \spi_mosi_ready64_prev3_e_0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27342\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_mosi_ready64_prevZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47754\,
            ce => \N__32515\,
            sr => \_gnd_net_\
        );

    \spi_mosi_ready64_prev2_e_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27333\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_mosi_ready64_prevZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47754\,
            ce => \N__32515\,
            sr => \_gnd_net_\
        );

    \spi_mosi_ready64_prev3_e_0_RNICM2C1_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27341\,
            in1 => \N__27332\,
            in2 => \N__27324\,
            in3 => \N__27311\,
            lcout => \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1\,
            ltout => \spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sPointer_RNI85NC1_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27291\,
            in3 => \N__29192\,
            lcout => un1_spointer11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_rpi_ibuf_RNIIUT3_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32516\,
            lcout => \LED3_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.data_in_reg_i_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29526\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47765\,
            ce => \N__27348\,
            sr => \N__53009\
        );

    \spi_slave_inst.data_in_reg_i_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29481\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47765\,
            ce => \N__27348\,
            sr => \N__53009\
        );

    \spi_slave_inst.data_in_reg_i_2_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29421\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47765\,
            ce => \N__27348\,
            sr => \N__53009\
        );

    \spi_slave_inst.data_in_reg_i_3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30009\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47765\,
            ce => \N__27348\,
            sr => \N__53009\
        );

    \spi_slave_inst.data_in_reg_i_4_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29952\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47765\,
            ce => \N__27348\,
            sr => \N__53009\
        );

    \spi_slave_inst.data_in_reg_i_5_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29799\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47765\,
            ce => \N__27348\,
            sr => \N__53009\
        );

    \spi_slave_inst.data_in_reg_i_6_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27720\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47765\,
            ce => \N__27348\,
            sr => \N__53009\
        );

    \spi_slave_inst.data_in_reg_i_7_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27669\,
            lcout => \spi_slave_inst.data_in_reg_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47765\,
            ce => \N__27348\,
            sr => \N__53009\
        );

    \sEEACQ_0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51080\,
            lcout => \sEEACQZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47779\,
            ce => \N__28911\,
            sr => \N__53001\
        );

    \sEEACQ_1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50664\,
            lcout => \sEEACQZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47779\,
            ce => \N__28911\,
            sr => \N__53001\
        );

    \sEEACQ_2_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50274\,
            lcout => \sEEACQZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47779\,
            ce => \N__28911\,
            sr => \N__53001\
        );

    \sEEACQ_3_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49689\,
            lcout => \sEEACQZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47779\,
            ce => \N__28911\,
            sr => \N__53001\
        );

    \sEEACQ_4_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49368\,
            lcout => \sEEACQZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47779\,
            ce => \N__28911\,
            sr => \N__53001\
        );

    \sEEACQ_5_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47046\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEACQZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47779\,
            ce => \N__28911\,
            sr => \N__53001\
        );

    \sEEACQ_6_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48274\,
            lcout => \sEEACQZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47779\,
            ce => \N__28911\,
            sr => \N__53001\
        );

    \sEEACQ_7_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48705\,
            lcout => \sEEACQZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47779\,
            ce => \N__28911\,
            sr => \N__53001\
        );

    \spi_data_miso_6_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__27765\,
            in1 => \N__29852\,
            in2 => \N__27741\,
            in3 => \N__29937\,
            lcout => \spi_data_misoZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47794\,
            ce => \N__29780\,
            sr => \N__52992\
        );

    \spi_data_miso_7_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111111101010"
        )
    port map (
            in0 => \N__29938\,
            in1 => \N__27711\,
            in2 => \N__29868\,
            in3 => \N__27687\,
            lcout => \spi_data_misoZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47794\,
            ce => \N__29780\,
            sr => \N__52992\
        );

    \RAM_nWE_obuf_RNO_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__27617\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29939\,
            lcout => \RAM_nWE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sADC_clk_prev_RNIM9TK_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__32351\,
            in1 => \N__27635\,
            in2 => \_gnd_net_\,
            in3 => \N__27616\,
            lcout => \sRAM_ADD_0_sqmuxa_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_rpi_ibuf_RNI4GQD1_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__32350\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27575\,
            lcout => \N_1470_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sRead_data_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000100"
        )
    port map (
            in0 => \N__29933\,
            in1 => \N__29851\,
            in2 => \N__27486\,
            in3 => \N__27470\,
            lcout => \sRead_dataZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47805\,
            ce => 'H',
            sr => \N__52987\
        );

    \sCounterRAM_RNISREI1_7_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27456\,
            in1 => \N__27438\,
            in2 => \N__27417\,
            in3 => \N__27396\,
            lcout => OPEN,
            ltout => \spi_data_miso_0_sqmuxa_2_i_o2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterRAM_RNIS8L63_1_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28038\,
            in1 => \N__28020\,
            in2 => \N__27999\,
            in3 => \N__27996\,
            lcout => \N_75\,
            ltout => \N_75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_23_c_RNIGRPG4_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110101111"
        )
    port map (
            in0 => \N__27858\,
            in1 => \N__32217\,
            in2 => \N__27984\,
            in3 => \N__31916\,
            lcout => \N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sSPI_MSB0LSB1_RNINK761_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27979\,
            in2 => \_gnd_net_\,
            in3 => \N__27897\,
            lcout => \N_88\,
            ltout => \N_88_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPointerReset_RNILL2C1_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101011111010"
        )
    port map (
            in0 => \N__33434\,
            in1 => \N__31915\,
            in2 => \N__27852\,
            in3 => \N__32216\,
            lcout => \N_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_9_RNO_0_15_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__31684\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27806\,
            lcout => OPEN,
            ltout => \N_93_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_9_15_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__31885\,
            in1 => \N__32214\,
            in2 => \N__27825\,
            in3 => \N__32354\,
            lcout => \RAM_DATA_cl_9Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47815\,
            ce => 'H',
            sr => \N__52982\
        );

    \RAM_DATA_cl_RNO_0_15_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__31685\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27776\,
            lcout => OPEN,
            ltout => \N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_15_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__31883\,
            in1 => \N__32212\,
            in2 => \N__27795\,
            in3 => \N__32352\,
            lcout => \RAM_DATA_clZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47815\,
            ce => 'H',
            sr => \N__52982\
        );

    \RAM_DATA_cl_8_RNO_0_15_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__31683\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28310\,
            lcout => OPEN,
            ltout => \N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_8_15_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__31884\,
            in1 => \N__32213\,
            in2 => \N__28329\,
            in3 => \N__32353\,
            lcout => \RAM_DATA_cl_8Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47815\,
            ce => 'H',
            sr => \N__52982\
        );

    \un4_sacqtime_cry_23_c_RNITTS3_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32211\,
            in2 => \_gnd_net_\,
            in3 => \N__31882\,
            lcout => \un4_sacqtime_cry_23_c_RNITTSZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sRAM_ADD_14_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__33015\,
            in1 => \N__32196\,
            in2 => \N__28299\,
            in3 => \N__31960\,
            lcout => \RAM_ADD_c_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47823\,
            ce => \N__30267\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_15_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__31957\,
            in1 => \N__32994\,
            in2 => \N__32226\,
            in3 => \N__28248\,
            lcout => \RAM_ADD_c_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47823\,
            ce => \N__30267\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_16_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__28209\,
            in1 => \N__32973\,
            in2 => \N__32221\,
            in3 => \N__31961\,
            lcout => \RAM_ADD_c_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47823\,
            ce => \N__30267\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_17_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__31958\,
            in1 => \N__28164\,
            in2 => \N__32227\,
            in3 => \N__32952\,
            lcout => \RAM_ADD_c_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47823\,
            ce => \N__30267\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_18_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__33327\,
            in1 => \N__32197\,
            in2 => \N__28125\,
            in3 => \N__31962\,
            lcout => \RAM_ADD_c_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47823\,
            ce => \N__30267\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_2_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__31959\,
            in1 => \N__28080\,
            in2 => \N__32228\,
            in3 => \N__32925\,
            lcout => \RAM_ADD_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47823\,
            ce => \N__30267\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_3_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__31956\,
            in1 => \N__32198\,
            in2 => \N__28689\,
            in3 => \N__32904\,
            lcout => \RAM_ADD_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47823\,
            ce => \N__30267\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_4_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__32883\,
            in1 => \N__31955\,
            in2 => \N__32229\,
            in3 => \N__28650\,
            lcout => \RAM_ADD_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47823\,
            ce => \N__30267\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_5_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__28605\,
            in1 => \N__32163\,
            in2 => \N__32859\,
            in3 => \N__31912\,
            lcout => \RAM_ADD_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => \N__30263\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_6_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__31910\,
            in1 => \N__28560\,
            in2 => \N__32219\,
            in3 => \N__32838\,
            lcout => \RAM_ADD_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => \N__30263\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_7_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__32820\,
            in1 => \N__32164\,
            in2 => \N__28512\,
            in3 => \N__31913\,
            lcout => \RAM_ADD_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => \N__30263\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_8_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__31911\,
            in1 => \N__28464\,
            in2 => \N__32220\,
            in3 => \N__32802\,
            lcout => \RAM_ADD_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => \N__30263\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_9_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__32781\,
            in1 => \N__32165\,
            in2 => \N__28419\,
            in3 => \N__31914\,
            lcout => \RAM_ADD_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47833\,
            ce => \N__30263\,
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_15_15_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__31963\,
            in1 => \N__32444\,
            in2 => \N__32218\,
            in3 => \N__28371\,
            lcout => \RAM_DATA_cl_15Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47840\,
            ce => 'H',
            sr => \N__52972\
        );

    \RAM_DATA_cl_13_15_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__30492\,
            in1 => \N__32159\,
            in2 => \N__32504\,
            in3 => \N__31964\,
            lcout => \RAM_DATA_cl_13Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47840\,
            ce => 'H',
            sr => \N__52972\
        );

    \RAM_DATA_cl_1_15_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__30528\,
            in1 => \N__32151\,
            in2 => \N__32505\,
            in3 => \N__31965\,
            lcout => \RAM_DATA_cl_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47848\,
            ce => 'H',
            sr => \N__52968\
        );

    \RAM_DATA_cl_2_15_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__30459\,
            in1 => \N__32152\,
            in2 => \N__32506\,
            in3 => \N__31966\,
            lcout => \RAM_DATA_cl_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47848\,
            ce => 'H',
            sr => \N__52968\
        );

    \spi_slave_inst.spi_cs_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__33285\,
            in1 => \N__38564\,
            in2 => \_gnd_net_\,
            in3 => \N__52425\,
            lcout => \spi_slave_inst.spi_csZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.spi_sclk_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28719\,
            in1 => \N__38565\,
            in2 => \_gnd_net_\,
            in3 => \N__52343\,
            lcout => spi_sclk,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_0_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53241\,
            ce => \N__42233\,
            sr => \N__53090\
        );

    \spi_slave_inst.rxdata_reg_i_0_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30795\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => spi_data_mosi_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => \N__28767\,
            sr => \N__53079\
        );

    \spi_slave_inst.rxdata_reg_i_1_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30783\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => spi_data_mosi_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => \N__28767\,
            sr => \N__53079\
        );

    \spi_slave_inst.rxdata_reg_i_2_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30771\,
            lcout => spi_data_mosi_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => \N__28767\,
            sr => \N__53079\
        );

    \spi_slave_inst.rxdata_reg_i_3_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30759\,
            lcout => spi_data_mosi_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => \N__28767\,
            sr => \N__53079\
        );

    \spi_slave_inst.rxdata_reg_i_4_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30747\,
            lcout => spi_data_mosi_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => \N__28767\,
            sr => \N__53079\
        );

    \spi_slave_inst.rxdata_reg_i_5_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30735\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => spi_data_mosi_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => \N__28767\,
            sr => \N__53079\
        );

    \spi_slave_inst.rxdata_reg_i_6_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30723\,
            lcout => spi_data_mosi_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => \N__28767\,
            sr => \N__53079\
        );

    \spi_slave_inst.rxdata_reg_i_7_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30711\,
            lcout => spi_data_mosi_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47834\,
            ce => \N__28767\,
            sr => \N__53079\
        );

    \spi_slave_inst.rx_done_reg1_i_RNID541_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28805\,
            in2 => \_gnd_net_\,
            in3 => \N__28794\,
            lcout => \spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rxdata_reg_i_RNINNBS_2_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__48910\,
            in1 => \N__49415\,
            in2 => \N__47948\,
            in3 => \N__49906\,
            lcout => \spi_slave_inst.un1_spointer11_2_0_a2_0_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_master_inst.spi_data_path_u1.data_in_10_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39468\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53244\,
            ce => \N__28841\,
            sr => \N__53057\
        );

    \spi_master_inst.spi_data_path_u1.data_in_13_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37731\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53244\,
            ce => \N__28841\,
            sr => \N__53057\
        );

    \spi_master_inst.spi_data_path_u1.data_in_4_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41202\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53244\,
            ce => \N__28841\,
            sr => \N__53057\
        );

    \spi_master_inst.spi_data_path_u1.data_in_5_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33768\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53244\,
            ce => \N__28841\,
            sr => \N__53057\
        );

    \spi_master_inst.spi_data_path_u1.data_in_0_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28899\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53244\,
            ce => \N__28841\,
            sr => \N__53057\
        );

    \spi_master_inst.spi_data_path_u1.data_in_7_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37425\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53244\,
            ce => \N__28841\,
            sr => \N__53057\
        );

    \spi_master_inst.spi_data_path_u1.data_in_8_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40917\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53244\,
            ce => \N__28841\,
            sr => \N__53057\
        );

    \spi_master_inst.spi_data_path_u1.data_in_9_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39171\,
            lcout => \spi_master_inst.spi_data_path_u1.data_inZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53244\,
            ce => \N__28841\,
            sr => \N__53057\
        );

    \sDAC_mem_4_1_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50454\,
            lcout => \sDAC_mem_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47806\,
            ce => \N__39635\,
            sr => \N__53047\
        );

    \sDAC_mem_4_4_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48988\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47806\,
            ce => \N__39635\,
            sr => \N__53047\
        );

    \sDAC_mem_23_0_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50881\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_23Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47795\,
            ce => \N__28988\,
            sr => \N__53038\
        );

    \sDAC_mem_23_1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50455\,
            lcout => \sDAC_mem_23Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47795\,
            ce => \N__28988\,
            sr => \N__53038\
        );

    \sDAC_mem_23_2_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50023\,
            lcout => \sDAC_mem_23Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47795\,
            ce => \N__28988\,
            sr => \N__53038\
        );

    \sDAC_mem_23_3_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49572\,
            lcout => \sDAC_mem_23Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47795\,
            ce => \N__28988\,
            sr => \N__53038\
        );

    \sDAC_mem_23_4_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49076\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_23Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47795\,
            ce => \N__28988\,
            sr => \N__53038\
        );

    \sDAC_mem_23_5_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46861\,
            lcout => \sDAC_mem_23Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47795\,
            ce => \N__28988\,
            sr => \N__53038\
        );

    \sDAC_mem_23_6_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48160\,
            lcout => \sDAC_mem_23Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47795\,
            ce => \N__28988\,
            sr => \N__53038\
        );

    \sDAC_mem_33_0_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51025\,
            lcout => \sDAC_mem_33Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47780\,
            ce => \N__30858\,
            sr => \N__53027\
        );

    \sDAC_mem_33_1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50456\,
            lcout => \sDAC_mem_33Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47780\,
            ce => \N__30858\,
            sr => \N__53027\
        );

    \sDAC_mem_33_2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50024\,
            lcout => \sDAC_mem_33Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47780\,
            ce => \N__30858\,
            sr => \N__53027\
        );

    \sDAC_mem_33_3_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49573\,
            lcout => \sDAC_mem_33Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47780\,
            ce => \N__30858\,
            sr => \N__53027\
        );

    \sDAC_mem_33_4_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49131\,
            lcout => \sDAC_mem_33Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47780\,
            ce => \N__30858\,
            sr => \N__53027\
        );

    \sDAC_mem_33_5_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46958\,
            lcout => \sDAC_mem_33Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47780\,
            ce => \N__30858\,
            sr => \N__53027\
        );

    \sDAC_mem_33_6_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48161\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_33Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47780\,
            ce => \N__30858\,
            sr => \N__53027\
        );

    \sDAC_mem_33_7_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48597\,
            lcout => \sDAC_mem_33Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47780\,
            ce => \N__30858\,
            sr => \N__53027\
        );

    \sDAC_mem_1_0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51026\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47766\,
            ce => \N__42031\,
            sr => \N__53019\
        );

    \sDAC_mem_1_1_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50457\,
            lcout => \sDAC_mem_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47766\,
            ce => \N__42031\,
            sr => \N__53019\
        );

    \sDAC_mem_1_2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50025\,
            lcout => \sDAC_mem_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47766\,
            ce => \N__42031\,
            sr => \N__53019\
        );

    \sDAC_mem_1_7_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48598\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47766\,
            ce => \N__42031\,
            sr => \N__53019\
        );

    \sAddress_RNI25GS1_1_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__44871\,
            in1 => \N__31071\,
            in2 => \N__40355\,
            in3 => \N__44723\,
            lcout => un1_spointer11_5_0_2,
            ltout => \un1_spointer11_5_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_0_2_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__40518\,
            in1 => \N__44953\,
            in2 => \N__28914\,
            in3 => \N__40325\,
            lcout => \sAddress_RNIA6242_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_1_2_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__40323\,
            in1 => \N__40516\,
            in2 => \N__44961\,
            in3 => \N__30991\,
            lcout => \sAddress_RNIA6242_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_6_1_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__43142\,
            in1 => \N__44553\,
            in2 => \_gnd_net_\,
            in3 => \N__44444\,
            lcout => \sDAC_mem_32_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_16_3_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40324\,
            in1 => \N__40517\,
            in2 => \N__44571\,
            in3 => \N__43141\,
            lcout => \sDAC_mem_23_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sPointer_RNI5LBD1_0_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__29176\,
            in1 => \N__43856\,
            in2 => \_gnd_net_\,
            in3 => \N__29127\,
            lcout => \N_275\,
            ltout => \N_275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_rpi_ibuf_RNIHQCR1_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32558\,
            in2 => \N__28971\,
            in3 => \N__31070\,
            lcout => \N_360\,
            ltout => \N_360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEPointerReset_RNO_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__44549\,
            in1 => \N__44443\,
            in2 => \N__28968\,
            in3 => \N__28965\,
            lcout => \N_132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_0_0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40329\,
            in1 => \N__31073\,
            in2 => \N__28935\,
            in3 => \N__44716\,
            lcout => \sAddress_RNIA6242_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIAM2A_1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001010000"
        )
    port map (
            in0 => \N__44959\,
            in1 => \N__40328\,
            in2 => \N__40539\,
            in3 => \N__44870\,
            lcout => un1_spointer11_7_0_tz,
            ltout => \un1_spointer11_7_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNID9242_3_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40519\,
            in1 => \N__31074\,
            in2 => \N__28926\,
            in3 => \N__44717\,
            lcout => \sAddress_RNID9242Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_0_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__50873\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43860\,
            lcout => \sAddressZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47741\,
            ce => \N__43771\,
            sr => \N__53006\
        );

    \sAddress_3_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__43861\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49571\,
            lcout => \sAddressZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47741\,
            ce => \N__43771\,
            sr => \N__53006\
        );

    \sAddress_5_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46957\,
            in2 => \_gnd_net_\,
            in3 => \N__43862\,
            lcout => \sAddressZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47741\,
            ce => \N__43771\,
            sr => \N__53006\
        );

    \spi_slave_inst.rxdata_reg_i_RNILLBS_1_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__46956\,
            in1 => \N__50560\,
            in2 => \N__48672\,
            in3 => \N__50872\,
            lcout => OPEN,
            ltout => \spi_slave_inst.un1_spointer11_2_0_a2_0_6_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.rxdata_reg_i_RNIH2363_1_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__29229\,
            in1 => \N__29144\,
            in2 => \N__29220\,
            in3 => \N__29129\,
            lcout => un1_spointer11_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_5_3_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__40532\,
            in1 => \N__40334\,
            in2 => \N__46207\,
            in3 => \N__43145\,
            lcout => \sDAC_mem_22_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI5B15_1_1_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44958\,
            in2 => \_gnd_net_\,
            in3 => \N__44868\,
            lcout => \N_285\,
            ltout => \N_285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_18_3_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40531\,
            in1 => \N__40333\,
            in2 => \N__29199\,
            in3 => \N__43143\,
            lcout => \sDAC_mem_21_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_5_1_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__43144\,
            in1 => \N__46184\,
            in2 => \_gnd_net_\,
            in3 => \N__46068\,
            lcout => \sDAC_mem_29_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigInternal_RNO_1_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__46067\,
            in1 => \N__43260\,
            in2 => \N__29196\,
            in3 => \N__31090\,
            lcout => OPEN,
            ltout => \N_116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigInternal_RNO_0_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51078\,
            in2 => \N__29148\,
            in3 => \N__29040\,
            lcout => OPEN,
            ltout => \N_117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEETrigInternal_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29041\,
            in1 => \N__29145\,
            in2 => \N__29133\,
            in3 => \N__29130\,
            lcout => \sEETrigInternalZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47755\,
            ce => 'H',
            sr => \N__52998\
        );

    \sEEPoff_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51133\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPoffZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47767\,
            ce => \N__30975\,
            sr => \N__52991\
        );

    \sEEPoff_1_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50572\,
            lcout => \sEEPoffZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47767\,
            ce => \N__30975\,
            sr => \N__52991\
        );

    \sEEPoff_2_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50026\,
            lcout => \sEEPoffZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47767\,
            ce => \N__30975\,
            sr => \N__52991\
        );

    \sEEPoff_3_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49574\,
            lcout => \sEEPoffZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47767\,
            ce => \N__30975\,
            sr => \N__52991\
        );

    \sEEPoff_4_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49130\,
            lcout => \sEEPoffZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47767\,
            ce => \N__30975\,
            sr => \N__52991\
        );

    \sEEPoff_5_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47045\,
            lcout => \sEEPoffZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47767\,
            ce => \N__30975\,
            sr => \N__52991\
        );

    \sEEPoff_6_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48272\,
            lcout => \sEEPoffZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47767\,
            ce => \N__30975\,
            sr => \N__52991\
        );

    \sEEPoff_7_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48575\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPoffZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47767\,
            ce => \N__30975\,
            sr => \N__52991\
        );

    \sEEPoff_10_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50180\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPoffZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47781\,
            ce => \N__29337\,
            sr => \N__52986\
        );

    \sEEPoff_11_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49575\,
            lcout => \sEEPoffZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47781\,
            ce => \N__29337\,
            sr => \N__52986\
        );

    \sEEPoff_12_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49129\,
            lcout => \sEEPoffZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47781\,
            ce => \N__29337\,
            sr => \N__52986\
        );

    \sEEPoff_13_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47053\,
            lcout => \sEEPoffZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47781\,
            ce => \N__29337\,
            sr => \N__52986\
        );

    \sEEPoff_14_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48273\,
            lcout => \sEEPoffZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47781\,
            ce => \N__29337\,
            sr => \N__52986\
        );

    \sEEPoff_15_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEPoffZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47781\,
            ce => \N__29337\,
            sr => \N__52986\
        );

    \sEEPoff_8_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51079\,
            lcout => \sEEPoffZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47781\,
            ce => \N__29337\,
            sr => \N__52986\
        );

    \sEEPoff_9_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50573\,
            lcout => \sEEPoffZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47781\,
            ce => \N__29337\,
            sr => \N__52986\
        );

    \sCounterADC_0_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38225\,
            in1 => \N__38267\,
            in2 => \_gnd_net_\,
            in3 => \N__29322\,
            lcout => \sCounterADCZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \sCounterADC_cry_0\,
            clk => \N__47796\,
            ce => \N__29940\,
            sr => \N__52981\
        );

    \sCounterADC_1_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38203\,
            in1 => \N__38282\,
            in2 => \_gnd_net_\,
            in3 => \N__29319\,
            lcout => \sCounterADCZ0Z_1\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_0\,
            carryout => \sCounterADC_cry_1\,
            clk => \N__47796\,
            ce => \N__29940\,
            sr => \N__52981\
        );

    \sCounterADC_2_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38226\,
            in1 => \N__34350\,
            in2 => \_gnd_net_\,
            in3 => \N__29589\,
            lcout => \sCounterADCZ0Z_2\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_1\,
            carryout => \sCounterADC_cry_2\,
            clk => \N__47796\,
            ce => \N__29940\,
            sr => \N__52981\
        );

    \sCounterADC_3_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38204\,
            in1 => \N__34364\,
            in2 => \_gnd_net_\,
            in3 => \N__29586\,
            lcout => \sCounterADCZ0Z_3\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_2\,
            carryout => \sCounterADC_cry_3\,
            clk => \N__47796\,
            ce => \N__29940\,
            sr => \N__52981\
        );

    \sCounterADC_4_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38227\,
            in1 => \N__34304\,
            in2 => \_gnd_net_\,
            in3 => \N__29583\,
            lcout => \sCounterADCZ0Z_4\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_3\,
            carryout => \sCounterADC_cry_4\,
            clk => \N__47796\,
            ce => \N__29940\,
            sr => \N__52981\
        );

    \sCounterADC_5_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38205\,
            in1 => \N__34320\,
            in2 => \_gnd_net_\,
            in3 => \N__29580\,
            lcout => \sCounterADCZ0Z_5\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_4\,
            carryout => \sCounterADC_cry_5\,
            clk => \N__47796\,
            ce => \N__29940\,
            sr => \N__52981\
        );

    \sCounterADC_6_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38228\,
            in1 => \N__34274\,
            in2 => \_gnd_net_\,
            in3 => \N__29577\,
            lcout => \sCounterADCZ0Z_6\,
            ltout => OPEN,
            carryin => \sCounterADC_cry_5\,
            carryout => \sCounterADC_cry_6\,
            clk => \N__47796\,
            ce => \N__29940\,
            sr => \N__52981\
        );

    \sCounterADC_7_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38206\,
            in1 => \N__34259\,
            in2 => \_gnd_net_\,
            in3 => \N__29574\,
            lcout => \sCounterADCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47796\,
            ce => \N__29940\,
            sr => \N__52981\
        );

    \spi_data_miso_0_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__29571\,
            in1 => \N__29856\,
            in2 => \N__29547\,
            in3 => \N__29920\,
            lcout => \spi_data_misoZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47807\,
            ce => \N__29787\,
            sr => \N__52978\
        );

    \spi_data_miso_1_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__29921\,
            in1 => \N__29514\,
            in2 => \N__29869\,
            in3 => \N__29499\,
            lcout => \spi_data_misoZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47807\,
            ce => \N__29787\,
            sr => \N__52978\
        );

    \spi_data_miso_2_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__29469\,
            in1 => \N__29860\,
            in2 => \N__29445\,
            in3 => \N__29922\,
            lcout => \spi_data_misoZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47807\,
            ce => \N__29787\,
            sr => \N__52978\
        );

    \spi_data_miso_3_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__29923\,
            in1 => \N__30051\,
            in2 => \N__29870\,
            in3 => \N__30030\,
            lcout => \spi_data_misoZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47807\,
            ce => \N__29787\,
            sr => \N__52978\
        );

    \spi_data_miso_4_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__29997\,
            in1 => \N__29864\,
            in2 => \N__29976\,
            in3 => \N__29924\,
            lcout => \spi_data_misoZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47807\,
            ce => \N__29787\,
            sr => \N__52978\
        );

    \spi_data_miso_5_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__29925\,
            in1 => \N__29889\,
            in2 => \N__29871\,
            in3 => \N__29823\,
            lcout => \spi_data_misoZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47807\,
            ce => \N__29787\,
            sr => \N__52978\
        );

    \sRAM_ADD_0_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__31936\,
            in1 => \N__29763\,
            in2 => \N__31623\,
            in3 => \N__32184\,
            lcout => \RAM_ADD_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47816\,
            ce => \N__30262\,
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_23_c_RNIQQ6O1_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100110011"
        )
    port map (
            in0 => \N__32179\,
            in1 => \N__29718\,
            in2 => \N__29703\,
            in3 => \N__31934\,
            lcout => \N_67_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un4_sacqtime_cry_23_c_RNIJ7QO_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31935\,
            in1 => \N__29699\,
            in2 => \_gnd_net_\,
            in3 => \N__32180\,
            lcout => \N_31_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sRAM_ADD_1_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__32183\,
            in1 => \N__29688\,
            in2 => \N__31605\,
            in3 => \N__31941\,
            lcout => \RAM_ADD_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47816\,
            ce => \N__30262\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_10_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__31937\,
            in1 => \N__33096\,
            in2 => \N__29646\,
            in3 => \N__32185\,
            lcout => \RAM_ADD_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47816\,
            ce => \N__30262\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_11_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__32181\,
            in1 => \N__30405\,
            in2 => \N__33078\,
            in3 => \N__31939\,
            lcout => \RAM_ADD_c_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47816\,
            ce => \N__30262\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_12_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__31938\,
            in1 => \N__33057\,
            in2 => \N__30354\,
            in3 => \N__32186\,
            lcout => \RAM_ADD_c_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47816\,
            ce => \N__30262\,
            sr => \_gnd_net_\
        );

    \sRAM_ADD_13_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__32182\,
            in1 => \N__30309\,
            in2 => \N__33036\,
            in3 => \N__31940\,
            lcout => \RAM_ADD_c_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47816\,
            ce => \N__30262\,
            sr => \_gnd_net_\
        );

    \RAM_DATA_1_3_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30240\,
            lcout => \RAM_DATA_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => \N__31181\,
            sr => \N__52970\
        );

    \RAM_DATA_1_0_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30204\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RAM_DATA_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => \N__31181\,
            sr => \N__52970\
        );

    \RAM_DATA_1_5_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30165\,
            lcout => \RAM_DATA_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => \N__31181\,
            sr => \N__52970\
        );

    \RAM_DATA_1_1_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30123\,
            lcout => \RAM_DATA_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => \N__31181\,
            sr => \N__52970\
        );

    \RAM_DATA_1_8_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30090\,
            lcout => \RAM_DATA_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => \N__31181\,
            sr => \N__52970\
        );

    \RAM_DATA_1_9_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30639\,
            lcout => \RAM_DATA_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => \N__31181\,
            sr => \N__52970\
        );

    \RAM_DATA_1_15_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37903\,
            lcout => \RAM_DATA_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => \N__31181\,
            sr => \N__52970\
        );

    \RAM_DATA_1_7_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \RAM_DATA_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47824\,
            ce => \N__31181\,
            sr => \N__52970\
        );

    \RAM_DATA_cl_1_RNO_0_15_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__30539\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31711\,
            lcout => \N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_13_RNO_0_15_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30503\,
            in2 => \_gnd_net_\,
            in3 => \N__31710\,
            lcout => \N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_3_RNO_0_15_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30431\,
            in2 => \_gnd_net_\,
            in3 => \N__31713\,
            lcout => \N_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_2_RNO_0_15_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30470\,
            in2 => \_gnd_net_\,
            in3 => \N__31712\,
            lcout => \N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_3_15_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__30453\,
            in1 => \N__32153\,
            in2 => \N__32675\,
            in3 => \N__31973\,
            lcout => \RAM_DATA_cl_3Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47841\,
            ce => 'H',
            sr => \N__52967\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_0_LC_13_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38552\,
            in1 => \N__52592\,
            in2 => \_gnd_net_\,
            in3 => \N__30420\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30697\,
            ce => \N__30672\,
            sr => \N__53110\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_5_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30746\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30700\,
            ce => \N__30671\,
            sr => \N__53097\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_1_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30794\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30700\,
            ce => \N__30671\,
            sr => \N__53097\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_2_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30782\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30700\,
            ce => \N__30671\,
            sr => \N__53097\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_3_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30770\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30700\,
            ce => \N__30671\,
            sr => \N__53097\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_4_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30758\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30700\,
            ce => \N__30671\,
            sr => \N__53097\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_6_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30734\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30700\,
            ce => \N__30671\,
            sr => \N__53097\
        );

    \spi_slave_inst.rx_shift_data_pos_sclk_i_7_LC_13_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30722\,
            lcout => \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__30700\,
            ce => \N__30671\,
            sr => \N__53097\
        );

    \sDAC_mem_38_1_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50422\,
            lcout => \sDAC_mem_38Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47817\,
            ce => \N__41868\,
            sr => \N__53084\
        );

    \sDAC_mem_6_2_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50005\,
            lcout => \sDAC_mem_6Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47808\,
            ce => \N__43078\,
            sr => \N__53072\
        );

    \sDAC_mem_6_5_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46793\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_6Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47808\,
            ce => \N__43078\,
            sr => \N__53072\
        );

    \sDAC_mem_6_7_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48671\,
            lcout => \sDAC_mem_6Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47808\,
            ce => \N__43078\,
            sr => \N__53072\
        );

    \sDAC_mem_2_0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51024\,
            lcout => \sDAC_mem_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47797\,
            ce => \N__37407\,
            sr => \N__53060\
        );

    \sDAC_mem_2_1_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50625\,
            lcout => \sDAC_mem_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47797\,
            ce => \N__37407\,
            sr => \N__53060\
        );

    \sDAC_mem_2_2_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50006\,
            lcout => \sDAC_mem_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47797\,
            ce => \N__37407\,
            sr => \N__53060\
        );

    \sDAC_mem_2_3_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49496\,
            lcout => \sDAC_mem_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47797\,
            ce => \N__37407\,
            sr => \N__53060\
        );

    \sDAC_mem_2_4_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48989\,
            lcout => \sDAC_mem_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47797\,
            ce => \N__37407\,
            sr => \N__53060\
        );

    \sDAC_mem_2_5_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46794\,
            lcout => \sDAC_mem_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47797\,
            ce => \N__37407\,
            sr => \N__53060\
        );

    \sDAC_mem_2_6_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48062\,
            lcout => \sDAC_mem_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47797\,
            ce => \N__37407\,
            sr => \N__53060\
        );

    \sDAC_mem_2_7_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48670\,
            lcout => \sDAC_mem_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47797\,
            ce => \N__37407\,
            sr => \N__53060\
        );

    \sDAC_mem_22_1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50691\,
            lcout => \sDAC_mem_22Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47782\,
            ce => \N__39824\,
            sr => \N__53050\
        );

    \sDAC_data_RNO_21_5_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52007\,
            in1 => \N__30849\,
            in2 => \_gnd_net_\,
            in3 => \N__30843\,
            lcout => \sDAC_data_RNO_21Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_22_2_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50091\,
            lcout => \sDAC_mem_22Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47782\,
            ce => \N__39824\,
            sr => \N__53050\
        );

    \sDAC_data_RNO_21_6_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__30837\,
            in1 => \_gnd_net_\,
            in2 => \N__52118\,
            in3 => \N__30831\,
            lcout => \sDAC_data_RNO_21Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_22_3_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49590\,
            lcout => \sDAC_mem_22Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47782\,
            ce => \N__39824\,
            sr => \N__53050\
        );

    \sDAC_data_RNO_21_7_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52008\,
            in1 => \N__30825\,
            in2 => \_gnd_net_\,
            in3 => \N__30819\,
            lcout => \sDAC_data_RNO_21Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_22_4_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49077\,
            lcout => \sDAC_mem_22Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47782\,
            ce => \N__39824\,
            sr => \N__53050\
        );

    \sAddress_RNIAM2A_3_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__46438\,
            in1 => \N__40534\,
            in2 => \_gnd_net_\,
            in3 => \N__40347\,
            lcout => \N_291\,
            ltout => \N_291_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_6_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30906\,
            in2 => \N__30813\,
            in3 => \N__44730\,
            lcout => \sEEPonPoff_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_20_3_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30871\,
            in2 => \_gnd_net_\,
            in3 => \N__43160\,
            lcout => \sDAC_mem_17_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_0_5_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__30870\,
            in1 => \N__46512\,
            in2 => \_gnd_net_\,
            in3 => \N__46328\,
            lcout => \sDAC_mem_1_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_2_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__44957\,
            in1 => \N__40348\,
            in2 => \N__40555\,
            in3 => \N__30996\,
            lcout => \sAddress_RNIA6242Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIQ63A_0_6_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__30954\,
            in1 => \N__46511\,
            in2 => \N__30933\,
            in3 => \N__44644\,
            lcout => \sEEPonPoff_1_sqmuxa_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_21_3_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__44731\,
            in1 => \N__30873\,
            in2 => \_gnd_net_\,
            in3 => \N__31105\,
            lcout => \sEEPon_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_5_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30872\,
            in1 => \N__46513\,
            in2 => \_gnd_net_\,
            in3 => \N__46329\,
            lcout => \sDAC_mem_33_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_17_0_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51027\,
            lcout => \sDAC_mem_17Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47756\,
            ce => \N__30960\,
            sr => \N__53031\
        );

    \sDAC_mem_17_1_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50693\,
            lcout => \sDAC_mem_17Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47756\,
            ce => \N__30960\,
            sr => \N__53031\
        );

    \sDAC_mem_17_2_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50092\,
            lcout => \sDAC_mem_17Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47756\,
            ce => \N__30960\,
            sr => \N__53031\
        );

    \sDAC_mem_17_3_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49591\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_17Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47756\,
            ce => \N__30960\,
            sr => \N__53031\
        );

    \sDAC_mem_17_4_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49075\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_17Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47756\,
            ce => \N__30960\,
            sr => \N__53031\
        );

    \sDAC_mem_17_5_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46897\,
            lcout => \sDAC_mem_17Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47756\,
            ce => \N__30960\,
            sr => \N__53031\
        );

    \sDAC_mem_17_6_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48124\,
            lcout => \sDAC_mem_17Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47756\,
            ce => \N__30960\,
            sr => \N__53031\
        );

    \sDAC_mem_17_7_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48668\,
            lcout => \sDAC_mem_17Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47756\,
            ce => \N__30960\,
            sr => \N__53031\
        );

    \sDAC_mem_32_0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51132\,
            lcout => \sDAC_mem_32Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47742\,
            ce => \N__31113\,
            sr => \N__53021\
        );

    \sDAC_mem_32_1_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50694\,
            lcout => \sDAC_mem_32Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47742\,
            ce => \N__31113\,
            sr => \N__53021\
        );

    \sDAC_mem_32_2_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50093\,
            lcout => \sDAC_mem_32Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47742\,
            ce => \N__31113\,
            sr => \N__53021\
        );

    \sDAC_mem_32_3_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49592\,
            lcout => \sDAC_mem_32Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47742\,
            ce => \N__31113\,
            sr => \N__53021\
        );

    \sDAC_mem_32_4_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49078\,
            lcout => \sDAC_mem_32Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47742\,
            ce => \N__31113\,
            sr => \N__53021\
        );

    \sDAC_mem_32_5_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46898\,
            lcout => \sDAC_mem_32Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47742\,
            ce => \N__31113\,
            sr => \N__53021\
        );

    \sDAC_mem_32_6_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48254\,
            lcout => \sDAC_mem_32Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47742\,
            ce => \N__31113\,
            sr => \N__53021\
        );

    \sDAC_mem_32_7_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48669\,
            lcout => \sDAC_mem_32Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47742\,
            ce => \N__31113\,
            sr => \N__53021\
        );

    \sAddress_RNI9IH12_0_6_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__44694\,
            in1 => \N__46096\,
            in2 => \N__44595\,
            in3 => \N__31104\,
            lcout => \sEETrigCounter_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI5B15_3_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40495\,
            in2 => \_gnd_net_\,
            in3 => \N__40304\,
            lcout => \N_1480\,
            ltout => \N_1480_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_7_1_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001000"
        )
    port map (
            in0 => \N__43139\,
            in1 => \N__44592\,
            in2 => \N__30999\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_31_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_9_3_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__40512\,
            in1 => \N__40306\,
            in2 => \N__46450\,
            in3 => \N__43140\,
            lcout => \sDAC_mem_18_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIA6242_2_2_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__40305\,
            in1 => \N__44960\,
            in2 => \N__40533\,
            in3 => \N__30992\,
            lcout => \sAddress_RNIA6242_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIVREN1_0_4_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__46486\,
            in1 => \N__44637\,
            in2 => \N__44797\,
            in3 => \N__44693\,
            lcout => \N_280\,
            ltout => \N_280_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_3_3_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__44588\,
            in1 => \N__40511\,
            in2 => \N__30963\,
            in3 => \N__40335\,
            lcout => \sDAC_mem_24_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_14_3_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__40336\,
            in1 => \N__43269\,
            in2 => \N__40540\,
            in3 => \N__43138\,
            lcout => \sDAC_mem_19_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_19_0_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51134\,
            lcout => \sDAC_mem_19Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47743\,
            ce => \N__31122\,
            sr => \N__53010\
        );

    \sDAC_mem_19_1_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50574\,
            lcout => \sDAC_mem_19Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47743\,
            ce => \N__31122\,
            sr => \N__53010\
        );

    \sDAC_mem_19_2_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50179\,
            lcout => \sDAC_mem_19Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47743\,
            ce => \N__31122\,
            sr => \N__53010\
        );

    \sDAC_mem_19_3_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49702\,
            lcout => \sDAC_mem_19Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47743\,
            ce => \N__31122\,
            sr => \N__53010\
        );

    \sDAC_mem_19_4_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49145\,
            lcout => \sDAC_mem_19Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47743\,
            ce => \N__31122\,
            sr => \N__53010\
        );

    \sDAC_mem_19_5_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46993\,
            lcout => \sDAC_mem_19Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47743\,
            ce => \N__31122\,
            sr => \N__53010\
        );

    \sDAC_mem_19_6_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48236\,
            lcout => \sDAC_mem_19Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47743\,
            ce => \N__31122\,
            sr => \N__53010\
        );

    \sDAC_mem_19_7_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48817\,
            lcout => \sDAC_mem_19Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47743\,
            ce => \N__31122\,
            sr => \N__53010\
        );

    \sDAC_mem_18_3_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49703\,
            lcout => \sDAC_mem_18Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47757\,
            ce => \N__34089\,
            sr => \N__53002\
        );

    \sDAC_data_RNO_30_7_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__52150\,
            in1 => \N__31152\,
            in2 => \_gnd_net_\,
            in3 => \N__31158\,
            lcout => \sDAC_data_RNO_30Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_18_4_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49307\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_18Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47757\,
            ce => \N__34089\,
            sr => \N__53002\
        );

    \sDAC_data_RNO_30_8_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__52151\,
            in1 => \N__31140\,
            in2 => \_gnd_net_\,
            in3 => \N__31146\,
            lcout => \sDAC_data_RNO_30Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_18_5_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46994\,
            lcout => \sDAC_mem_18Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47757\,
            ce => \N__34089\,
            sr => \N__53002\
        );

    \sDAC_data_RNO_30_9_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__52152\,
            in1 => \N__31128\,
            in2 => \_gnd_net_\,
            in3 => \N__31134\,
            lcout => \sDAC_data_RNO_30Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_18_6_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48237\,
            lcout => \sDAC_mem_18Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47757\,
            ce => \N__34089\,
            sr => \N__53002\
        );

    \sDAC_mem_24_0_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51216\,
            lcout => \sDAC_mem_24Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47768\,
            ce => \N__39954\,
            sr => \N__52993\
        );

    \sDAC_mem_24_1_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50732\,
            lcout => \sDAC_mem_24Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47768\,
            ce => \N__39954\,
            sr => \N__52993\
        );

    \sDAC_mem_24_3_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49704\,
            lcout => \sDAC_mem_24Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47768\,
            ce => \N__39954\,
            sr => \N__52993\
        );

    \sDAC_mem_24_4_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49144\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_24Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47768\,
            ce => \N__39954\,
            sr => \N__52993\
        );

    \sDAC_mem_24_6_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48303\,
            lcout => \sDAC_mem_24Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47768\,
            ce => \N__39954\,
            sr => \N__52993\
        );

    \sEEACQ_10_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50257\,
            lcout => \sEEACQZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47783\,
            ce => \N__31170\,
            sr => \N__52988\
        );

    \sEEACQ_11_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49786\,
            lcout => \sEEACQZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47783\,
            ce => \N__31170\,
            sr => \N__52988\
        );

    \sEEACQ_12_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49226\,
            lcout => \sEEACQZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47783\,
            ce => \N__31170\,
            sr => \N__52988\
        );

    \sEEACQ_13_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47119\,
            lcout => \sEEACQZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47783\,
            ce => \N__31170\,
            sr => \N__52988\
        );

    \sEEACQ_14_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48304\,
            lcout => \sEEACQZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47783\,
            ce => \N__31170\,
            sr => \N__52988\
        );

    \sEEACQ_15_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48667\,
            lcout => \sEEACQZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47783\,
            ce => \N__31170\,
            sr => \N__52988\
        );

    \sEEACQ_8_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51262\,
            lcout => \sEEACQZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47783\,
            ce => \N__31170\,
            sr => \N__52988\
        );

    \sEEACQ_9_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50734\,
            lcout => \sEEACQZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47783\,
            ce => \N__31170\,
            sr => \N__52988\
        );

    \RAM_DATA_1_4_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RAM_DATA_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47798\,
            ce => \N__31182\,
            sr => \N__52983\
        );

    \RAM_DATA_1_6_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31554\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RAM_DATA_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47798\,
            ce => \N__31182\,
            sr => \N__52983\
        );

    \RAM_DATA_1_10_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31521\,
            lcout => \RAM_DATA_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47798\,
            ce => \N__31182\,
            sr => \N__52983\
        );

    \RAM_DATA_1_11_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31476\,
            lcout => \RAM_DATA_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47798\,
            ce => \N__31182\,
            sr => \N__52983\
        );

    \RAM_DATA_1_12_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RAM_DATA_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47798\,
            ce => \N__31182\,
            sr => \N__52983\
        );

    \RAM_DATA_1_13_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31389\,
            lcout => \RAM_DATA_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47798\,
            ce => \N__31182\,
            sr => \N__52983\
        );

    \RAM_DATA_1_14_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31301\,
            lcout => \RAM_DATA_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47798\,
            ce => \N__31182\,
            sr => \N__52983\
        );

    \RAM_DATA_1_2_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31215\,
            lcout => \RAM_DATA_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47798\,
            ce => \N__31182\,
            sr => \N__52983\
        );

    \RAM_DATA_cl_4_15_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__31629\,
            in1 => \N__32222\,
            in2 => \N__32546\,
            in3 => \N__31945\,
            lcout => \RAM_DATA_cl_4Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47809\,
            ce => 'H',
            sr => \N__52980\
        );

    \RAM_DATA_cl_5_RNO_0_15_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32735\,
            in2 => \_gnd_net_\,
            in3 => \N__31695\,
            lcout => OPEN,
            ltout => \N_107_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_5_15_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32493\,
            in1 => \N__32223\,
            in2 => \N__32757\,
            in3 => \N__31946\,
            lcout => \RAM_DATA_cl_5Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47809\,
            ce => 'H',
            sr => \N__52980\
        );

    \RAM_DATA_cl_6_RNO_0_15_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32702\,
            in2 => \_gnd_net_\,
            in3 => \N__31696\,
            lcout => OPEN,
            ltout => \N_108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_6_15_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32494\,
            in1 => \N__32224\,
            in2 => \N__32724\,
            in3 => \N__31947\,
            lcout => \RAM_DATA_cl_6Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47809\,
            ce => 'H',
            sr => \N__52980\
        );

    \RAM_DATA_cl_7_RNO_0_15_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31757\,
            in2 => \_gnd_net_\,
            in3 => \N__31697\,
            lcout => OPEN,
            ltout => \N_95_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RAM_DATA_cl_7_15_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32495\,
            in1 => \N__32225\,
            in2 => \N__31980\,
            in3 => \N__31948\,
            lcout => \RAM_DATA_cl_7Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47809\,
            ce => 'H',
            sr => \N__52980\
        );

    \RAM_DATA_cl_4_RNO_0_15_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31724\,
            in2 => \_gnd_net_\,
            in3 => \N__31694\,
            lcout => \N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sRAM_pointer_write_0_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33556\,
            in1 => \N__31619\,
            in2 => \_gnd_net_\,
            in3 => \N__31608\,
            lcout => \sRAM_pointer_writeZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \sRAM_pointer_write_cry_0\,
            clk => \N__47818\,
            ce => \N__33306\,
            sr => \N__52976\
        );

    \sRAM_pointer_write_1_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33552\,
            in1 => \N__31601\,
            in2 => \_gnd_net_\,
            in3 => \N__32928\,
            lcout => \sRAM_pointer_writeZ0Z_1\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_0\,
            carryout => \sRAM_pointer_write_cry_1\,
            clk => \N__47818\,
            ce => \N__33306\,
            sr => \N__52976\
        );

    \sRAM_pointer_write_2_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33557\,
            in1 => \N__32918\,
            in2 => \_gnd_net_\,
            in3 => \N__32907\,
            lcout => \sRAM_pointer_writeZ0Z_2\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_1\,
            carryout => \sRAM_pointer_write_cry_2\,
            clk => \N__47818\,
            ce => \N__33306\,
            sr => \N__52976\
        );

    \sRAM_pointer_write_3_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33553\,
            in1 => \N__32897\,
            in2 => \_gnd_net_\,
            in3 => \N__32886\,
            lcout => \sRAM_pointer_writeZ0Z_3\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_2\,
            carryout => \sRAM_pointer_write_cry_3\,
            clk => \N__47818\,
            ce => \N__33306\,
            sr => \N__52976\
        );

    \sRAM_pointer_write_4_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33558\,
            in1 => \N__32873\,
            in2 => \_gnd_net_\,
            in3 => \N__32862\,
            lcout => \sRAM_pointer_writeZ0Z_4\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_3\,
            carryout => \sRAM_pointer_write_cry_4\,
            clk => \N__47818\,
            ce => \N__33306\,
            sr => \N__52976\
        );

    \sRAM_pointer_write_5_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33554\,
            in1 => \N__32852\,
            in2 => \_gnd_net_\,
            in3 => \N__32841\,
            lcout => \sRAM_pointer_writeZ0Z_5\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_4\,
            carryout => \sRAM_pointer_write_cry_5\,
            clk => \N__47818\,
            ce => \N__33306\,
            sr => \N__52976\
        );

    \sRAM_pointer_write_6_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33559\,
            in1 => \N__32834\,
            in2 => \_gnd_net_\,
            in3 => \N__32823\,
            lcout => \sRAM_pointer_writeZ0Z_6\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_5\,
            carryout => \sRAM_pointer_write_cry_6\,
            clk => \N__47818\,
            ce => \N__33306\,
            sr => \N__52976\
        );

    \sRAM_pointer_write_7_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33555\,
            in1 => \N__32816\,
            in2 => \_gnd_net_\,
            in3 => \N__32805\,
            lcout => \sRAM_pointer_writeZ0Z_7\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_6\,
            carryout => \sRAM_pointer_write_cry_7\,
            clk => \N__47818\,
            ce => \N__33306\,
            sr => \N__52976\
        );

    \sRAM_pointer_write_8_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33567\,
            in1 => \N__32795\,
            in2 => \_gnd_net_\,
            in3 => \N__32784\,
            lcout => \sRAM_pointer_writeZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \sRAM_pointer_write_cry_8\,
            clk => \N__47825\,
            ce => \N__33305\,
            sr => \N__52973\
        );

    \sRAM_pointer_write_9_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33563\,
            in1 => \N__32771\,
            in2 => \_gnd_net_\,
            in3 => \N__32760\,
            lcout => \sRAM_pointer_writeZ0Z_9\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_8\,
            carryout => \sRAM_pointer_write_cry_9\,
            clk => \N__47825\,
            ce => \N__33305\,
            sr => \N__52973\
        );

    \sRAM_pointer_write_10_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33564\,
            in1 => \N__33092\,
            in2 => \_gnd_net_\,
            in3 => \N__33081\,
            lcout => \sRAM_pointer_writeZ0Z_10\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_9\,
            carryout => \sRAM_pointer_write_cry_10\,
            clk => \N__47825\,
            ce => \N__33305\,
            sr => \N__52973\
        );

    \sRAM_pointer_write_11_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33560\,
            in1 => \N__33071\,
            in2 => \_gnd_net_\,
            in3 => \N__33060\,
            lcout => \sRAM_pointer_writeZ0Z_11\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_10\,
            carryout => \sRAM_pointer_write_cry_11\,
            clk => \N__47825\,
            ce => \N__33305\,
            sr => \N__52973\
        );

    \sRAM_pointer_write_12_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33565\,
            in1 => \N__33050\,
            in2 => \_gnd_net_\,
            in3 => \N__33039\,
            lcout => \sRAM_pointer_writeZ0Z_12\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_11\,
            carryout => \sRAM_pointer_write_cry_12\,
            clk => \N__47825\,
            ce => \N__33305\,
            sr => \N__52973\
        );

    \sRAM_pointer_write_13_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33561\,
            in1 => \N__33029\,
            in2 => \_gnd_net_\,
            in3 => \N__33018\,
            lcout => \sRAM_pointer_writeZ0Z_13\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_12\,
            carryout => \sRAM_pointer_write_cry_13\,
            clk => \N__47825\,
            ce => \N__33305\,
            sr => \N__52973\
        );

    \sRAM_pointer_write_14_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33566\,
            in1 => \N__33008\,
            in2 => \_gnd_net_\,
            in3 => \N__32997\,
            lcout => \sRAM_pointer_writeZ0Z_14\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_13\,
            carryout => \sRAM_pointer_write_cry_14\,
            clk => \N__47825\,
            ce => \N__33305\,
            sr => \N__52973\
        );

    \sRAM_pointer_write_15_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33562\,
            in1 => \N__32987\,
            in2 => \_gnd_net_\,
            in3 => \N__32976\,
            lcout => \sRAM_pointer_writeZ0Z_15\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_14\,
            carryout => \sRAM_pointer_write_cry_15\,
            clk => \N__47825\,
            ce => \N__33305\,
            sr => \N__52973\
        );

    \sRAM_pointer_write_16_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33542\,
            in1 => \N__32969\,
            in2 => \_gnd_net_\,
            in3 => \N__32955\,
            lcout => \sRAM_pointer_writeZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => \sRAM_pointer_write_cry_16\,
            clk => \N__47835\,
            ce => \N__33304\,
            sr => \N__52969\
        );

    \sRAM_pointer_write_17_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33541\,
            in1 => \N__32942\,
            in2 => \_gnd_net_\,
            in3 => \N__32931\,
            lcout => \sRAM_pointer_writeZ0Z_17\,
            ltout => OPEN,
            carryin => \sRAM_pointer_write_cry_16\,
            carryout => \sRAM_pointer_write_cry_17\,
            clk => \N__47835\,
            ce => \N__33304\,
            sr => \N__52969\
        );

    \sRAM_pointer_write_18_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33543\,
            in1 => \N__33320\,
            in2 => \_gnd_net_\,
            in3 => \N__33330\,
            lcout => \sRAM_pointer_writeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47835\,
            ce => \N__33304\,
            sr => \N__52969\
        );

    \sDAC_mem_pointer_RNIF3GH_6_LC_14_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37272\,
            in2 => \_gnd_net_\,
            in3 => \N__37278\,
            lcout => un17_sdacdyn_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1_1_LC_14_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001101"
        )
    port map (
            in0 => \N__33277\,
            in1 => \N__38553\,
            in2 => \N__37188\,
            in3 => \N__52415\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNIOASC_5_LC_14_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__37103\,
            in1 => \N__37118\,
            in2 => \N__37244\,
            in3 => \N__37343\,
            lcout => OPEN,
            ltout => \spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNI1DAJ_1_LC_14_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__37138\,
            in1 => \_gnd_net_\,
            in2 => \N__33234\,
            in3 => \N__37207\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_i6\,
            ltout => \spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_done_neg_sclk_i_LC_14_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33213\,
            in2 => \N__33162\,
            in3 => \N__33149\,
            lcout => \spi_slave_inst.tx_done_neg_sclk_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi_slave_inst.tx_done_neg_sclk_iC_net\,
            ce => 'H',
            sr => \N__53125\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNIKKJ63_0_LC_14_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__38554\,
            in1 => \N__38594\,
            in2 => \N__33138\,
            in3 => \N__52314\,
            lcout => spi_miso_rpi_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_13_3_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52156\,
            in1 => \N__41661\,
            in2 => \N__43666\,
            in3 => \N__33606\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_3_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52161\,
            in1 => \N__40068\,
            in2 => \N__33099\,
            in3 => \N__37296\,
            lcout => \sDAC_data_RNO_5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_6_0_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50986\,
            lcout => \sDAC_mem_6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47810\,
            ce => \N__43071\,
            sr => \N__53098\
        );

    \sDAC_data_RNO_13_4_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52160\,
            in1 => \N__33600\,
            in2 => \N__43668\,
            in3 => \N__33591\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_4_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52157\,
            in1 => \N__40059\,
            in2 => \N__33594\,
            in3 => \N__37290\,
            lcout => \sDAC_data_RNO_5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_6_1_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50600\,
            lcout => \sDAC_mem_6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47810\,
            ce => \N__43071\,
            sr => \N__53098\
        );

    \sDAC_data_RNO_13_5_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52158\,
            in1 => \N__41646\,
            in2 => \N__43667\,
            in3 => \N__33585\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_5_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__40182\,
            in1 => \N__52159\,
            in2 => \N__33579\,
            in3 => \N__37368\,
            lcout => \sDAC_data_RNO_5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_12_5_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__51910\,
            in1 => \N__38733\,
            in2 => \N__43673\,
            in3 => \N__33573\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_5_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52138\,
            in1 => \N__38769\,
            in2 => \N__33576\,
            in3 => \N__37359\,
            lcout => \sDAC_data_RNO_4Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_4_2_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50106\,
            lcout => \sDAC_mem_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47799\,
            ce => \N__39627\,
            sr => \N__53085\
        );

    \sDAC_data_RNO_12_6_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52137\,
            in1 => \N__38721\,
            in2 => \N__43671\,
            in3 => \N__33648\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_6_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51907\,
            in1 => \N__38760\,
            in2 => \N__33651\,
            in3 => \N__37353\,
            lcout => \sDAC_data_RNO_4Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_4_3_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47799\,
            ce => \N__39627\,
            sr => \N__53085\
        );

    \sDAC_data_RNO_12_7_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__51908\,
            in1 => \N__38709\,
            in2 => \N__43672\,
            in3 => \N__33642\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_7_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__37413\,
            in1 => \N__38751\,
            in2 => \N__33630\,
            in3 => \N__51909\,
            lcout => \sDAC_data_RNO_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_3_0_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51040\,
            lcout => \sDAC_mem_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47784\,
            ce => \N__42960\,
            sr => \N__53073\
        );

    \sDAC_data_RNO_28_3_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__43606\,
            in1 => \N__51902\,
            in2 => \N__33627\,
            in3 => \N__37332\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_3_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51903\,
            in1 => \N__40230\,
            in2 => \N__33618\,
            in3 => \N__33615\,
            lcout => \sDAC_data_RNO_15Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_5_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43607\,
            in1 => \N__44184\,
            in2 => \_gnd_net_\,
            in3 => \N__44319\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_5_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__51904\,
            in1 => \_gnd_net_\,
            in2 => \N__33609\,
            in3 => \N__45207\,
            lcout => \sDAC_data_RNO_8Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_5_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__38742\,
            in1 => \N__51905\,
            in2 => \N__43665\,
            in3 => \N__41832\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_5_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51906\,
            in1 => \N__43974\,
            in2 => \N__33717\,
            in3 => \N__47193\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_7Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_5_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101100010"
        )
    port map (
            in0 => \N__45874\,
            in1 => \N__34065\,
            in2 => \N__33714\,
            in3 => \N__33711\,
            lcout => \sDAC_data_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_5_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__33705\,
            in1 => \N__41919\,
            in2 => \N__45908\,
            in3 => \N__33693\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_10Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_5_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__42528\,
            in1 => \N__42638\,
            in2 => \N__33696\,
            in3 => \N__38412\,
            lcout => \sDAC_data_2_41_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_5_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__45861\,
            in1 => \N__45518\,
            in2 => \N__36681\,
            in3 => \N__34104\,
            lcout => \sDAC_data_2_32_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_5_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__45519\,
            in1 => \N__45865\,
            in2 => \N__33918\,
            in3 => \N__33738\,
            lcout => OPEN,
            ltout => \sDAC_data_2_14_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_5_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__33687\,
            in1 => \N__45866\,
            in2 => \N__33678\,
            in3 => \N__33675\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_5_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__42529\,
            in1 => \N__33666\,
            in2 => \N__33660\,
            in3 => \N__33657\,
            lcout => OPEN,
            ltout => \sDAC_data_2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_5_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45990\,
            in2 => \N__33771\,
            in3 => \N__42381\,
            lcout => \sDAC_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53248\,
            ce => \N__42230\,
            sr => \N__53061\
        );

    \sDAC_mem_3_2_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47758\,
            ce => \N__42977\,
            sr => \N__53051\
        );

    \sDAC_data_RNO_28_5_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__51815\,
            in1 => \N__37320\,
            in2 => \N__43621\,
            in3 => \N__33756\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_5_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51818\,
            in1 => \N__40221\,
            in2 => \N__33747\,
            in3 => \N__33744\,
            lcout => \sDAC_data_RNO_15Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_7_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__51814\,
            in1 => \N__41808\,
            in2 => \N__43620\,
            in3 => \N__38829\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_7_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51817\,
            in1 => \N__44259\,
            in2 => \N__33732\,
            in3 => \N__47166\,
            lcout => \sDAC_data_RNO_7Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_7_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43542\,
            in1 => \N__44157\,
            in2 => \_gnd_net_\,
            in3 => \N__44292\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_7_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51816\,
            in2 => \N__33729\,
            in3 => \N__45180\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_8Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_7_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011000110010"
        )
    port map (
            in0 => \N__45783\,
            in1 => \N__43914\,
            in2 => \N__33726\,
            in3 => \N__33723\,
            lcout => \sDAC_data_RNO_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_27_8_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__43520\,
            in1 => \N__51555\,
            in2 => \N__33834\,
            in3 => \N__33849\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_27Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_8_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__33864\,
            in1 => \_gnd_net_\,
            in2 => \N__33852\,
            in3 => \N__33840\,
            lcout => \sDAC_data_RNO_14Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_26_8_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__43518\,
            in1 => \N__51553\,
            in2 => \N__33833\,
            in3 => \N__33848\,
            lcout => \sDAC_data_RNO_26Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_1_5_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47016\,
            lcout => \sDAC_mem_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47744\,
            ce => \N__42032\,
            sr => \N__53041\
        );

    \sDAC_data_RNO_26_9_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__43519\,
            in1 => \N__51554\,
            in2 => \N__33804\,
            in3 => \N__33780\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_9_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33819\,
            in2 => \N__33807\,
            in3 => \N__33786\,
            lcout => \sDAC_data_RNO_14Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_27_9_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__43517\,
            in1 => \N__51552\,
            in2 => \N__33803\,
            in3 => \N__33779\,
            lcout => \sDAC_data_RNO_27Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_1_6_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48233\,
            lcout => \sDAC_mem_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47744\,
            ce => \N__42032\,
            sr => \N__53041\
        );

    \sDAC_mem_3_6_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48255\,
            lcout => \sDAC_mem_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47733\,
            ce => \N__42978\,
            sr => \N__53032\
        );

    \sDAC_data_RNO_28_9_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__43514\,
            in1 => \N__51599\,
            in2 => \N__34008\,
            in3 => \N__37308\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_9_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51601\,
            in1 => \N__40722\,
            in2 => \N__33993\,
            in3 => \N__33990\,
            lcout => \sDAC_data_RNO_15Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_26_4_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__43515\,
            in1 => \N__51600\,
            in2 => \N__33969\,
            in3 => \N__33947\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_4_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33984\,
            in2 => \N__33972\,
            in3 => \N__33939\,
            lcout => \sDAC_data_RNO_14Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_27_4_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__43513\,
            in1 => \N__51598\,
            in2 => \N__33968\,
            in3 => \N__33948\,
            lcout => \sDAC_data_RNO_27Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_26_5_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__51602\,
            in1 => \N__43516\,
            in2 => \N__33906\,
            in3 => \N__33891\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_5_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__33933\,
            in1 => \_gnd_net_\,
            in2 => \N__33921\,
            in3 => \N__33873\,
            lcout => \sDAC_data_RNO_14Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_27_3_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__43501\,
            in1 => \N__52083\,
            in2 => \N__39296\,
            in3 => \N__39263\,
            lcout => \sDAC_data_RNO_27Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_27_5_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__52082\,
            in1 => \N__33902\,
            in2 => \N__43550\,
            in3 => \N__33890\,
            lcout => \sDAC_data_RNO_27Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_10_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43502\,
            in1 => \N__44355\,
            in2 => \_gnd_net_\,
            in3 => \N__34038\,
            lcout => \sDAC_data_RNO_17Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_pointer_RNIAIV21_3_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__52081\,
            in1 => \N__45639\,
            in2 => \N__42614\,
            in3 => \N__45372\,
            lcout => OPEN,
            ltout => \op_le_op_le_un15_sdacdynlt4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_pointer_RNI4LV52_4_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000000"
        )
    port map (
            in0 => \N__43500\,
            in1 => \N__42447\,
            in2 => \N__34050\,
            in3 => \N__34047\,
            lcout => un17_sdacdyn_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_10_7_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48777\,
            lcout => \sDAC_mem_10Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47724\,
            ce => \N__45000\,
            sr => \N__53022\
        );

    \sDAC_data_RNO_9_10_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001011111"
        )
    port map (
            in0 => \N__47274\,
            in1 => \N__51288\,
            in2 => \N__45807\,
            in3 => \N__45373\,
            lcout => \sDAC_data_2_24_ns_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_30_10_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34026\,
            in1 => \N__51597\,
            in2 => \_gnd_net_\,
            in3 => \N__34032\,
            lcout => \sDAC_data_RNO_30Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_18_7_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48816\,
            lcout => \sDAC_mem_18Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47734\,
            ce => \N__34088\,
            sr => \N__53017\
        );

    \sDAC_data_RNO_30_3_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34014\,
            in1 => \N__51596\,
            in2 => \_gnd_net_\,
            in3 => \N__34020\,
            lcout => \sDAC_data_RNO_30Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_18_0_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51246\,
            lcout => \sDAC_mem_18Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47734\,
            ce => \N__34088\,
            sr => \N__53017\
        );

    \sDAC_data_RNO_30_4_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51594\,
            in2 => \N__34125\,
            in3 => \N__34116\,
            lcout => \sDAC_data_RNO_30Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_18_1_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50575\,
            lcout => \sDAC_mem_18Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47734\,
            ce => \N__34088\,
            sr => \N__53017\
        );

    \sDAC_data_RNO_30_5_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34095\,
            in1 => \N__51595\,
            in2 => \_gnd_net_\,
            in3 => \N__34110\,
            lcout => \sDAC_data_RNO_30Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_18_2_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50261\,
            lcout => \sDAC_mem_18Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47734\,
            ce => \N__34088\,
            sr => \N__53017\
        );

    \sDAC_data_RNO_19_5_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43740\,
            in1 => \N__51865\,
            in2 => \_gnd_net_\,
            in3 => \N__45090\,
            lcout => \sDAC_data_RNO_19Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_5_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51866\,
            in1 => \N__49857\,
            in2 => \_gnd_net_\,
            in3 => \N__34137\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_5_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110011101"
        )
    port map (
            in0 => \N__45421\,
            in1 => \N__45859\,
            in2 => \N__34074\,
            in3 => \N__34071\,
            lcout => \sDAC_data_2_24_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_6_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51867\,
            in1 => \N__49383\,
            in2 => \_gnd_net_\,
            in3 => \N__34131\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_6_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110011101"
        )
    port map (
            in0 => \N__45422\,
            in1 => \N__45860\,
            in2 => \N__34053\,
            in3 => \N__34143\,
            lcout => \sDAC_data_2_24_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_19_6_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51864\,
            in1 => \N__45075\,
            in2 => \_gnd_net_\,
            in3 => \N__43728\,
            lcout => \sDAC_data_RNO_19Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_12_2_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50105\,
            lcout => \sDAC_mem_12Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47745\,
            ce => \N__47384\,
            sr => \N__53011\
        );

    \sDAC_mem_12_3_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49795\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_12Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47745\,
            ce => \N__47384\,
            sr => \N__53011\
        );

    \sDAC_mem_31_0_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51261\,
            lcout => \sDAC_mem_31Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47759\,
            ce => \N__34380\,
            sr => \N__53003\
        );

    \sDAC_mem_31_1_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50733\,
            lcout => \sDAC_mem_31Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47759\,
            ce => \N__34380\,
            sr => \N__53003\
        );

    \sDAC_mem_31_2_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50262\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_31Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47759\,
            ce => \N__34380\,
            sr => \N__53003\
        );

    \sDAC_mem_31_3_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49796\,
            lcout => \sDAC_mem_31Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47759\,
            ce => \N__34380\,
            sr => \N__53003\
        );

    \sDAC_mem_31_4_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49222\,
            lcout => \sDAC_mem_31Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47759\,
            ce => \N__34380\,
            sr => \N__53003\
        );

    \sDAC_mem_31_5_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47073\,
            lcout => \sDAC_mem_31Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47759\,
            ce => \N__34380\,
            sr => \N__53003\
        );

    \sDAC_mem_31_6_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48324\,
            lcout => \sDAC_mem_31Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47759\,
            ce => \N__34380\,
            sr => \N__53003\
        );

    \sDAC_mem_31_7_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48842\,
            lcout => \sDAC_mem_31Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47759\,
            ce => \N__34380\,
            sr => \N__53003\
        );

    \sEEADC_freq_RNI4KIA1_2_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__34335\,
            in1 => \N__34365\,
            in2 => \N__34329\,
            in3 => \N__34349\,
            lcout => \un11_sacqtime_NE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEADC_freq_2_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50264\,
            lcout => \sEEADC_freqZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47769\,
            ce => \N__44127\,
            sr => \_gnd_net_\
        );

    \sEEADC_freq_3_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEADC_freqZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47769\,
            ce => \N__44127\,
            sr => \_gnd_net_\
        );

    \sEEADC_freq_RNICSIA1_4_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__34290\,
            in1 => \N__34319\,
            in2 => \N__34284\,
            in3 => \N__34305\,
            lcout => \un11_sacqtime_NE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEADC_freq_4_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49165\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEADC_freqZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47769\,
            ce => \N__44127\,
            sr => \_gnd_net_\
        );

    \sEEADC_freq_5_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47126\,
            lcout => \sEEADC_freqZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47769\,
            ce => \N__44127\,
            sr => \_gnd_net_\
        );

    \sEEADC_freq_RNIK4JA1_6_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__34275\,
            in1 => \N__41451\,
            in2 => \N__41442\,
            in3 => \N__34260\,
            lcout => \un11_sacqtime_NE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_0_c_inv_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35088\,
            in2 => \N__34244\,
            in3 => \N__34161\,
            lcout => \sEEACQ_i_0\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => un5_sdacdyn_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_1_c_inv_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35082\,
            in1 => \N__35062\,
            in2 => \N__34977\,
            in3 => \_gnd_net_\,
            lcout => \sEEACQ_i_1\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_0,
            carryout => un5_sdacdyn_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_2_c_inv_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34956\,
            in2 => \N__34866\,
            in3 => \N__34884\,
            lcout => \sEEACQ_i_2\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_1,
            carryout => un5_sdacdyn_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_3_c_inv_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34856\,
            in2 => \N__34761\,
            in3 => \N__34779\,
            lcout => \sEEACQ_i_3\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_2,
            carryout => un5_sdacdyn_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_4_c_inv_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34752\,
            in1 => \N__34734\,
            in2 => \N__36884\,
            in3 => \_gnd_net_\,
            lcout => \sEEACQ_i_4\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_3,
            carryout => un5_sdacdyn_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_5_c_inv_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34726\,
            in2 => \N__34629\,
            in3 => \N__34647\,
            lcout => \sEEACQ_i_5\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_4,
            carryout => un5_sdacdyn_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_6_c_inv_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34612\,
            in2 => \N__34503\,
            in3 => \N__34521\,
            lcout => \sEEACQ_i_6\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_5,
            carryout => un5_sdacdyn_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_7_c_inv_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34386\,
            in2 => \N__34493\,
            in3 => \N__34404\,
            lcout => \sEEACQ_i_7\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_6,
            carryout => un5_sdacdyn_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_8_c_inv_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35775\,
            in2 => \N__35888\,
            in3 => \N__35793\,
            lcout => \sEEACQ_i_8\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => un5_sdacdyn_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_9_c_inv_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35769\,
            in2 => \N__35664\,
            in3 => \N__35682\,
            lcout => \sEEACQ_i_9\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_8,
            carryout => un5_sdacdyn_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_10_c_inv_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35646\,
            in2 => \N__35550\,
            in3 => \N__35571\,
            lcout => \sEEACQ_i_10\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_9,
            carryout => un5_sdacdyn_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_11_c_inv_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35540\,
            in2 => \N__35445\,
            in3 => \N__35463\,
            lcout => \sEEACQ_i_11\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_10,
            carryout => un5_sdacdyn_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_12_c_inv_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35436\,
            in1 => \N__35409\,
            in2 => \N__35328\,
            in3 => \_gnd_net_\,
            lcout => \sEEACQ_i_12\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_11,
            carryout => un5_sdacdyn_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_13_c_inv_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35214\,
            in2 => \N__35319\,
            in3 => \N__35235\,
            lcout => \sEEACQ_i_13\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_12,
            carryout => un5_sdacdyn_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_14_c_inv_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35203\,
            in2 => \N__35097\,
            in3 => \N__35115\,
            lcout => \sEEACQ_i_14\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_13,
            carryout => un5_sdacdyn_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_15_c_inv_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36660\,
            in2 => \N__36555\,
            in3 => \N__36573\,
            lcout => \sEEACQ_i_15\,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_14,
            carryout => un5_sdacdyn_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_16_c_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36541\,
            in2 => \N__38075\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => un5_sdacdyn_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_17_c_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36442\,
            in2 => \N__38079\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_16,
            carryout => un5_sdacdyn_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_18_c_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36347\,
            in2 => \N__38076\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_17,
            carryout => un5_sdacdyn_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_19_c_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36255\,
            in2 => \N__38080\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_18,
            carryout => un5_sdacdyn_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_20_c_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36170\,
            in2 => \N__38077\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_19,
            carryout => un5_sdacdyn_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_21_c_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36081\,
            in2 => \N__38081\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_20,
            carryout => un5_sdacdyn_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_22_c_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35994\,
            in2 => \N__38078\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_21,
            carryout => un5_sdacdyn_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_23_c_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37087\,
            in2 => \N__38082\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_sdacdyn_cry_22,
            carryout => un5_sdacdyn_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_sdacdyn_cry_23_c_RNIELG28_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__36993\,
            in1 => \N__36978\,
            in2 => \N__36888\,
            in3 => \N__36723\,
            lcout => \un5_sdacdyn_cry_23_c_RNIELGZ0Z28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_pointer_0_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__51541\,
            in1 => \N__42298\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_pointerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53278\,
            ce => \N__42232\,
            sr => \N__52977\
        );

    \sDAC_data_RNO_31_6_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51540\,
            in1 => \N__36720\,
            in2 => \_gnd_net_\,
            in3 => \N__40098\,
            lcout => \sDAC_data_RNO_31Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_31_9_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36708\,
            in1 => \N__51539\,
            in2 => \_gnd_net_\,
            in3 => \N__40107\,
            lcout => \sDAC_data_RNO_31Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_32_3_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51537\,
            in1 => \N__45261\,
            in2 => \_gnd_net_\,
            in3 => \N__38112\,
            lcout => \sDAC_data_RNO_32Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_32_9_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51538\,
            in1 => \N__41487\,
            in2 => \_gnd_net_\,
            in3 => \N__38094\,
            lcout => \sDAC_data_RNO_32Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_16_7_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48808\,
            lcout => \sDAC_mem_16Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47826\,
            ce => \N__46635\,
            sr => \N__52974\
        );

    \sDAC_mem_16_0_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51276\,
            lcout => \sDAC_mem_16Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47826\,
            ce => \N__46635\,
            sr => \N__52974\
        );

    \sDAC_data_RNO_29_5_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36696\,
            in1 => \N__51480\,
            in2 => \_gnd_net_\,
            in3 => \N__37284\,
            lcout => \sDAC_data_RNO_29Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_16_2_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50310\,
            lcout => \sDAC_mem_16Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47826\,
            ce => \N__46635\,
            sr => \N__52974\
        );

    \sDAC_mem_pointer_6_LC_15_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_mem_pointerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53242\,
            ce => \N__42231\,
            sr => \N__53137\
        );

    \sDAC_mem_pointer_7_LC_15_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_mem_pointerZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53242\,
            ce => \N__42231\,
            sr => \N__53137\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_0_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37186\,
            in1 => \N__37240\,
            in2 => \N__37266\,
            in3 => \N__37265\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_2_0_\,
            carryout => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0\,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53132\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_1_LC_15_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37185\,
            in1 => \N__37208\,
            in2 => \_gnd_net_\,
            in3 => \N__37191\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0\,
            carryout => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1\,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53132\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_2_LC_15_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37187\,
            in1 => \N__37139\,
            in2 => \_gnd_net_\,
            in3 => \N__37122\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1\,
            carryout => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2\,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53132\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_3_LC_15_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37119\,
            in2 => \_gnd_net_\,
            in3 => \N__37107\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2\,
            carryout => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3\,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53132\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_4_LC_15_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37104\,
            in2 => \_gnd_net_\,
            in3 => \N__37092\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4\,
            ltout => OPEN,
            carryin => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3\,
            carryout => \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4\,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53132\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_5_LC_15_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37344\,
            in2 => \_gnd_net_\,
            in3 => \N__37347\,
            lcout => \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net\,
            ce => 'H',
            sr => \N__53132\
        );

    \sDAC_mem_34_0_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50882\,
            lcout => \sDAC_mem_34Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__40089\,
            sr => \N__53126\
        );

    \sDAC_mem_34_2_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50004\,
            lcout => \sDAC_mem_34Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__40089\,
            sr => \N__53126\
        );

    \sDAC_mem_34_4_LC_15_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49188\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_34Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__40089\,
            sr => \N__53126\
        );

    \sDAC_mem_34_5_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46769\,
            lcout => \sDAC_mem_34Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__40089\,
            sr => \N__53126\
        );

    \sDAC_mem_34_6_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_34Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__40089\,
            sr => \N__53126\
        );

    \sDAC_mem_34_7_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48545\,
            lcout => \sDAC_mem_34Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47811\,
            ce => \N__40089\,
            sr => \N__53126\
        );

    \sDAC_mem_7_0_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50987\,
            lcout => \sDAC_mem_7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47800\,
            ce => \N__37383\,
            sr => \N__53111\
        );

    \sDAC_mem_7_1_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50601\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_7Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47800\,
            ce => \N__37383\,
            sr => \N__53111\
        );

    \sDAC_mem_7_2_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50107\,
            lcout => \sDAC_mem_7Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47800\,
            ce => \N__37383\,
            sr => \N__53111\
        );

    \sDAC_mem_7_3_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49609\,
            lcout => \sDAC_mem_7Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47800\,
            ce => \N__37383\,
            sr => \N__53111\
        );

    \sDAC_mem_7_4_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_7Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47800\,
            ce => \N__37383\,
            sr => \N__53111\
        );

    \sDAC_mem_7_5_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46876\,
            lcout => \sDAC_mem_7Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47800\,
            ce => \N__37383\,
            sr => \N__53111\
        );

    \sDAC_mem_7_6_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48189\,
            lcout => \sDAC_mem_7Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47800\,
            ce => \N__37383\,
            sr => \N__53111\
        );

    \sDAC_mem_7_7_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48746\,
            lcout => \sDAC_mem_7Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47800\,
            ce => \N__37383\,
            sr => \N__53111\
        );

    \sDAC_mem_5_0_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51099\,
            lcout => \sDAC_mem_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47785\,
            ce => \N__37395\,
            sr => \N__53099\
        );

    \sDAC_mem_5_1_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50685\,
            lcout => \sDAC_mem_5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47785\,
            ce => \N__37395\,
            sr => \N__53099\
        );

    \sDAC_mem_5_2_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50108\,
            lcout => \sDAC_mem_5Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47785\,
            ce => \N__37395\,
            sr => \N__53099\
        );

    \sDAC_mem_5_3_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49610\,
            lcout => \sDAC_mem_5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47785\,
            ce => \N__37395\,
            sr => \N__53099\
        );

    \sDAC_mem_5_4_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47785\,
            ce => \N__37395\,
            sr => \N__53099\
        );

    \sDAC_mem_5_5_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46878\,
            lcout => \sDAC_mem_5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47785\,
            ce => \N__37395\,
            sr => \N__53099\
        );

    \sDAC_mem_5_6_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48191\,
            lcout => \sDAC_mem_5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47785\,
            ce => \N__37395\,
            sr => \N__53099\
        );

    \sDAC_mem_5_7_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48747\,
            lcout => \sDAC_mem_5Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47785\,
            ce => \N__37395\,
            sr => \N__53099\
        );

    \sAddress_RNI9IH12_10_3_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__40584\,
            in1 => \N__40398\,
            in2 => \N__46449\,
            in3 => \N__37494\,
            lcout => \sDAC_mem_2_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_17_3_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__37490\,
            in1 => \N__40585\,
            in2 => \N__46246\,
            in3 => \N__40401\,
            lcout => \sDAC_mem_5_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_15_3_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40583\,
            in1 => \N__40397\,
            in2 => \N__44586\,
            in3 => \N__37489\,
            lcout => \sDAC_mem_7_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_2_3_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__37492\,
            in1 => \N__40586\,
            in2 => \N__44587\,
            in3 => \N__40402\,
            lcout => \sDAC_mem_8_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_19_3_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__43282\,
            in1 => \N__40396\,
            in2 => \N__40604\,
            in3 => \N__37491\,
            lcout => \sDAC_mem_3_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_4_3_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__37493\,
            in1 => \N__40582\,
            in2 => \N__46245\,
            in3 => \N__40399\,
            lcout => \sDAC_mem_6_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIVREN1_1_4_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__46528\,
            in1 => \N__44645\,
            in2 => \N__44808\,
            in3 => \N__44741\,
            lcout => \N_279\,
            ltout => \N_279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_6_3_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__40575\,
            in1 => \N__40400\,
            in2 => \N__37473\,
            in3 => \N__43283\,
            lcout => \sDAC_mem_4_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_7_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__37470\,
            in1 => \N__38790\,
            in2 => \N__45875\,
            in3 => \N__38862\,
            lcout => \sDAC_data_RNO_10Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_7_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__45803\,
            in1 => \N__45520\,
            in2 => \N__42093\,
            in3 => \N__39072\,
            lcout => OPEN,
            ltout => \sDAC_data_2_14_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_7_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__45867\,
            in1 => \N__38892\,
            in2 => \N__37461\,
            in3 => \N__37458\,
            lcout => \sDAC_data_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_7_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010101110101"
        )
    port map (
            in0 => \N__42631\,
            in1 => \N__38469\,
            in2 => \N__42534\,
            in3 => \N__37449\,
            lcout => OPEN,
            ltout => \sDAC_data_2_41_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_7_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111000001110"
        )
    port map (
            in0 => \N__42518\,
            in1 => \N__37443\,
            in2 => \N__37437\,
            in3 => \N__37434\,
            lcout => OPEN,
            ltout => \sDAC_data_2_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_7_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__45960\,
            in1 => \_gnd_net_\,
            in2 => \N__37428\,
            in3 => \N__42382\,
            lcout => \sDAC_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53252\,
            ce => \N__42229\,
            sr => \N__53074\
        );

    \sDAC_data_RNO_17_9_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43581\,
            in1 => \N__44367\,
            in2 => \_gnd_net_\,
            in3 => \N__44271\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_9_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51808\,
            in2 => \N__37539\,
            in3 => \N__45156\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_8Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_9_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011000110010"
        )
    port map (
            in0 => \N__45751\,
            in1 => \N__38295\,
            in2 => \N__37536\,
            in3 => \N__37530\,
            lcout => \sDAC_data_RNO_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_3_4_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49260\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47746\,
            ce => \N__42961\,
            sr => \N__53062\
        );

    \sDAC_data_RNO_16_9_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__38817\,
            in1 => \N__43580\,
            in2 => \N__52012\,
            in3 => \N__41796\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_9_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52119\,
            in1 => \N__44232\,
            in2 => \N__37533\,
            in3 => \N__46650\,
            lcout => \sDAC_data_RNO_7Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_29_7_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37524\,
            in1 => \N__52014\,
            in2 => \_gnd_net_\,
            in3 => \N__37515\,
            lcout => \sDAC_data_RNO_29Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_16_4_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49360\,
            lcout => \sDAC_mem_16Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47735\,
            ce => \N__46629\,
            sr => \N__53052\
        );

    \sDAC_data_RNO_29_8_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37509\,
            in1 => \N__52013\,
            in2 => \_gnd_net_\,
            in3 => \N__37500\,
            lcout => \sDAC_data_RNO_29Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_16_5_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47017\,
            lcout => \sDAC_mem_16Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47735\,
            ce => \N__46629\,
            sr => \N__53052\
        );

    \sDAC_data_RNO_29_9_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37569\,
            in1 => \N__52015\,
            in2 => \_gnd_net_\,
            in3 => \N__37560\,
            lcout => \sDAC_data_RNO_29Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_16_6_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48234\,
            lcout => \sDAC_mem_16Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47735\,
            ce => \N__46629\,
            sr => \N__53052\
        );

    \sDAC_mem_pointer_RNI3NFH_1_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52041\,
            in2 => \N__45491\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_10_0_\,
            carryout => \sDAC_mem_pointer_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_pointer_2_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__42373\,
            in1 => \N__45717\,
            in2 => \_gnd_net_\,
            in3 => \N__37554\,
            lcout => \sDAC_mem_pointerZ0Z_2\,
            ltout => OPEN,
            carryin => \sDAC_mem_pointer_0_cry_1\,
            carryout => \sDAC_mem_pointer_0_cry_2\,
            clk => \N__53254\,
            ce => \N__42225\,
            sr => \N__53042\
        );

    \sDAC_mem_pointer_3_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__42376\,
            in1 => \N__42623\,
            in2 => \_gnd_net_\,
            in3 => \N__37551\,
            lcout => \sDAC_mem_pointerZ0Z_3\,
            ltout => OPEN,
            carryin => \sDAC_mem_pointer_0_cry_2\,
            carryout => \sDAC_mem_pointer_0_cry_3\,
            clk => \N__53254\,
            ce => \N__42225\,
            sr => \N__53042\
        );

    \sDAC_mem_pointer_4_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__42374\,
            in1 => \N__42483\,
            in2 => \_gnd_net_\,
            in3 => \N__37548\,
            lcout => \sDAC_mem_pointerZ0Z_4\,
            ltout => OPEN,
            carryin => \sDAC_mem_pointer_0_cry_3\,
            carryout => \sDAC_mem_pointer_0_cry_4\,
            clk => \N__53254\,
            ce => \N__42225\,
            sr => \N__53042\
        );

    \sDAC_mem_pointer_5_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__43479\,
            in1 => \N__42375\,
            in2 => \_gnd_net_\,
            in3 => \N__37545\,
            lcout => \sDAC_mem_pointerZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53254\,
            ce => \N__42225\,
            sr => \N__53042\
        );

    \sDAC_data_RNO_23_9_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52017\,
            in1 => \N__38355\,
            in2 => \_gnd_net_\,
            in3 => \N__37629\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_23Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_9_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__45709\,
            in1 => \N__38169\,
            in2 => \N__37542\,
            in3 => \N__38121\,
            lcout => \sDAC_data_RNO_11Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_10_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37653\,
            in1 => \N__52019\,
            in2 => \_gnd_net_\,
            in3 => \N__45141\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_8Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_10_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011000110010"
        )
    port map (
            in0 => \N__45710\,
            in1 => \N__37647\,
            in2 => \N__37641\,
            in3 => \N__37635\,
            lcout => \sDAC_data_RNO_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_10_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52016\,
            in1 => \N__41997\,
            in2 => \N__43575\,
            in3 => \N__38808\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_10_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52018\,
            in1 => \N__44220\,
            in2 => \N__37638\,
            in3 => \N__47340\,
            lcout => \sDAC_data_RNO_7Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_28_6_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48310\,
            lcout => \sDAC_mem_28Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47718\,
            ce => \N__41772\,
            sr => \N__53033\
        );

    \sDAC_mem_pointer_1_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__45424\,
            in1 => \N__52064\,
            in2 => \_gnd_net_\,
            in3 => \N__42379\,
            lcout => \sDAC_mem_pointerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53263\,
            ce => \N__42228\,
            sr => \N__53023\
        );

    \sDAC_data_1_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53263\,
            ce => \N__42228\,
            sr => \N__53023\
        );

    \sDAC_data_11_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53263\,
            ce => \N__42228\,
            sr => \N__53023\
        );

    \sDAC_data_12_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38018\,
            lcout => \sDAC_dataZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53263\,
            ce => \N__42228\,
            sr => \N__53023\
        );

    \sDAC_data_13_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__38019\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_dataZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53263\,
            ce => \N__42228\,
            sr => \N__53023\
        );

    \sDAC_data_14_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53263\,
            ce => \N__42228\,
            sr => \N__53023\
        );

    \sDAC_data_15_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \GNDG0\,
            lcout => \sDAC_dataZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53263\,
            ce => \N__42228\,
            sr => \N__53023\
        );

    \sDAC_data_RNO_31_8_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40128\,
            in1 => \N__51880\,
            in2 => \_gnd_net_\,
            in3 => \N__38157\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_31Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_25_8_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__45848\,
            in1 => \N__45415\,
            in2 => \N__37683\,
            in3 => \N__37677\,
            lcout => OPEN,
            ltout => \sDAC_data_2_39_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_8_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__45828\,
            in1 => \N__37659\,
            in2 => \N__37680\,
            in3 => \N__37671\,
            lcout => \sDAC_data_RNO_11Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_32_8_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51878\,
            in1 => \N__41499\,
            in2 => \_gnd_net_\,
            in3 => \N__38100\,
            lcout => \sDAC_data_RNO_32Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_8_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51881\,
            in1 => \N__38364\,
            in2 => \_gnd_net_\,
            in3 => \N__41511\,
            lcout => \sDAC_data_RNO_23Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_8_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51879\,
            in1 => \N__37665\,
            in2 => \_gnd_net_\,
            in3 => \N__39708\,
            lcout => \sDAC_data_RNO_24Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_24_5_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47117\,
            lcout => \sDAC_mem_24Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47736\,
            ce => \N__39971\,
            sr => \N__53018\
        );

    \sDAC_data_RNO_25_9_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__45847\,
            in1 => \N__45414\,
            in2 => \N__38151\,
            in3 => \N__38133\,
            lcout => \sDAC_data_2_39_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_26_0_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51247\,
            lcout => \sDAC_mem_26Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47747\,
            ce => \N__39528\,
            sr => \N__53012\
        );

    \sDAC_mem_26_1_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50723\,
            lcout => \sDAC_mem_26Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47747\,
            ce => \N__39528\,
            sr => \N__53012\
        );

    \sDAC_mem_26_2_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50263\,
            lcout => \sDAC_mem_26Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47747\,
            ce => \N__39528\,
            sr => \N__53012\
        );

    \sDAC_mem_26_3_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49797\,
            lcout => \sDAC_mem_26Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47747\,
            ce => \N__39528\,
            sr => \N__53012\
        );

    \sDAC_mem_26_4_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49177\,
            lcout => \sDAC_mem_26Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47747\,
            ce => \N__39528\,
            sr => \N__53012\
        );

    \sDAC_mem_26_5_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47074\,
            lcout => \sDAC_mem_26Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47747\,
            ce => \N__39528\,
            sr => \N__53012\
        );

    \sDAC_mem_26_6_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48311\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_26Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47747\,
            ce => \N__39528\,
            sr => \N__53012\
        );

    \sDAC_mem_26_7_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48843\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_26Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47747\,
            ce => \N__39528\,
            sr => \N__53012\
        );

    \sDAC_data_RNO_19_9_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52112\,
            in1 => \N__45036\,
            in2 => \_gnd_net_\,
            in3 => \N__43947\,
            lcout => \sDAC_data_RNO_19Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_9_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52114\,
            in1 => \N__45234\,
            in2 => \_gnd_net_\,
            in3 => \N__47868\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_9_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__45736\,
            in1 => \N__45439\,
            in2 => \N__38304\,
            in3 => \N__38301\,
            lcout => \sDAC_data_2_24_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEADC_freq_RNISBIA1_0_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__41460\,
            in1 => \N__38283\,
            in2 => \N__44142\,
            in3 => \N__38268\,
            lcout => OPEN,
            ltout => \un11_sacqtime_NE_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEADC_freq_RNI01BA5_0_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__38253\,
            in1 => \N__38247\,
            in2 => \N__38241\,
            in3 => \N__38238\,
            lcout => \un11_sacqtime_NE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_9_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38175\,
            in1 => \N__52113\,
            in2 => \_gnd_net_\,
            in3 => \N__39699\,
            lcout => \sDAC_data_RNO_24Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_29_0_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51253\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_29Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47770\,
            ce => \N__38346\,
            sr => \N__52994\
        );

    \sDAC_mem_29_1_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50754\,
            lcout => \sDAC_mem_29Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47770\,
            ce => \N__38346\,
            sr => \N__52994\
        );

    \sDAC_mem_29_2_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50300\,
            lcout => \sDAC_mem_29Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47770\,
            ce => \N__38346\,
            sr => \N__52994\
        );

    \sDAC_mem_29_3_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49835\,
            lcout => \sDAC_mem_29Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47770\,
            ce => \N__38346\,
            sr => \N__52994\
        );

    \sDAC_mem_29_4_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49326\,
            lcout => \sDAC_mem_29Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47770\,
            ce => \N__38346\,
            sr => \N__52994\
        );

    \sDAC_mem_29_5_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__47134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_29Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47770\,
            ce => \N__38346\,
            sr => \N__52994\
        );

    \sDAC_mem_29_6_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48337\,
            lcout => \sDAC_mem_29Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47770\,
            ce => \N__38346\,
            sr => \N__52994\
        );

    \sDAC_mem_29_7_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48830\,
            lcout => \sDAC_mem_29Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47770\,
            ce => \N__38346\,
            sr => \N__52994\
        );

    \sDAC_data_RNO_11_6_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__38424\,
            in1 => \N__38325\,
            in2 => \N__45841\,
            in3 => \N__38664\,
            lcout => \sDAC_data_RNO_11Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_6_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52075\,
            in1 => \N__38331\,
            in2 => \_gnd_net_\,
            in3 => \N__38457\,
            lcout => \sDAC_data_RNO_23Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_31_7_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51892\,
            in1 => \N__38319\,
            in2 => \_gnd_net_\,
            in3 => \N__39897\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_31Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_25_7_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__45440\,
            in1 => \N__45746\,
            in2 => \N__38307\,
            in3 => \N__38442\,
            lcout => OPEN,
            ltout => \sDAC_data_2_39_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_7_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__39744\,
            in1 => \N__45750\,
            in2 => \N__38472\,
            in3 => \N__38649\,
            lcout => \sDAC_data_RNO_11Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_28_3_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_28Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47786\,
            ce => \N__41778\,
            sr => \N__52989\
        );

    \sDAC_data_RNO_32_7_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51891\,
            in1 => \N__41226\,
            in2 => \_gnd_net_\,
            in3 => \N__38451\,
            lcout => \sDAC_data_RNO_32Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_6_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52074\,
            in1 => \N__38436\,
            in2 => \_gnd_net_\,
            in3 => \N__39720\,
            lcout => \sDAC_data_RNO_24Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_31_5_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51495\,
            in1 => \N__38679\,
            in2 => \_gnd_net_\,
            in3 => \N__40134\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_31Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_25_5_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__45734\,
            in1 => \N__45521\,
            in2 => \N__38418\,
            in3 => \N__38388\,
            lcout => OPEN,
            ltout => \sDAC_data_2_39_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_5_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__45737\,
            in1 => \N__38685\,
            in2 => \N__38415\,
            in3 => \N__38370\,
            lcout => \sDAC_data_RNO_11Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_32_5_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41256\,
            in1 => \N__51493\,
            in2 => \_gnd_net_\,
            in3 => \N__38397\,
            lcout => \sDAC_data_RNO_32Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_5_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51494\,
            in1 => \N__38379\,
            in2 => \_gnd_net_\,
            in3 => \N__41535\,
            lcout => \sDAC_data_RNO_23Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_5_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51501\,
            in1 => \N__38697\,
            in2 => \_gnd_net_\,
            in3 => \N__39729\,
            lcout => \sDAC_data_RNO_24Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_24_2_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50301\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_24Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47801\,
            ce => \N__39972\,
            sr => \N__52984\
        );

    \sDAC_data_RNO_25_6_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__45735\,
            in1 => \N__45522\,
            in2 => \N__38673\,
            in3 => \N__38631\,
            lcout => \sDAC_data_2_39_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_7_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51502\,
            in1 => \N__38658\,
            in2 => \_gnd_net_\,
            in3 => \N__41523\,
            lcout => \sDAC_data_RNO_23Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_32_6_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51478\,
            in1 => \N__41241\,
            in2 => \_gnd_net_\,
            in3 => \N__38640\,
            lcout => \sDAC_data_RNO_32Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_31_3_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__38625\,
            in1 => \N__51477\,
            in2 => \_gnd_net_\,
            in3 => \N__40113\,
            lcout => \sDAC_data_RNO_31Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_29_6_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51479\,
            in1 => \N__38610\,
            in2 => \_gnd_net_\,
            in3 => \N__44055\,
            lcout => \sDAC_data_RNO_29Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ00Q2_0_LC_16_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__38595\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38563\,
            lcout => spi_miso_ft_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_8_3_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__40613\,
            in1 => \N__40641\,
            in2 => \N__46452\,
            in3 => \N__40417\,
            lcout => \sDAC_mem_34_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_36_0_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51082\,
            lcout => \sDAC_mem_36Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47787\,
            ce => \N__40656\,
            sr => \N__53127\
        );

    \sDAC_mem_36_1_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50677\,
            lcout => \sDAC_mem_36Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47787\,
            ce => \N__40656\,
            sr => \N__53127\
        );

    \sDAC_mem_36_2_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50151\,
            lcout => \sDAC_mem_36Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47787\,
            ce => \N__40656\,
            sr => \N__53127\
        );

    \sDAC_mem_36_3_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49661\,
            lcout => \sDAC_mem_36Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47787\,
            ce => \N__40656\,
            sr => \N__53127\
        );

    \sDAC_mem_36_4_LC_16_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49109\,
            lcout => \sDAC_mem_36Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47787\,
            ce => \N__40656\,
            sr => \N__53127\
        );

    \sDAC_mem_36_5_LC_16_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46877\,
            lcout => \sDAC_mem_36Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47787\,
            ce => \N__40656\,
            sr => \N__53127\
        );

    \sDAC_mem_36_6_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48190\,
            lcout => \sDAC_mem_36Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47787\,
            ce => \N__40656\,
            sr => \N__53127\
        );

    \sDAC_mem_36_7_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48737\,
            lcout => \sDAC_mem_36Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47787\,
            ce => \N__40656\,
            sr => \N__53127\
        );

    \sDAC_mem_37_0_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51100\,
            lcout => \sDAC_mem_37Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47771\,
            ce => \N__40149\,
            sr => \N__53112\
        );

    \sDAC_mem_37_1_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50686\,
            lcout => \sDAC_mem_37Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47771\,
            ce => \N__40149\,
            sr => \N__53112\
        );

    \sDAC_mem_37_2_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50240\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_37Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47771\,
            ce => \N__40149\,
            sr => \N__53112\
        );

    \sDAC_mem_37_3_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49765\,
            lcout => \sDAC_mem_37Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47771\,
            ce => \N__40149\,
            sr => \N__53112\
        );

    \sDAC_mem_37_4_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49110\,
            lcout => \sDAC_mem_37Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47771\,
            ce => \N__40149\,
            sr => \N__53112\
        );

    \sDAC_mem_37_5_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46879\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_37Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47771\,
            ce => \N__40149\,
            sr => \N__53112\
        );

    \sDAC_mem_37_6_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48192\,
            lcout => \sDAC_mem_37Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47771\,
            ce => \N__40149\,
            sr => \N__53112\
        );

    \sDAC_mem_37_7_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48738\,
            lcout => \sDAC_mem_37Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47771\,
            ce => \N__40149\,
            sr => \N__53112\
        );

    \sDAC_mem_8_0_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51101\,
            lcout => \sDAC_mem_8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47760\,
            ce => \N__38796\,
            sr => \N__53100\
        );

    \sDAC_mem_8_1_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50687\,
            lcout => \sDAC_mem_8Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47760\,
            ce => \N__38796\,
            sr => \N__53100\
        );

    \sDAC_mem_8_2_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50241\,
            lcout => \sDAC_mem_8Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47760\,
            ce => \N__38796\,
            sr => \N__53100\
        );

    \sDAC_mem_8_3_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49766\,
            lcout => \sDAC_mem_8Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47760\,
            ce => \N__38796\,
            sr => \N__53100\
        );

    \sDAC_mem_8_4_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49358\,
            lcout => \sDAC_mem_8Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47760\,
            ce => \N__38796\,
            sr => \N__53100\
        );

    \sDAC_mem_8_5_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46880\,
            lcout => \sDAC_mem_8Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47760\,
            ce => \N__38796\,
            sr => \N__53100\
        );

    \sDAC_mem_8_6_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48211\,
            lcout => \sDAC_mem_8Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47760\,
            ce => \N__38796\,
            sr => \N__53100\
        );

    \sDAC_mem_8_7_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48740\,
            lcout => \sDAC_mem_8Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47760\,
            ce => \N__38796\,
            sr => \N__53100\
        );

    \sDAC_data_RNO_20_7_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52002\,
            in1 => \N__40704\,
            in2 => \_gnd_net_\,
            in3 => \N__38781\,
            lcout => \sDAC_data_RNO_20Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_20_4_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49111\,
            lcout => \sDAC_mem_20Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47748\,
            ce => \N__44029\,
            sr => \N__53086\
        );

    \sDAC_data_RNO_20_8_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40698\,
            in1 => \N__51999\,
            in2 => \_gnd_net_\,
            in3 => \N__38775\,
            lcout => \sDAC_data_RNO_20Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_20_5_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46881\,
            lcout => \sDAC_mem_20Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47748\,
            ce => \N__44029\,
            sr => \N__53086\
        );

    \sDAC_data_RNO_20_9_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52001\,
            in1 => \N__40692\,
            in2 => \_gnd_net_\,
            in3 => \N__38961\,
            lcout => \sDAC_data_RNO_20Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_20_6_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48212\,
            lcout => \sDAC_mem_20Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47748\,
            ce => \N__44029\,
            sr => \N__53086\
        );

    \sDAC_data_RNO_21_10_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52000\,
            in1 => \N__38955\,
            in2 => \_gnd_net_\,
            in3 => \N__38946\,
            lcout => \sDAC_data_RNO_21Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_21_3_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51998\,
            in1 => \N__38931\,
            in2 => \_gnd_net_\,
            in3 => \N__38922\,
            lcout => \sDAC_data_RNO_21Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_13_7_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52122\,
            in1 => \N__41625\,
            in2 => \N__43669\,
            in3 => \N__40824\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_7_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51811\,
            in1 => \N__40173\,
            in2 => \N__38907\,
            in3 => \N__38904\,
            lcout => \sDAC_data_RNO_5Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_7_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__45490\,
            in1 => \N__45799\,
            in2 => \N__38886\,
            in3 => \N__38868\,
            lcout => \sDAC_data_2_32_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_7_3_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__40416\,
            in1 => \N__43281\,
            in2 => \N__40603\,
            in3 => \N__43190\,
            lcout => \sDAC_mem_20_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_28_7_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__51809\,
            in1 => \N__43624\,
            in2 => \N__38856\,
            in3 => \N__38841\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_7_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__39081\,
            in1 => \N__51810\,
            in2 => \N__39075\,
            in3 => \N__40209\,
            lcout => \sDAC_data_RNO_15Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_12_8_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52116\,
            in1 => \N__39066\,
            in2 => \N__43565\,
            in3 => \N__39033\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_8_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52105\,
            in1 => \N__39057\,
            in2 => \N__39048\,
            in3 => \N__39045\,
            lcout => \sDAC_data_RNO_4Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_4_5_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47088\,
            lcout => \sDAC_mem_4Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47725\,
            ce => \N__39631\,
            sr => \N__53063\
        );

    \sDAC_data_RNO_12_9_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52106\,
            in1 => \N__39027\,
            in2 => \N__43686\,
            in3 => \N__38994\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_9_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52117\,
            in1 => \N__39018\,
            in2 => \N__39009\,
            in3 => \N__39006\,
            lcout => \sDAC_data_RNO_4Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_4_6_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48235\,
            lcout => \sDAC_mem_4Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47725\,
            ce => \N__39631\,
            sr => \N__53063\
        );

    \sDAC_data_RNO_13_10_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52115\,
            in1 => \N__41880\,
            in2 => \N__43564\,
            in3 => \N__38988\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_10_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52104\,
            in1 => \N__40161\,
            in2 => \N__38976\,
            in3 => \N__38973\,
            lcout => \sDAC_data_RNO_5Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_9_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__42726\,
            in1 => \N__39195\,
            in2 => \N__45808\,
            in3 => \N__39132\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_9_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__42517\,
            in1 => \N__39189\,
            in2 => \N__39177\,
            in3 => \N__39087\,
            lcout => OPEN,
            ltout => \sDAC_data_2_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_9_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47250\,
            in2 => \N__39174\,
            in3 => \N__42380\,
            lcout => \sDAC_dataZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53257\,
            ce => \N__42222\,
            sr => \N__53053\
        );

    \sDAC_data_RNO_6_9_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__45533\,
            in1 => \N__45712\,
            in2 => \N__39156\,
            in3 => \N__39144\,
            lcout => \sDAC_data_2_14_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_9_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__45711\,
            in1 => \N__39126\,
            in2 => \N__45534\,
            in3 => \N__39120\,
            lcout => OPEN,
            ltout => \sDAC_data_2_32_ns_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_9_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__45716\,
            in1 => \N__39843\,
            in2 => \N__39108\,
            in3 => \N__39105\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_10Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_9_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__42479\,
            in1 => \N__42610\,
            in2 => \N__39096\,
            in3 => \N__39093\,
            lcout => \sDAC_data_2_41_ns_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_3_5_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47089\,
            lcout => \sDAC_mem_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47713\,
            ce => \N__42984\,
            sr => \N__53043\
        );

    \sDAC_data_RNO_28_8_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__43450\,
            in1 => \N__52092\,
            in2 => \N__39399\,
            in3 => \N__39384\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_8_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52093\,
            in1 => \N__40194\,
            in2 => \N__39369\,
            in3 => \N__39366\,
            lcout => \sDAC_data_RNO_15Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_26_10_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__43449\,
            in1 => \N__52094\,
            in2 => \N__39342\,
            in3 => \N__39320\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_10_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39360\,
            in2 => \N__39345\,
            in3 => \N__39306\,
            lcout => \sDAC_data_RNO_14Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_27_10_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__43448\,
            in1 => \N__52091\,
            in2 => \N__39341\,
            in3 => \N__39321\,
            lcout => \sDAC_data_RNO_27Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_26_3_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__52095\,
            in1 => \N__43451\,
            in2 => \N__39300\,
            in3 => \N__39270\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_3_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39252\,
            in2 => \N__39237\,
            in3 => \N__39234\,
            lcout => \sDAC_data_RNO_14Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_10_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__39537\,
            in1 => \N__39225\,
            in2 => \N__45882\,
            in3 => \N__39201\,
            lcout => \sDAC_data_RNO_10Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_10_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__45728\,
            in1 => \N__45423\,
            in2 => \N__39213\,
            in3 => \N__41322\,
            lcout => \sDAC_data_2_32_ns_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_10_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__39513\,
            in1 => \N__45729\,
            in2 => \N__42849\,
            in3 => \N__45523\,
            lcout => OPEN,
            ltout => \sDAC_data_2_14_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_10_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__45730\,
            in1 => \N__39504\,
            in2 => \N__39495\,
            in3 => \N__39411\,
            lcout => \sDAC_data_RNO_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_10_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001110111"
        )
    port map (
            in0 => \N__42532\,
            in1 => \N__39492\,
            in2 => \N__40044\,
            in3 => \N__42630\,
            lcout => OPEN,
            ltout => \sDAC_data_2_41_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_10_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111000001110"
        )
    port map (
            in0 => \N__42533\,
            in1 => \N__39486\,
            in2 => \N__39480\,
            in3 => \N__39477\,
            lcout => OPEN,
            ltout => \sDAC_data_2_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_10_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46587\,
            in2 => \N__39471\,
            in3 => \N__42378\,
            lcout => \sDAC_dataZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53268\,
            ce => \N__42227\,
            sr => \N__53034\
        );

    \sDAC_data_RNO_12_10_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__51971\,
            in1 => \N__39450\,
            in2 => \N__43634\,
            in3 => \N__39405\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_10_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51996\,
            in1 => \N__39438\,
            in2 => \N__39426\,
            in3 => \N__39423\,
            lcout => \sDAC_data_RNO_4Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_4_7_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47726\,
            ce => \N__39639\,
            sr => \N__53024\
        );

    \sDAC_data_RNO_12_3_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__51997\,
            in1 => \N__39687\,
            in2 => \N__43635\,
            in3 => \N__39645\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_3_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51972\,
            in1 => \N__39675\,
            in2 => \N__39660\,
            in3 => \N__39657\,
            lcout => \sDAC_data_RNO_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_4_0_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51252\,
            lcout => \sDAC_mem_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47726\,
            ce => \N__39639\,
            sr => \N__53024\
        );

    \sDAC_data_RNO_12_4_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__51970\,
            in1 => \N__39597\,
            in2 => \N__43633\,
            in3 => \N__39588\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_am_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_4_4_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__51995\,
            in1 => \N__39570\,
            in2 => \N__39555\,
            in3 => \N__39552\,
            lcout => \sDAC_data_RNO_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_20_10_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51985\,
            in1 => \N__40686\,
            in2 => \_gnd_net_\,
            in3 => \N__44046\,
            lcout => \sDAC_data_RNO_20Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_4_1_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__44410\,
            in1 => \N__46244\,
            in2 => \_gnd_net_\,
            in3 => \N__43179\,
            lcout => \sDAC_mem_30_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_2_1_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__43178\,
            in1 => \N__44409\,
            in2 => \_gnd_net_\,
            in3 => \N__43254\,
            lcout => \sDAC_mem_28_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_0_1_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__44411\,
            in1 => \N__46418\,
            in2 => \_gnd_net_\,
            in3 => \N__43177\,
            lcout => \sDAC_mem_26_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI5B15_0_3_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40541\,
            in2 => \_gnd_net_\,
            in3 => \N__40359\,
            lcout => \N_142\,
            ltout => \N_142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_rpi_ibuf_RNIRGF52_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46243\,
            in2 => \N__39732\,
            in3 => \N__46044\,
            lcout => \sEEADC_freq_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_30_0_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51248\,
            lcout => \sDAC_mem_30Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47749\,
            ce => \N__39693\,
            sr => \N__53013\
        );

    \sDAC_mem_30_1_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50724\,
            lcout => \sDAC_mem_30Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47749\,
            ce => \N__39693\,
            sr => \N__53013\
        );

    \sDAC_mem_30_2_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50178\,
            lcout => \sDAC_mem_30Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47749\,
            ce => \N__39693\,
            sr => \N__53013\
        );

    \sDAC_mem_30_3_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49836\,
            lcout => \sDAC_mem_30Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47749\,
            ce => \N__39693\,
            sr => \N__53013\
        );

    \sDAC_mem_30_4_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49091\,
            lcout => \sDAC_mem_30Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47749\,
            ce => \N__39693\,
            sr => \N__53013\
        );

    \sDAC_mem_30_5_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47135\,
            lcout => \sDAC_mem_30Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47749\,
            ce => \N__39693\,
            sr => \N__53013\
        );

    \sDAC_mem_30_6_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48338\,
            lcout => \sDAC_mem_30Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47749\,
            ce => \N__39693\,
            sr => \N__53013\
        );

    \sDAC_mem_30_7_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48831\,
            lcout => \sDAC_mem_30Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47749\,
            ce => \N__39693\,
            sr => \N__53013\
        );

    \sDAC_data_RNO_21_8_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51888\,
            in1 => \N__39885\,
            in2 => \_gnd_net_\,
            in3 => \N__39867\,
            lcout => \sDAC_data_RNO_21Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_22_5_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47136\,
            lcout => \sDAC_mem_22Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47761\,
            ce => \N__39825\,
            sr => \N__53004\
        );

    \sDAC_data_RNO_21_9_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51889\,
            in1 => \N__39861\,
            in2 => \_gnd_net_\,
            in3 => \N__39831\,
            lcout => \sDAC_data_RNO_21Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_22_6_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48339\,
            lcout => \sDAC_mem_22Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47761\,
            ce => \N__39825\,
            sr => \N__53004\
        );

    \sDAC_data_RNO_23_4_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39786\,
            in1 => \N__51886\,
            in2 => \_gnd_net_\,
            in3 => \N__41541\,
            lcout => \sDAC_data_RNO_23Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_4_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51887\,
            in1 => \N__39780\,
            in2 => \_gnd_net_\,
            in3 => \N__39774\,
            lcout => \sDAC_data_RNO_24Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_7_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51885\,
            in1 => \N__39762\,
            in2 => \_gnd_net_\,
            in3 => \N__39750\,
            lcout => \sDAC_data_RNO_24Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_31_10_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51895\,
            in1 => \N__39978\,
            in2 => \_gnd_net_\,
            in3 => \N__39891\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_31Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_25_10_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__45877\,
            in1 => \N__45481\,
            in2 => \N__39735\,
            in3 => \N__40023\,
            lcout => OPEN,
            ltout => \sDAC_data_2_39_ns_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_10_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__45878\,
            in1 => \N__39984\,
            in2 => \N__40047\,
            in3 => \N__40011\,
            lcout => \sDAC_data_RNO_11Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_32_10_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51893\,
            in2 => \N__41472\,
            in3 => \N__40032\,
            lcout => \sDAC_data_RNO_32Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_10_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51894\,
            in1 => \N__40017\,
            in2 => \_gnd_net_\,
            in3 => \N__41784\,
            lcout => \sDAC_data_RNO_23Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_10_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51896\,
            in1 => \N__40005\,
            in2 => \_gnd_net_\,
            in3 => \N__39993\,
            lcout => \sDAC_data_RNO_24Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_24_7_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48799\,
            lcout => \sDAC_mem_24Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47772\,
            ce => \N__39967\,
            sr => \N__52995\
        );

    \sDAC_data_RNO_25_3_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__45876\,
            in1 => \N__45480\,
            in2 => \N__39921\,
            in3 => \N__39906\,
            lcout => \sDAC_data_2_39_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_25_4_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49327\,
            lcout => \sDAC_mem_25Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47788\,
            ce => \N__41723\,
            sr => \N__52990\
        );

    \sDAC_mem_25_7_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48801\,
            lcout => \sDAC_mem_25Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47788\,
            ce => \N__41723\,
            sr => \N__52990\
        );

    \sDAC_mem_25_2_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50299\,
            lcout => \sDAC_mem_25Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47788\,
            ce => \N__41723\,
            sr => \N__52990\
        );

    \sDAC_mem_25_5_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47131\,
            lcout => \sDAC_mem_25Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47788\,
            ce => \N__41723\,
            sr => \N__52990\
        );

    \sDAC_mem_25_0_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51271\,
            lcout => \sDAC_mem_25Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47802\,
            ce => \N__41727\,
            sr => \N__52985\
        );

    \sDAC_mem_25_6_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48342\,
            lcout => \sDAC_mem_25Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47802\,
            ce => \N__41727\,
            sr => \N__52985\
        );

    \sDAC_mem_25_3_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49833\,
            lcout => \sDAC_mem_25Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47802\,
            ce => \N__41727\,
            sr => \N__52985\
        );

    \sDAC_mem_34_1_LC_17_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50500\,
            lcout => \sDAC_mem_34Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47789\,
            ce => \N__40088\,
            sr => \N__53138\
        );

    \sDAC_mem_34_3_LC_17_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49626\,
            lcout => \sDAC_mem_34Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47789\,
            ce => \N__40088\,
            sr => \N__53138\
        );

    \sDAC_mem_39_0_LC_17_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51083\,
            lcout => \sDAC_mem_39Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47773\,
            ce => \N__40140\,
            sr => \N__53133\
        );

    \sDAC_mem_39_1_LC_17_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50678\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_39Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47773\,
            ce => \N__40140\,
            sr => \N__53133\
        );

    \sDAC_mem_39_2_LC_17_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50255\,
            lcout => \sDAC_mem_39Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47773\,
            ce => \N__40140\,
            sr => \N__53133\
        );

    \sDAC_mem_39_3_LC_17_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49784\,
            lcout => \sDAC_mem_39Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47773\,
            ce => \N__40140\,
            sr => \N__53133\
        );

    \sDAC_mem_39_4_LC_17_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49357\,
            lcout => \sDAC_mem_39Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47773\,
            ce => \N__40140\,
            sr => \N__53133\
        );

    \sDAC_mem_39_5_LC_17_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46985\,
            lcout => \sDAC_mem_39Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47773\,
            ce => \N__40140\,
            sr => \N__53133\
        );

    \sDAC_mem_39_6_LC_17_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48210\,
            lcout => \sDAC_mem_39Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47773\,
            ce => \N__40140\,
            sr => \N__53133\
        );

    \sDAC_mem_39_7_LC_17_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48739\,
            lcout => \sDAC_mem_39Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47773\,
            ce => \N__40140\,
            sr => \N__53133\
        );

    \sAddress_RNI9IH12_0_3_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__40609\,
            in1 => \N__40407\,
            in2 => \N__44593\,
            in3 => \N__40633\,
            lcout => \sDAC_mem_40_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_13_3_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__40636\,
            in1 => \N__46250\,
            in2 => \N__40418\,
            in3 => \N__40610\,
            lcout => \sDAC_mem_37_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_12_3_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__40611\,
            in1 => \N__40412\,
            in2 => \N__44594\,
            in3 => \N__40635\,
            lcout => \sDAC_mem_39_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_11_3_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__40634\,
            in1 => \N__40612\,
            in2 => \N__40419\,
            in3 => \N__43255\,
            lcout => \sDAC_mem_35_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_3_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__43256\,
            in1 => \N__40406\,
            in2 => \N__40614\,
            in3 => \N__40637\,
            lcout => \sDAC_mem_36_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIVREN1_4_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46573\,
            in1 => \N__44649\,
            in2 => \N__44807\,
            in3 => \N__44750\,
            lcout => \N_288\,
            ltout => \N_288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_1_3_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__40608\,
            in1 => \N__46249\,
            in2 => \N__40422\,
            in3 => \N__40408\,
            lcout => \sDAC_mem_38_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_35_0_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51155\,
            lcout => \sDAC_mem_35Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47750\,
            ce => \N__40710\,
            sr => \N__53113\
        );

    \sDAC_mem_35_1_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50707\,
            lcout => \sDAC_mem_35Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47750\,
            ce => \N__40710\,
            sr => \N__53113\
        );

    \sDAC_mem_35_2_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50242\,
            lcout => \sDAC_mem_35Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47750\,
            ce => \N__40710\,
            sr => \N__53113\
        );

    \sDAC_mem_35_3_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49767\,
            lcout => \sDAC_mem_35Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47750\,
            ce => \N__40710\,
            sr => \N__53113\
        );

    \sDAC_mem_35_4_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49356\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_35Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47750\,
            ce => \N__40710\,
            sr => \N__53113\
        );

    \sDAC_mem_35_5_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46986\,
            lcout => \sDAC_mem_35Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47750\,
            ce => \N__40710\,
            sr => \N__53113\
        );

    \sDAC_mem_35_6_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48213\,
            lcout => \sDAC_mem_35Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47750\,
            ce => \N__40710\,
            sr => \N__53113\
        );

    \sDAC_mem_35_7_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48797\,
            lcout => \sDAC_mem_35Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47750\,
            ce => \N__40710\,
            sr => \N__53113\
        );

    \sDAC_mem_21_0_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51157\,
            lcout => \sDAC_mem_21Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47737\,
            ce => \N__40674\,
            sr => \N__53101\
        );

    \sDAC_mem_21_1_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50708\,
            lcout => \sDAC_mem_21Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47737\,
            ce => \N__40674\,
            sr => \N__53101\
        );

    \sDAC_mem_21_2_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50243\,
            lcout => \sDAC_mem_21Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47737\,
            ce => \N__40674\,
            sr => \N__53101\
        );

    \sDAC_mem_21_3_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49768\,
            lcout => \sDAC_mem_21Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47737\,
            ce => \N__40674\,
            sr => \N__53101\
        );

    \sDAC_mem_21_4_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49207\,
            lcout => \sDAC_mem_21Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47737\,
            ce => \N__40674\,
            sr => \N__53101\
        );

    \sDAC_mem_21_5_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46983\,
            lcout => \sDAC_mem_21Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47737\,
            ce => \N__40674\,
            sr => \N__53101\
        );

    \sDAC_mem_21_6_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48214\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_21Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47737\,
            ce => \N__40674\,
            sr => \N__53101\
        );

    \sDAC_mem_21_7_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48741\,
            lcout => \sDAC_mem_21Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47737\,
            ce => \N__40674\,
            sr => \N__53101\
        );

    \sDAC_data_RNO_13_6_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__41634\,
            in1 => \N__51812\,
            in2 => \N__43636\,
            in3 => \N__40830\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_6_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__40857\,
            in1 => \N__52120\,
            in2 => \N__40845\,
            in3 => \N__40842\,
            lcout => \sDAC_data_RNO_5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_6_3_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49769\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_6Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47727\,
            ce => \N__43085\,
            sr => \N__53087\
        );

    \sDAC_mem_6_4_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49312\,
            lcout => \sDAC_mem_6Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47727\,
            ce => \N__43085\,
            sr => \N__53087\
        );

    \sDAC_data_RNO_13_8_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__41889\,
            in1 => \N__51813\,
            in2 => \N__43637\,
            in3 => \N__40818\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_8_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__40806\,
            in1 => \N__52121\,
            in2 => \N__40794\,
            in3 => \N__40791\,
            lcout => \sDAC_data_RNO_5Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_8_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__40779\,
            in1 => \N__45870\,
            in2 => \N__40734\,
            in3 => \N__40767\,
            lcout => \sDAC_data_RNO_10Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_8_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__45868\,
            in1 => \N__45526\,
            in2 => \N__40758\,
            in3 => \N__40746\,
            lcout => \sDAC_data_2_32_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_8_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__45527\,
            in1 => \N__45869\,
            in2 => \N__40989\,
            in3 => \N__40977\,
            lcout => OPEN,
            ltout => \sDAC_data_2_14_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_8_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__45871\,
            in1 => \N__40968\,
            in2 => \N__40962\,
            in3 => \N__40959\,
            lcout => \sDAC_data_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_8_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101010101"
        )
    port map (
            in0 => \N__42639\,
            in1 => \N__40953\,
            in2 => \N__40947\,
            in3 => \N__42525\,
            lcout => OPEN,
            ltout => \sDAC_data_2_41_ns_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_8_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111000001110"
        )
    port map (
            in0 => \N__42526\,
            in1 => \N__42771\,
            in2 => \N__40929\,
            in3 => \N__40926\,
            lcout => OPEN,
            ltout => \sDAC_data_2_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_8_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47262\,
            in2 => \N__40920\,
            in3 => \N__42383\,
            lcout => \sDAC_dataZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53258\,
            ce => \N__42223\,
            sr => \N__53075\
        );

    \sDAC_mem_3_1_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50740\,
            lcout => \sDAC_mem_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47714\,
            ce => \N__42985\,
            sr => \N__53064\
        );

    \sDAC_data_RNO_28_4_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__52109\,
            in1 => \N__43628\,
            in2 => \N__40899\,
            in3 => \N__40884\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_4_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52107\,
            in1 => \N__40875\,
            in2 => \N__40866\,
            in3 => \N__40863\,
            lcout => \sDAC_data_RNO_15Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_6_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43629\,
            in1 => \N__44172\,
            in2 => \_gnd_net_\,
            in3 => \N__44304\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_6_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52110\,
            in2 => \N__41103\,
            in3 => \N__45192\,
            lcout => \sDAC_data_RNO_8Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_6_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52111\,
            in1 => \N__41820\,
            in2 => \N__43670\,
            in3 => \N__41100\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_6_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52108\,
            in1 => \N__43959\,
            in2 => \N__41088\,
            in3 => \N__47178\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_7Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_6_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101100010"
        )
    port map (
            in0 => \N__45873\,
            in1 => \N__41085\,
            in2 => \N__41073\,
            in3 => \N__41070\,
            lcout => \sDAC_data_RNO_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_4_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__41265\,
            in1 => \N__41943\,
            in2 => \N__45945\,
            in3 => \N__41049\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_10Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_4_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110011101"
        )
    port map (
            in0 => \N__42641\,
            in1 => \N__42531\,
            in2 => \N__41064\,
            in3 => \N__41577\,
            lcout => \sDAC_data_2_41_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_4_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__45938\,
            in1 => \N__45528\,
            in2 => \N__41676\,
            in3 => \N__41061\,
            lcout => \sDAC_data_2_32_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_4_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__45529\,
            in1 => \N__45942\,
            in2 => \N__41043\,
            in3 => \N__41031\,
            lcout => OPEN,
            ltout => \sDAC_data_2_14_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_4_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__45943\,
            in1 => \N__41019\,
            in2 => \N__41004\,
            in3 => \N__41001\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_4_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__42530\,
            in1 => \N__43299\,
            in2 => \N__41214\,
            in3 => \N__41211\,
            lcout => OPEN,
            ltout => \sDAC_data_2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_4_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46002\,
            in2 => \N__41205\,
            in3 => \N__42366\,
            lcout => \sDAC_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53269\,
            ce => \N__42224\,
            sr => \N__53054\
        );

    \sDAC_data_RNO_10_3_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__41190\,
            in1 => \N__41967\,
            in2 => \N__45909\,
            in3 => \N__41166\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_10Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_3_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__42522\,
            in1 => \N__42642\,
            in2 => \N__41178\,
            in3 => \N__41385\,
            lcout => \sDAC_data_2_41_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_3_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__45883\,
            in1 => \N__45457\,
            in2 => \N__44070\,
            in3 => \N__41175\,
            lcout => \sDAC_data_2_32_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_3_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__45458\,
            in1 => \N__45887\,
            in2 => \N__41160\,
            in3 => \N__41142\,
            lcout => OPEN,
            ltout => \sDAC_data_2_14_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_1_3_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__45888\,
            in1 => \N__41136\,
            in2 => \N__41121\,
            in3 => \N__41118\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_3_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__42523\,
            in1 => \N__43002\,
            in2 => \N__41112\,
            in3 => \N__41109\,
            lcout => OPEN,
            ltout => \sDAC_data_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_3_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__42377\,
            in1 => \N__46017\,
            in2 => \N__41373\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53271\,
            ce => \N__42226\,
            sr => \N__53044\
        );

    \sDAC_data_RNO_29_10_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41352\,
            in1 => \N__51993\,
            in2 => \_gnd_net_\,
            in3 => \N__41337\,
            lcout => \sDAC_data_RNO_29Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_30_6_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41316\,
            in1 => \N__51994\,
            in2 => \_gnd_net_\,
            in3 => \N__41304\,
            lcout => \sDAC_data_RNO_30Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_3_5_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__44430\,
            in1 => \N__46574\,
            in2 => \N__46251\,
            in3 => \N__46322\,
            lcout => \sDAC_mem_14_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_21_4_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52153\,
            in1 => \N__41295\,
            in2 => \_gnd_net_\,
            in3 => \N__41280\,
            lcout => \sDAC_data_RNO_21Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_27_1_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50761\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_27Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47728\,
            ce => \N__45245\,
            sr => \N__53025\
        );

    \sDAC_mem_27_2_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50174\,
            lcout => \sDAC_mem_27Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47728\,
            ce => \N__45245\,
            sr => \N__53025\
        );

    \sDAC_mem_27_3_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49794\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_27Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47728\,
            ce => \N__45245\,
            sr => \N__53025\
        );

    \sDAC_mem_27_4_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49231\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_27Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47728\,
            ce => \N__45245\,
            sr => \N__53025\
        );

    \sDAC_mem_27_5_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47081\,
            lcout => \sDAC_mem_27Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47728\,
            ce => \N__45245\,
            sr => \N__53025\
        );

    \sDAC_mem_27_6_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48331\,
            lcout => \sDAC_mem_27Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47728\,
            ce => \N__45245\,
            sr => \N__53025\
        );

    \sDAC_mem_27_7_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48841\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_27Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47728\,
            ce => \N__45245\,
            sr => \N__53025\
        );

    \sEEADC_freq_0_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51269\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEADC_freqZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47738\,
            ce => \N__44122\,
            sr => \_gnd_net_\
        );

    \sEEADC_freq_6_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48332\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEADC_freqZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47738\,
            ce => \N__44122\,
            sr => \_gnd_net_\
        );

    \sEEADC_freq_7_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48818\,
            lcout => \sEEADC_freqZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47738\,
            ce => \N__44122\,
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_24_3_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51771\,
            in1 => \N__41427\,
            in2 => \_gnd_net_\,
            in3 => \N__41415\,
            lcout => \sDAC_data_RNO_24Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_23_3_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52073\,
            in1 => \N__41409\,
            in2 => \_gnd_net_\,
            in3 => \N__41613\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_23Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_3_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__45879\,
            in1 => \N__41400\,
            in2 => \N__41394\,
            in3 => \N__41391\,
            lcout => \sDAC_data_RNO_11Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_28_0_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51272\,
            lcout => \sDAC_mem_28Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47751\,
            ce => \N__41777\,
            sr => \N__53014\
        );

    \sDAC_data_RNO_31_4_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51772\,
            in1 => \N__41607\,
            in2 => \_gnd_net_\,
            in3 => \N__41736\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_31Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_25_4_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__45881\,
            in1 => \N__45501\,
            in2 => \N__41595\,
            in3 => \N__41547\,
            lcout => OPEN,
            ltout => \sDAC_data_2_39_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_11_4_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__45880\,
            in1 => \N__41592\,
            in2 => \N__41586\,
            in3 => \N__41583\,
            lcout => \sDAC_data_RNO_11Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_32_4_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41568\,
            in1 => \N__51770\,
            in2 => \_gnd_net_\,
            in3 => \N__41556\,
            lcout => \sDAC_data_RNO_32Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_28_1_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50771\,
            lcout => \sDAC_mem_28Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47762\,
            ce => \N__41776\,
            sr => \N__53005\
        );

    \sDAC_mem_28_2_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50256\,
            lcout => \sDAC_mem_28Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47762\,
            ce => \N__41776\,
            sr => \N__53005\
        );

    \sDAC_mem_28_4_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49305\,
            lcout => \sDAC_mem_28Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47762\,
            ce => \N__41776\,
            sr => \N__53005\
        );

    \sDAC_mem_28_5_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47133\,
            lcout => \sDAC_mem_28Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47762\,
            ce => \N__41776\,
            sr => \N__53005\
        );

    \sDAC_mem_28_7_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48800\,
            lcout => \sDAC_mem_28Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47762\,
            ce => \N__41776\,
            sr => \N__53005\
        );

    \sAddress_RNI9IH12_1_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__46428\,
            in1 => \N__46132\,
            in2 => \_gnd_net_\,
            in3 => \N__43189\,
            lcout => \sDAC_mem_25_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_25_1_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50772\,
            lcout => \sDAC_mem_25Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47774\,
            ce => \N__41716\,
            sr => \N__52996\
        );

    \sDAC_data_RNO_29_4_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41694\,
            in1 => \N__51551\,
            in2 => \_gnd_net_\,
            in3 => \N__45219\,
            lcout => \sDAC_data_RNO_29Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_38_6_LC_18_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48227\,
            lcout => \sDAC_mem_38Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47763\,
            ce => \N__41867\,
            sr => \N__53139\
        );

    \sDAC_mem_38_0_LC_18_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51156\,
            lcout => \sDAC_mem_38Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47752\,
            ce => \N__41866\,
            sr => \N__53134\
        );

    \sDAC_mem_38_2_LC_18_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50078\,
            lcout => \sDAC_mem_38Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47752\,
            ce => \N__41866\,
            sr => \N__53134\
        );

    \sDAC_mem_38_3_LC_18_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49734\,
            lcout => \sDAC_mem_38Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47752\,
            ce => \N__41866\,
            sr => \N__53134\
        );

    \sDAC_mem_38_4_LC_18_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49362\,
            lcout => \sDAC_mem_38Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47752\,
            ce => \N__41866\,
            sr => \N__53134\
        );

    \sDAC_mem_38_5_LC_18_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47099\,
            lcout => \sDAC_mem_38Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47752\,
            ce => \N__41866\,
            sr => \N__53134\
        );

    \sDAC_mem_38_7_LC_18_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48742\,
            lcout => \sDAC_mem_38Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47752\,
            ce => \N__41866\,
            sr => \N__53134\
        );

    \sDAC_mem_40_0_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51158\,
            lcout => \sDAC_mem_40Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47739\,
            ce => \N__41985\,
            sr => \N__53128\
        );

    \sDAC_mem_40_1_LC_18_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50709\,
            lcout => \sDAC_mem_40Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47739\,
            ce => \N__41985\,
            sr => \N__53128\
        );

    \sDAC_mem_40_2_LC_18_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50079\,
            lcout => \sDAC_mem_40Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47739\,
            ce => \N__41985\,
            sr => \N__53128\
        );

    \sDAC_mem_40_3_LC_18_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49735\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_40Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47739\,
            ce => \N__41985\,
            sr => \N__53128\
        );

    \sDAC_mem_40_4_LC_18_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49363\,
            lcout => \sDAC_mem_40Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47739\,
            ce => \N__41985\,
            sr => \N__53128\
        );

    \sDAC_mem_40_5_LC_18_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47071\,
            lcout => \sDAC_mem_40Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47739\,
            ce => \N__41985\,
            sr => \N__53128\
        );

    \sDAC_mem_40_6_LC_18_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48228\,
            lcout => \sDAC_mem_40Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47739\,
            ce => \N__41985\,
            sr => \N__53128\
        );

    \sDAC_mem_40_7_LC_18_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48743\,
            lcout => \sDAC_mem_40Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47739\,
            ce => \N__41985\,
            sr => \N__53128\
        );

    \sDAC_data_RNO_20_3_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52003\,
            in1 => \N__41973\,
            in2 => \_gnd_net_\,
            in3 => \N__41955\,
            lcout => \sDAC_data_RNO_20Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_20_0_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51164\,
            lcout => \sDAC_mem_20Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47729\,
            ce => \N__44030\,
            sr => \N__53114\
        );

    \sDAC_data_RNO_20_4_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52004\,
            in1 => \N__41949\,
            in2 => \_gnd_net_\,
            in3 => \N__41931\,
            lcout => \sDAC_data_RNO_20Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_20_1_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50710\,
            lcout => \sDAC_mem_20Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47729\,
            ce => \N__44030\,
            sr => \N__53114\
        );

    \sDAC_data_RNO_20_5_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52005\,
            in1 => \N__41925\,
            in2 => \_gnd_net_\,
            in3 => \N__41910\,
            lcout => \sDAC_data_RNO_20Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_20_2_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50080\,
            lcout => \sDAC_mem_20Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47729\,
            ce => \N__44030\,
            sr => \N__53114\
        );

    \sDAC_data_RNO_20_6_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52006\,
            in1 => \N__41904\,
            in2 => \_gnd_net_\,
            in3 => \N__41895\,
            lcout => \sDAC_data_RNO_20Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_20_3_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49736\,
            lcout => \sDAC_mem_20Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47729\,
            ce => \N__44030\,
            sr => \N__53114\
        );

    \sDAC_data_RNO_26_6_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__43579\,
            in1 => \N__51804\,
            in2 => \N__42144\,
            in3 => \N__42114\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_6_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42159\,
            in2 => \N__42147\,
            in3 => \N__42120\,
            lcout => \sDAC_data_RNO_14Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_27_6_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__43577\,
            in1 => \N__51802\,
            in2 => \N__42143\,
            in3 => \N__42113\,
            lcout => \sDAC_data_RNO_27Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_1_3_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49824\,
            lcout => \sDAC_mem_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47719\,
            ce => \N__42039\,
            sr => \N__53102\
        );

    \sDAC_data_RNO_26_7_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__43578\,
            in1 => \N__51803\,
            in2 => \N__42078\,
            in3 => \N__42048\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_26Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_14_7_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42105\,
            in2 => \N__42096\,
            in3 => \N__42054\,
            lcout => \sDAC_data_RNO_14Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_27_7_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__43576\,
            in1 => \N__51801\,
            in2 => \N__42077\,
            in3 => \N__42047\,
            lcout => \sDAC_data_RNO_27Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_1_4_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49334\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47719\,
            ce => \N__42039\,
            sr => \N__53102\
        );

    \sDAC_data_RNO_1_6_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__42015\,
            in1 => \N__42009\,
            in2 => \N__45944\,
            in3 => \N__42708\,
            lcout => \sDAC_data_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_6_6_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__45932\,
            in1 => \N__45524\,
            in2 => \N__42816\,
            in3 => \N__42714\,
            lcout => \sDAC_data_2_14_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_22_6_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__45525\,
            in1 => \N__45933\,
            in2 => \N__42702\,
            in3 => \N__42681\,
            lcout => OPEN,
            ltout => \sDAC_data_2_32_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_10_6_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__45934\,
            in1 => \N__42669\,
            in2 => \N__42654\,
            in3 => \N__42651\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_10Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_3_6_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__42524\,
            in1 => \N__42640\,
            in2 => \N__42555\,
            in3 => \N__42552\,
            lcout => OPEN,
            ltout => \sDAC_data_2_41_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_0_6_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111000001110"
        )
    port map (
            in0 => \N__42527\,
            in1 => \N__42399\,
            in2 => \N__42393\,
            in3 => \N__42390\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_6_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__42384\,
            in1 => \N__45975\,
            in2 => \N__42255\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53264\,
            ce => \N__42221\,
            sr => \N__53088\
        );

    \sDAC_mem_3_3_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49818\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47708\,
            ce => \N__42992\,
            sr => \N__53076\
        );

    \sDAC_data_RNO_28_6_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__43543\,
            in1 => \N__52141\,
            in2 => \N__42186\,
            in3 => \N__42171\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_6_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52142\,
            in1 => \N__42837\,
            in2 => \N__42825\,
            in3 => \N__42822\,
            lcout => \sDAC_data_RNO_15Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_8_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__44376\,
            in1 => \_gnd_net_\,
            in2 => \N__43622\,
            in3 => \N__44277\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_8_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__52143\,
            in1 => \N__45165\,
            in2 => \N__42807\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_data_RNO_8Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_8_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52144\,
            in1 => \N__42804\,
            in2 => \N__43623\,
            in3 => \N__42795\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_8_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__46662\,
            in1 => \N__52145\,
            in2 => \N__42783\,
            in3 => \N__44244\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_7Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_8_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101100010"
        )
    port map (
            in0 => \N__45872\,
            in1 => \N__43896\,
            in2 => \N__42780\,
            in3 => \N__42777\,
            lcout => \sDAC_data_RNO_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_13_9_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52154\,
            in1 => \N__42765\,
            in2 => \N__43689\,
            in3 => \N__43095\,
            lcout => OPEN,
            ltout => \sDAC_data_2_13_bm_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_5_9_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52079\,
            in1 => \N__42756\,
            in2 => \N__42744\,
            in3 => \N__42741\,
            lcout => \sDAC_data_RNO_5Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_6_6_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48329\,
            lcout => \sDAC_mem_6Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47704\,
            ce => \N__43089\,
            sr => \N__53065\
        );

    \sDAC_data_RNO_16_3_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__52078\,
            in1 => \N__43041\,
            in2 => \N__43688\,
            in3 => \N__43032\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_3_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52155\,
            in1 => \N__43998\,
            in2 => \N__43017\,
            in3 => \N__47217\,
            lcout => \sDAC_data_RNO_7Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_3_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43682\,
            in1 => \N__44208\,
            in2 => \_gnd_net_\,
            in3 => \N__44340\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_3_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52080\,
            in2 => \N__43014\,
            in3 => \N__45012\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_8Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_3_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001010100"
        )
    port map (
            in0 => \N__45099\,
            in1 => \N__45931\,
            in2 => \N__43011\,
            in3 => \N__43008\,
            lcout => \sDAC_data_RNO_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_3_7_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48778\,
            lcout => \sDAC_mem_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47709\,
            ce => \N__42996\,
            sr => \N__53055\
        );

    \sDAC_data_RNO_28_10_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__43674\,
            in1 => \N__52065\,
            in2 => \N__42906\,
            in3 => \N__42885\,
            lcout => OPEN,
            ltout => \sDAC_data_2_6_bm_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_15_10_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__52067\,
            in1 => \N__42870\,
            in2 => \N__42858\,
            in3 => \N__42855\,
            lcout => \sDAC_data_RNO_15Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_16_4_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__43716\,
            in1 => \N__52066\,
            in2 => \N__43687\,
            in3 => \N__43707\,
            lcout => OPEN,
            ltout => \sDAC_data_2_20_am_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_7_4_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__43986\,
            in1 => \N__47205\,
            in2 => \N__43692\,
            in3 => \N__52139\,
            lcout => \sDAC_data_RNO_7Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_17_4_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43678\,
            in1 => \N__44196\,
            in2 => \_gnd_net_\,
            in3 => \N__44331\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_17Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_8_4_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52140\,
            in2 => \N__43311\,
            in3 => \N__45006\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_8Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_2_4_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001010100"
        )
    port map (
            in0 => \N__45300\,
            in1 => \N__45889\,
            in2 => \N__43308\,
            in3 => \N__43305\,
            lcout => \sDAC_data_RNO_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI5B15_2_1_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44896\,
            in2 => \_gnd_net_\,
            in3 => \N__44831\,
            lcout => \N_284\,
            ltout => \N_284_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_4_5_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__46321\,
            in1 => \N__44445\,
            in2 => \N__43290\,
            in3 => \N__46569\,
            lcout => \sDAC_mem_12_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_8_5_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__43226\,
            in1 => \N__46119\,
            in2 => \N__46575\,
            in3 => \N__46320\,
            lcout => \sDAC_mem_11_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_3_1_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__46118\,
            in1 => \N__43225\,
            in2 => \_gnd_net_\,
            in3 => \N__43191\,
            lcout => \sDAC_mem_27_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_1_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50672\,
            in2 => \_gnd_net_\,
            in3 => \N__43868\,
            lcout => \sAddressZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47715\,
            ce => \N__43779\,
            sr => \N__53045\
        );

    \sAddress_RNI5B15_1_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44897\,
            in2 => \_gnd_net_\,
            in3 => \N__44832\,
            lcout => \N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_2_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50077\,
            in2 => \_gnd_net_\,
            in3 => \N__43869\,
            lcout => \sAddressZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47715\,
            ce => \N__43779\,
            sr => \N__53045\
        );

    \sDAC_mem_14_0_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51268\,
            lcout => \sDAC_mem_14Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47720\,
            ce => \N__43935\,
            sr => \N__53035\
        );

    \sDAC_mem_14_1_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50762\,
            lcout => \sDAC_mem_14Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47720\,
            ce => \N__43935\,
            sr => \N__53035\
        );

    \sDAC_mem_14_2_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50090\,
            lcout => \sDAC_mem_14Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47720\,
            ce => \N__43935\,
            sr => \N__53035\
        );

    \sDAC_mem_14_3_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49842\,
            lcout => \sDAC_mem_14Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47720\,
            ce => \N__43935\,
            sr => \N__53035\
        );

    \sDAC_mem_14_4_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49308\,
            lcout => \sDAC_mem_14Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47720\,
            ce => \N__43935\,
            sr => \N__53035\
        );

    \sDAC_mem_14_5_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47132\,
            lcout => \sDAC_mem_14Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47720\,
            ce => \N__43935\,
            sr => \N__53035\
        );

    \sDAC_mem_14_6_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48340\,
            lcout => \sDAC_mem_14Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47720\,
            ce => \N__43935\,
            sr => \N__53035\
        );

    \sDAC_mem_14_7_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48786\,
            lcout => \sDAC_mem_14Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47720\,
            ce => \N__43935\,
            sr => \N__53035\
        );

    \sDAC_data_RNO_19_7_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51973\,
            in1 => \N__45060\,
            in2 => \_gnd_net_\,
            in3 => \N__43929\,
            lcout => \sDAC_data_RNO_19Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_7_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51983\,
            in1 => \N__48885\,
            in2 => \_gnd_net_\,
            in3 => \N__43887\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_7_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__45890\,
            in1 => \N__45492\,
            in2 => \N__43923\,
            in3 => \N__43920\,
            lcout => \sDAC_data_2_24_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_8_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51984\,
            in1 => \N__45225\,
            in2 => \_gnd_net_\,
            in3 => \N__44148\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_8_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__45891\,
            in1 => \N__45493\,
            in2 => \N__43899\,
            in3 => \N__43875\,
            lcout => \sDAC_data_2_24_ns_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_12_4_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49166\,
            lcout => \sDAC_mem_12Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47730\,
            ce => \N__47376\,
            sr => \N__53026\
        );

    \sDAC_data_RNO_19_8_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51974\,
            in1 => \N__45048\,
            in2 => \_gnd_net_\,
            in3 => \N__43881\,
            lcout => \sDAC_data_RNO_19Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_12_5_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47147\,
            lcout => \sDAC_mem_12Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47730\,
            ce => \N__47376\,
            sr => \N__53026\
        );

    \sEEADC_freq_1_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50673\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEADC_freqZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47740\,
            ce => \N__44126\,
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_29_3_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44094\,
            in1 => \N__51890\,
            in2 => \_gnd_net_\,
            in3 => \N__44082\,
            lcout => \sDAC_data_RNO_29Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_16_3_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49845\,
            lcout => \sDAC_mem_16Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47775\,
            ce => \N__46631\,
            sr => \N__52997\
        );

    \sDAC_mem_20_7_LC_19_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48744\,
            lcout => \sDAC_mem_20Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47731\,
            ce => \N__44031\,
            sr => \N__53135\
        );

    \sDAC_mem_41_0_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51239\,
            lcout => \sDAC_mem_41Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47721\,
            ce => \N__46263\,
            sr => \N__53129\
        );

    \sDAC_mem_41_1_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50580\,
            lcout => \sDAC_mem_41Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47721\,
            ce => \N__46263\,
            sr => \N__53129\
        );

    \sDAC_mem_41_2_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50230\,
            lcout => \sDAC_mem_41Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47721\,
            ce => \N__46263\,
            sr => \N__53129\
        );

    \sDAC_mem_41_3_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49737\,
            lcout => \sDAC_mem_41Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47721\,
            ce => \N__46263\,
            sr => \N__53129\
        );

    \sDAC_mem_41_4_LC_19_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49281\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_41Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47721\,
            ce => \N__46263\,
            sr => \N__53129\
        );

    \sDAC_mem_41_5_LC_19_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46984\,
            lcout => \sDAC_mem_41Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47721\,
            ce => \N__46263\,
            sr => \N__53129\
        );

    \sDAC_mem_41_6_LC_19_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48229\,
            lcout => \sDAC_mem_41Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47721\,
            ce => \N__46263\,
            sr => \N__53129\
        );

    \sDAC_mem_41_7_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48745\,
            lcout => \sDAC_mem_41Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47721\,
            ce => \N__46263\,
            sr => \N__53129\
        );

    \sDAC_mem_42_0_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51168\,
            lcout => \sDAC_mem_42Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47716\,
            ce => \N__44976\,
            sr => \N__53115\
        );

    \sDAC_mem_42_1_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50581\,
            lcout => \sDAC_mem_42Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47716\,
            ce => \N__44976\,
            sr => \N__53115\
        );

    \sDAC_mem_42_2_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50291\,
            lcout => \sDAC_mem_42Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47716\,
            ce => \N__44976\,
            sr => \N__53115\
        );

    \sDAC_mem_42_3_LC_19_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49825\,
            lcout => \sDAC_mem_42Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47716\,
            ce => \N__44976\,
            sr => \N__53115\
        );

    \sDAC_mem_42_4_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49335\,
            lcout => \sDAC_mem_42Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47716\,
            ce => \N__44976\,
            sr => \N__53115\
        );

    \sDAC_mem_42_5_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47137\,
            lcout => \sDAC_mem_42Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47716\,
            ce => \N__44976\,
            sr => \N__53115\
        );

    \sDAC_mem_42_6_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48278\,
            lcout => \sDAC_mem_42Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47716\,
            ce => \N__44976\,
            sr => \N__53115\
        );

    \sDAC_mem_42_7_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48833\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_42Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47716\,
            ce => \N__44976\,
            sr => \N__53115\
        );

    \sDAC_mem_10_0_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51240\,
            lcout => \sDAC_mem_10Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47710\,
            ce => \N__44993\,
            sr => \N__53103\
        );

    \sDAC_mem_10_1_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50582\,
            lcout => \sDAC_mem_10Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47710\,
            ce => \N__44993\,
            sr => \N__53103\
        );

    \sDAC_mem_10_2_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50286\,
            lcout => \sDAC_mem_10Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47710\,
            ce => \N__44993\,
            sr => \N__53103\
        );

    \sDAC_mem_10_3_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49811\,
            lcout => \sDAC_mem_10Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47710\,
            ce => \N__44993\,
            sr => \N__53103\
        );

    \sDAC_mem_10_4_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49336\,
            lcout => \sDAC_mem_10Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47710\,
            ce => \N__44993\,
            sr => \N__53103\
        );

    \sDAC_mem_10_5_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47138\,
            lcout => \sDAC_mem_10Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47710\,
            ce => \N__44993\,
            sr => \N__53103\
        );

    \sDAC_mem_10_6_LC_19_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48279\,
            lcout => \sDAC_mem_10Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47710\,
            ce => \N__44993\,
            sr => \N__53103\
        );

    \sAddress_RNI9IH12_10_5_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__46294\,
            in1 => \N__46413\,
            in2 => \N__44470\,
            in3 => \N__46563\,
            lcout => \sDAC_mem_10_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_6_5_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__46566\,
            in1 => \N__46123\,
            in2 => \N__44554\,
            in3 => \N__46292\,
            lcout => \sDAC_mem_15_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_5_5_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__46295\,
            in1 => \N__46414\,
            in2 => \N__44471\,
            in3 => \N__46564\,
            lcout => \sDAC_mem_42_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI5B15_0_1_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44931\,
            in2 => \_gnd_net_\,
            in3 => \N__44855\,
            lcout => \N_286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNIP2UK1_4_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__44778\,
            in1 => \N__44722\,
            in2 => \_gnd_net_\,
            in3 => \N__44636\,
            lcout => \N_278\,
            ltout => \N_278_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_2_5_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__46565\,
            in1 => \N__44539\,
            in2 => \N__44481\,
            in3 => \N__44459\,
            lcout => \sDAC_mem_16_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_9_5_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__46296\,
            in1 => \N__46412\,
            in2 => \N__46133\,
            in3 => \N__46568\,
            lcout => \sDAC_mem_9_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_7_5_LC_19_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__46567\,
            in1 => \N__46124\,
            in2 => \N__46247\,
            in3 => \N__46293\,
            lcout => \sDAC_mem_13_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_15_0_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51241\,
            lcout => \sDAC_mem_15Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47702\,
            ce => \N__45024\,
            sr => \N__53077\
        );

    \sDAC_mem_15_1_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50583\,
            lcout => \sDAC_mem_15Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47702\,
            ce => \N__45024\,
            sr => \N__53077\
        );

    \sDAC_mem_15_2_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50287\,
            lcout => \sDAC_mem_15Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47702\,
            ce => \N__45024\,
            sr => \N__53077\
        );

    \sDAC_mem_15_3_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49819\,
            lcout => \sDAC_mem_15Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47702\,
            ce => \N__45024\,
            sr => \N__53077\
        );

    \sDAC_mem_15_4_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49359\,
            lcout => \sDAC_mem_15Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47702\,
            ce => \N__45024\,
            sr => \N__53077\
        );

    \sDAC_mem_15_5_LC_19_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47150\,
            lcout => \sDAC_mem_15Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47702\,
            ce => \N__45024\,
            sr => \N__53077\
        );

    \sDAC_mem_15_6_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48330\,
            lcout => \sDAC_mem_15Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47702\,
            ce => \N__45024\,
            sr => \N__53077\
        );

    \sDAC_mem_15_7_LC_19_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48812\,
            lcout => \sDAC_mem_15Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47702\,
            ce => \N__45024\,
            sr => \N__53077\
        );

    \sDAC_mem_11_0_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51242\,
            lcout => \sDAC_mem_11Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47705\,
            ce => \N__45129\,
            sr => \N__53066\
        );

    \sDAC_mem_11_1_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50584\,
            lcout => \sDAC_mem_11Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47705\,
            ce => \N__45129\,
            sr => \N__53066\
        );

    \sDAC_mem_11_2_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50307\,
            lcout => \sDAC_mem_11Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47705\,
            ce => \N__45129\,
            sr => \N__53066\
        );

    \sDAC_mem_11_3_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49841\,
            lcout => \sDAC_mem_11Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47705\,
            ce => \N__45129\,
            sr => \N__53066\
        );

    \sDAC_mem_11_4_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49322\,
            lcout => \sDAC_mem_11Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47705\,
            ce => \N__45129\,
            sr => \N__53066\
        );

    \sDAC_mem_11_5_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47151\,
            lcout => \sDAC_mem_11Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47705\,
            ce => \N__45129\,
            sr => \N__53066\
        );

    \sDAC_mem_11_6_LC_19_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48325\,
            lcout => \sDAC_mem_11Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47705\,
            ce => \N__45129\,
            sr => \N__53066\
        );

    \sDAC_mem_11_7_LC_19_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48779\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_11Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47705\,
            ce => \N__45129\,
            sr => \N__53066\
        );

    \sDAC_data_RNO_19_3_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52146\,
            in1 => \N__45123\,
            in2 => \_gnd_net_\,
            in3 => \N__45114\,
            lcout => \sDAC_data_RNO_19Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_3_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52148\,
            in1 => \N__50778\,
            in2 => \_gnd_net_\,
            in3 => \N__45294\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_3_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__45910\,
            in1 => \N__45494\,
            in2 => \N__45108\,
            in3 => \N__45105\,
            lcout => \sDAC_data_2_24_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_4_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52149\,
            in1 => \N__50316\,
            in2 => \_gnd_net_\,
            in3 => \N__45267\,
            lcout => OPEN,
            ltout => \sDAC_data_RNO_18Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_9_4_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__45911\,
            in1 => \N__45495\,
            in2 => \N__45303\,
            in3 => \N__45273\,
            lcout => \sDAC_data_2_24_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_12_0_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51270\,
            lcout => \sDAC_mem_12Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47711\,
            ce => \N__47375\,
            sr => \N__53056\
        );

    \sDAC_data_RNO_19_4_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52147\,
            in1 => \N__45288\,
            in2 => \_gnd_net_\,
            in3 => \N__45279\,
            lcout => \sDAC_data_RNO_19Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_12_1_LC_19_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50585\,
            lcout => \sDAC_mem_12Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47711\,
            ce => \N__47375\,
            sr => \N__53056\
        );

    \sDAC_mem_27_0_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51081\,
            lcout => \sDAC_mem_27Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47717\,
            ce => \N__45246\,
            sr => \N__53046\
        );

    \sDAC_mem_13_6_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48232\,
            lcout => \sDAC_mem_13Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47722\,
            ce => \N__48867\,
            sr => \N__53036\
        );

    \sDAC_mem_13_5_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47148\,
            lcout => \sDAC_mem_13Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47722\,
            ce => \N__48867\,
            sr => \N__53036\
        );

    \sDAC_mem_16_1_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50674\,
            lcout => \sDAC_mem_16Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47753\,
            ce => \N__46630\,
            sr => \N__53015\
        );

    \sEEDAC_7_LC_20_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48729\,
            lcout => \sEEDACZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47732\,
            ce => \N__47238\,
            sr => \_gnd_net_\
        );

    \sAddress_RNI9IH12_1_5_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__46559\,
            in1 => \N__46134\,
            in2 => \N__46445\,
            in3 => \N__46319\,
            lcout => \sDAC_mem_41_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_rpi_ibuf_RNIRGF52_0_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__46248\,
            in1 => \N__46128\,
            in2 => \_gnd_net_\,
            in3 => \N__46043\,
            lcout => \sEEDAC_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sEEDAC_0_LC_20_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51181\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEDACZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47712\,
            ce => \N__47234\,
            sr => \_gnd_net_\
        );

    \sEEDAC_1_LC_20_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50725\,
            lcout => \sEEDACZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47712\,
            ce => \N__47234\,
            sr => \_gnd_net_\
        );

    \sEEDAC_2_LC_20_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50292\,
            lcout => \sEEDACZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47712\,
            ce => \N__47234\,
            sr => \_gnd_net_\
        );

    \sEEDAC_3_LC_20_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49826\,
            lcout => \sEEDACZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47712\,
            ce => \N__47234\,
            sr => \_gnd_net_\
        );

    \sEEDAC_4_LC_20_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49343\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sEEDACZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47712\,
            ce => \N__47234\,
            sr => \_gnd_net_\
        );

    \sEEDAC_5_LC_20_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47139\,
            lcout => \sEEDACZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47712\,
            ce => \N__47234\,
            sr => \_gnd_net_\
        );

    \sEEDAC_6_LC_20_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48280\,
            lcout => \sEEDACZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47712\,
            ce => \N__47234\,
            sr => \_gnd_net_\
        );

    \sDAC_mem_9_0_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50981\,
            lcout => \sDAC_mem_9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47706\,
            ce => \N__47325\,
            sr => \N__53116\
        );

    \sDAC_mem_9_1_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50753\,
            lcout => \sDAC_mem_9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47706\,
            ce => \N__47325\,
            sr => \N__53116\
        );

    \sDAC_mem_9_2_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50308\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_9Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47706\,
            ce => \N__47325\,
            sr => \N__53116\
        );

    \sDAC_mem_9_3_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49843\,
            lcout => \sDAC_mem_9Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47706\,
            ce => \N__47325\,
            sr => \N__53116\
        );

    \sDAC_mem_9_4_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49344\,
            lcout => \sDAC_mem_9Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47706\,
            ce => \N__47325\,
            sr => \N__53116\
        );

    \sDAC_mem_9_5_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47140\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_9Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47706\,
            ce => \N__47325\,
            sr => \N__53116\
        );

    \sDAC_mem_9_6_LC_20_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48281\,
            lcout => \sDAC_mem_9Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47706\,
            ce => \N__47325\,
            sr => \N__53116\
        );

    \sDAC_mem_9_7_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48718\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_9Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47706\,
            ce => \N__47325\,
            sr => \N__53116\
        );

    \sCounterDAC_6_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011001100110"
        )
    port map (
            in0 => \N__52176\,
            in1 => \N__52444\,
            in2 => \N__52253\,
            in3 => \N__53449\,
            lcout => \sCounterDACZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53274\,
            ce => 'H',
            sr => \N__53104\
        );

    \sCounterDAC_RNI7A77_1_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__52547\,
            in1 => \N__53357\,
            in2 => \N__53414\,
            in3 => \N__52524\,
            lcout => \N_14_3\,
            ltout => \N_14_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_spi_start_RNO_0_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__47286\,
            in1 => \N__52548\,
            in2 => \N__47313\,
            in3 => \N__52232\,
            lcout => OPEN,
            ltout => \N_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_spi_start_LC_20_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__47300\,
            in1 => \N__47280\,
            in2 => \N__47310\,
            in3 => \N__53337\,
            lcout => \sDAC_spi_startZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53274\,
            ce => 'H',
            sr => \N__53104\
        );

    \sCounterDAC_RNIPQJ3_3_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__53335\,
            in1 => \N__52199\,
            in2 => \_gnd_net_\,
            in3 => \N__52233\,
            lcout => \N_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_spi_start_RNO_2_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__52200\,
            in1 => \N__52520\,
            in2 => \_gnd_net_\,
            in3 => \N__53336\,
            lcout => un1_scounterdac8_i_a2_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_spi_start_RNO_1_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__53410\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53451\,
            lcout => un1_scounterdac8_i_a2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_18_10_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52077\,
            in1 => \N__48873\,
            in2 => \_gnd_net_\,
            in3 => \N__48351\,
            lcout => \sDAC_data_RNO_18Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_data_RNO_19_10_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52076\,
            in1 => \N__51306\,
            in2 => \_gnd_net_\,
            in3 => \N__51300\,
            lcout => \sDAC_data_RNO_19Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sDAC_mem_13_0_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50982\,
            lcout => \sDAC_mem_13Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47703\,
            ce => \N__48866\,
            sr => \N__53078\
        );

    \sDAC_mem_13_1_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50576\,
            lcout => \sDAC_mem_13Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47703\,
            ce => \N__48866\,
            sr => \N__53078\
        );

    \sDAC_mem_13_2_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_13Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47703\,
            ce => \N__48866\,
            sr => \N__53078\
        );

    \sDAC_mem_13_3_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49844\,
            lcout => \sDAC_mem_13Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47703\,
            ce => \N__48866\,
            sr => \N__53078\
        );

    \sDAC_mem_13_4_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49355\,
            lcout => \sDAC_mem_13Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47703\,
            ce => \N__48866\,
            sr => \N__53078\
        );

    \sDAC_mem_13_7_LC_20_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48719\,
            lcout => \sDAC_mem_13Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47703\,
            ce => \N__48866\,
            sr => \N__53078\
        );

    \sDAC_mem_12_7_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48728\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sDAC_mem_12Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47707\,
            ce => \N__47377\,
            sr => \N__53067\
        );

    \sDAC_mem_12_6_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48341\,
            lcout => \sDAC_mem_12Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47723\,
            ce => \N__47391\,
            sr => \N__53037\
        );

    \sCounterDAC_8_LC_22_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010100101010"
        )
    port map (
            in0 => \N__53298\,
            in1 => \N__53450\,
            in2 => \N__52260\,
            in3 => \N__53322\,
            lcout => \sCounterDACZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53275\,
            ce => 'H',
            sr => \N__53140\
        );

    \un2_scounterdac_cry_1_c_LC_22_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52512\,
            in2 => \N__53395\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_22_10_0_\,
            carryout => un2_scounterdac_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_2_LC_22_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52476\,
            in2 => \_gnd_net_\,
            in3 => \N__52236\,
            lcout => \sCounterDACZ0Z_2\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_1,
            carryout => un2_scounterdac_cry_2,
            clk => \N__53277\,
            ce => 'H',
            sr => \N__53130\
        );

    \sCounterDAC_3_LC_22_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52225\,
            in2 => \_gnd_net_\,
            in3 => \N__52206\,
            lcout => \sCounterDACZ0Z_3\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_2,
            carryout => un2_scounterdac_cry_3,
            clk => \N__53277\,
            ce => 'H',
            sr => \N__53130\
        );

    \sCounterDAC_4_LC_22_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52541\,
            in2 => \_gnd_net_\,
            in3 => \N__52203\,
            lcout => \sCounterDACZ0Z_4\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_3,
            carryout => un2_scounterdac_cry_4,
            clk => \N__53277\,
            ce => 'H',
            sr => \N__53130\
        );

    \sCounterDAC_5_LC_22_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52193\,
            in2 => \_gnd_net_\,
            in3 => \N__52179\,
            lcout => \sCounterDACZ0Z_5\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_4,
            carryout => un2_scounterdac_cry_5,
            clk => \N__53277\,
            ce => 'H',
            sr => \N__53130\
        );

    \un2_scounterdac_cry_5_THRU_LUT4_0_LC_22_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__52449\,
            in3 => \N__52167\,
            lcout => \un2_scounterdac_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_5,
            carryout => un2_scounterdac_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_7_LC_22_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52488\,
            in2 => \_gnd_net_\,
            in3 => \N__52164\,
            lcout => \sCounterDACZ0Z_7\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_6,
            carryout => un2_scounterdac_cry_7,
            clk => \N__53277\,
            ce => 'H',
            sr => \N__53130\
        );

    \un2_scounterdac_cry_7_THRU_LUT4_0_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53331\,
            in2 => \_gnd_net_\,
            in3 => \N__53289\,
            lcout => \un2_scounterdac_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => un2_scounterdac_cry_7,
            carryout => un2_scounterdac_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_9_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52463\,
            in2 => \_gnd_net_\,
            in3 => \N__53286\,
            lcout => \sCounterDACZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53279\,
            ce => 'H',
            sr => \N__53117\
        );

    \sCounterDAC_0_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53405\,
            lcout => \sCounterDACZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53279\,
            ce => 'H',
            sr => \N__53117\
        );

    \sCounterDAC_1_LC_22_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53406\,
            in2 => \_gnd_net_\,
            in3 => \N__52519\,
            lcout => \sCounterDACZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__53279\,
            ce => 'H',
            sr => \N__53117\
        );

    \spi_slave_inst.spi_mosi_flash_LC_23_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52304\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52596\,
            lcout => spi_mosi_flash_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_RNIB1D2_1_LC_23_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52540\,
            in2 => \_gnd_net_\,
            in3 => \N__52511\,
            lcout => op_eq_scounterdac10_0_a2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_RNI4HQ4_9_LC_23_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__52487\,
            in1 => \N__52475\,
            in2 => \N__52464\,
            in3 => \N__52445\,
            lcout => \N_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.spi_cs_flash_LC_24_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52296\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52414\,
            lcout => spi_cs_flash_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \spi_slave_inst.spi_sclk_flash_LC_24_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52347\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52297\,
            lcout => spi_sclk_flash_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sCounterDAC_RNIBR1C_0_LC_24_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__53457\,
            in1 => \N__53436\,
            in2 => \N__53415\,
            in3 => \N__53364\,
            lcout => op_eq_scounterdac10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
