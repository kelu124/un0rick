pll248M2_inst: pll248M2
port map(
          REFERENCECLK => ,
          PLLOUTCOREA => ,
          PLLOUTCOREB => ,
          PLLOUTGLOBALA => ,
          PLLOUTGLOBALB => ,
          RESET => 
        );
