// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 13 2018 07:24:18

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MATTY_MAIN_VHDL" view "INTERFACE"

module MATTY_MAIN_VHDL (
    RAM_DATA,
    RAM_ADD,
    spi_sclk_ft,
    button_trig,
    ADC9,
    spi_cs_ft,
    poff,
    RAM_nOE,
    ADC0,
    spi_mosi_flash,
    spi_miso_flash,
    trig_ft,
    spi_miso_rpi,
    RAM_nWE,
    DAC_cs,
    ADC6,
    spi_select,
    clk,
    ADC4,
    trig_rpi,
    top_tour2,
    spi_cs_rpi,
    DAC_sclk,
    ADC_clk,
    ADC3,
    trig_ext,
    spi_mosi_rpi,
    spi_mosi_ft,
    cs_rpi2flash,
    spi_cs_flash,
    pon,
    RAM_nCE,
    LED3,
    ADC1,
    reset_rpi,
    RAM_nLB,
    LED_MODE,
    ADC8,
    spi_sclk_rpi,
    ADC7,
    top_tour1,
    spi_miso_ft,
    button_mode,
    DAC_mosi,
    ADC5,
    reset_ft,
    LED_ACQ,
    spi_sclk_flash,
    reset_alim,
    RAM_nUB,
    ADC2);

    inout [15:0] RAM_DATA;
    output [18:0] RAM_ADD;
    input spi_sclk_ft;
    input button_trig;
    input ADC9;
    input spi_cs_ft;
    output poff;
    output RAM_nOE;
    input ADC0;
    output spi_mosi_flash;
    input spi_miso_flash;
    input trig_ft;
    output spi_miso_rpi;
    output RAM_nWE;
    output DAC_cs;
    input ADC6;
    input spi_select;
    input clk;
    input ADC4;
    input trig_rpi;
    input top_tour2;
    input spi_cs_rpi;
    output DAC_sclk;
    output ADC_clk;
    input ADC3;
    input trig_ext;
    input spi_mosi_rpi;
    input spi_mosi_ft;
    input cs_rpi2flash;
    output spi_cs_flash;
    output pon;
    output RAM_nCE;
    output LED3;
    input ADC1;
    input reset_rpi;
    output RAM_nLB;
    output LED_MODE;
    input ADC8;
    input spi_sclk_rpi;
    input ADC7;
    input top_tour1;
    output spi_miso_ft;
    input button_mode;
    output DAC_mosi;
    input ADC5;
    input reset_ft;
    output LED_ACQ;
    output spi_sclk_flash;
    input reset_alim;
    output RAM_nUB;
    input ADC2;

    wire N__54196;
    wire N__54195;
    wire N__54194;
    wire N__54187;
    wire N__54186;
    wire N__54185;
    wire N__54178;
    wire N__54177;
    wire N__54176;
    wire N__54169;
    wire N__54168;
    wire N__54167;
    wire N__54160;
    wire N__54159;
    wire N__54158;
    wire N__54151;
    wire N__54150;
    wire N__54149;
    wire N__54142;
    wire N__54141;
    wire N__54140;
    wire N__54133;
    wire N__54132;
    wire N__54131;
    wire N__54124;
    wire N__54123;
    wire N__54122;
    wire N__54115;
    wire N__54114;
    wire N__54113;
    wire N__54106;
    wire N__54105;
    wire N__54104;
    wire N__54097;
    wire N__54096;
    wire N__54095;
    wire N__54088;
    wire N__54087;
    wire N__54086;
    wire N__54079;
    wire N__54078;
    wire N__54077;
    wire N__54070;
    wire N__54069;
    wire N__54068;
    wire N__54061;
    wire N__54060;
    wire N__54059;
    wire N__54052;
    wire N__54051;
    wire N__54050;
    wire N__54043;
    wire N__54042;
    wire N__54041;
    wire N__54034;
    wire N__54033;
    wire N__54032;
    wire N__54025;
    wire N__54024;
    wire N__54023;
    wire N__54016;
    wire N__54015;
    wire N__54014;
    wire N__54007;
    wire N__54006;
    wire N__54005;
    wire N__53998;
    wire N__53997;
    wire N__53996;
    wire N__53989;
    wire N__53988;
    wire N__53987;
    wire N__53980;
    wire N__53979;
    wire N__53978;
    wire N__53971;
    wire N__53970;
    wire N__53969;
    wire N__53962;
    wire N__53961;
    wire N__53960;
    wire N__53953;
    wire N__53952;
    wire N__53951;
    wire N__53944;
    wire N__53943;
    wire N__53942;
    wire N__53935;
    wire N__53934;
    wire N__53933;
    wire N__53926;
    wire N__53925;
    wire N__53924;
    wire N__53917;
    wire N__53916;
    wire N__53915;
    wire N__53908;
    wire N__53907;
    wire N__53906;
    wire N__53899;
    wire N__53898;
    wire N__53897;
    wire N__53890;
    wire N__53889;
    wire N__53888;
    wire N__53881;
    wire N__53880;
    wire N__53879;
    wire N__53872;
    wire N__53871;
    wire N__53870;
    wire N__53863;
    wire N__53862;
    wire N__53861;
    wire N__53854;
    wire N__53853;
    wire N__53852;
    wire N__53845;
    wire N__53844;
    wire N__53843;
    wire N__53836;
    wire N__53835;
    wire N__53834;
    wire N__53827;
    wire N__53826;
    wire N__53825;
    wire N__53818;
    wire N__53817;
    wire N__53816;
    wire N__53809;
    wire N__53808;
    wire N__53807;
    wire N__53800;
    wire N__53799;
    wire N__53798;
    wire N__53791;
    wire N__53790;
    wire N__53789;
    wire N__53782;
    wire N__53781;
    wire N__53780;
    wire N__53773;
    wire N__53772;
    wire N__53771;
    wire N__53764;
    wire N__53763;
    wire N__53762;
    wire N__53755;
    wire N__53754;
    wire N__53753;
    wire N__53746;
    wire N__53745;
    wire N__53744;
    wire N__53737;
    wire N__53736;
    wire N__53735;
    wire N__53728;
    wire N__53727;
    wire N__53726;
    wire N__53719;
    wire N__53718;
    wire N__53717;
    wire N__53710;
    wire N__53709;
    wire N__53708;
    wire N__53701;
    wire N__53700;
    wire N__53699;
    wire N__53692;
    wire N__53691;
    wire N__53690;
    wire N__53683;
    wire N__53682;
    wire N__53681;
    wire N__53674;
    wire N__53673;
    wire N__53672;
    wire N__53665;
    wire N__53664;
    wire N__53663;
    wire N__53656;
    wire N__53655;
    wire N__53654;
    wire N__53647;
    wire N__53646;
    wire N__53645;
    wire N__53638;
    wire N__53637;
    wire N__53636;
    wire N__53629;
    wire N__53628;
    wire N__53627;
    wire N__53620;
    wire N__53619;
    wire N__53618;
    wire N__53611;
    wire N__53610;
    wire N__53609;
    wire N__53602;
    wire N__53601;
    wire N__53600;
    wire N__53593;
    wire N__53592;
    wire N__53591;
    wire N__53584;
    wire N__53583;
    wire N__53582;
    wire N__53575;
    wire N__53574;
    wire N__53573;
    wire N__53566;
    wire N__53565;
    wire N__53564;
    wire N__53557;
    wire N__53556;
    wire N__53555;
    wire N__53548;
    wire N__53547;
    wire N__53546;
    wire N__53539;
    wire N__53538;
    wire N__53537;
    wire N__53530;
    wire N__53529;
    wire N__53528;
    wire N__53521;
    wire N__53520;
    wire N__53519;
    wire N__53512;
    wire N__53511;
    wire N__53510;
    wire N__53503;
    wire N__53502;
    wire N__53501;
    wire N__53494;
    wire N__53493;
    wire N__53492;
    wire N__53485;
    wire N__53484;
    wire N__53483;
    wire N__53476;
    wire N__53475;
    wire N__53474;
    wire N__53457;
    wire N__53454;
    wire N__53451;
    wire N__53450;
    wire N__53449;
    wire N__53446;
    wire N__53443;
    wire N__53440;
    wire N__53437;
    wire N__53436;
    wire N__53433;
    wire N__53430;
    wire N__53427;
    wire N__53424;
    wire N__53415;
    wire N__53414;
    wire N__53411;
    wire N__53410;
    wire N__53407;
    wire N__53406;
    wire N__53405;
    wire N__53402;
    wire N__53399;
    wire N__53396;
    wire N__53395;
    wire N__53390;
    wire N__53387;
    wire N__53382;
    wire N__53379;
    wire N__53372;
    wire N__53369;
    wire N__53364;
    wire N__53361;
    wire N__53358;
    wire N__53357;
    wire N__53354;
    wire N__53351;
    wire N__53346;
    wire N__53343;
    wire N__53340;
    wire N__53337;
    wire N__53336;
    wire N__53335;
    wire N__53332;
    wire N__53331;
    wire N__53326;
    wire N__53323;
    wire N__53322;
    wire N__53319;
    wire N__53316;
    wire N__53313;
    wire N__53310;
    wire N__53305;
    wire N__53298;
    wire N__53295;
    wire N__53292;
    wire N__53289;
    wire N__53286;
    wire N__53283;
    wire N__53282;
    wire N__53281;
    wire N__53280;
    wire N__53279;
    wire N__53278;
    wire N__53277;
    wire N__53276;
    wire N__53275;
    wire N__53274;
    wire N__53273;
    wire N__53272;
    wire N__53271;
    wire N__53270;
    wire N__53269;
    wire N__53268;
    wire N__53267;
    wire N__53266;
    wire N__53265;
    wire N__53264;
    wire N__53263;
    wire N__53262;
    wire N__53261;
    wire N__53260;
    wire N__53259;
    wire N__53258;
    wire N__53257;
    wire N__53256;
    wire N__53255;
    wire N__53254;
    wire N__53253;
    wire N__53252;
    wire N__53251;
    wire N__53250;
    wire N__53249;
    wire N__53248;
    wire N__53247;
    wire N__53246;
    wire N__53245;
    wire N__53244;
    wire N__53243;
    wire N__53242;
    wire N__53241;
    wire N__53154;
    wire N__53151;
    wire N__53148;
    wire N__53147;
    wire N__53146;
    wire N__53145;
    wire N__53144;
    wire N__53143;
    wire N__53142;
    wire N__53141;
    wire N__53140;
    wire N__53139;
    wire N__53138;
    wire N__53137;
    wire N__53136;
    wire N__53135;
    wire N__53134;
    wire N__53133;
    wire N__53132;
    wire N__53131;
    wire N__53130;
    wire N__53129;
    wire N__53128;
    wire N__53127;
    wire N__53126;
    wire N__53125;
    wire N__53124;
    wire N__53123;
    wire N__53122;
    wire N__53121;
    wire N__53120;
    wire N__53119;
    wire N__53118;
    wire N__53117;
    wire N__53116;
    wire N__53115;
    wire N__53114;
    wire N__53113;
    wire N__53112;
    wire N__53111;
    wire N__53110;
    wire N__53109;
    wire N__53108;
    wire N__53107;
    wire N__53106;
    wire N__53105;
    wire N__53104;
    wire N__53103;
    wire N__53102;
    wire N__53101;
    wire N__53100;
    wire N__53099;
    wire N__53098;
    wire N__53097;
    wire N__53096;
    wire N__53095;
    wire N__53094;
    wire N__53093;
    wire N__53092;
    wire N__53091;
    wire N__53090;
    wire N__53089;
    wire N__53088;
    wire N__53087;
    wire N__53086;
    wire N__53085;
    wire N__53084;
    wire N__53083;
    wire N__53082;
    wire N__53081;
    wire N__53080;
    wire N__53079;
    wire N__53078;
    wire N__53077;
    wire N__53076;
    wire N__53075;
    wire N__53074;
    wire N__53073;
    wire N__53072;
    wire N__53071;
    wire N__53070;
    wire N__53069;
    wire N__53068;
    wire N__53067;
    wire N__53066;
    wire N__53065;
    wire N__53064;
    wire N__53063;
    wire N__53062;
    wire N__53061;
    wire N__53060;
    wire N__53059;
    wire N__53058;
    wire N__53057;
    wire N__53056;
    wire N__53055;
    wire N__53054;
    wire N__53053;
    wire N__53052;
    wire N__53051;
    wire N__53050;
    wire N__53049;
    wire N__53048;
    wire N__53047;
    wire N__53046;
    wire N__53045;
    wire N__53044;
    wire N__53043;
    wire N__53042;
    wire N__53041;
    wire N__53040;
    wire N__53039;
    wire N__53038;
    wire N__53037;
    wire N__53036;
    wire N__53035;
    wire N__53034;
    wire N__53033;
    wire N__53032;
    wire N__53031;
    wire N__53030;
    wire N__53029;
    wire N__53028;
    wire N__53027;
    wire N__53026;
    wire N__53025;
    wire N__53024;
    wire N__53023;
    wire N__53022;
    wire N__53021;
    wire N__53020;
    wire N__53019;
    wire N__53018;
    wire N__53017;
    wire N__53016;
    wire N__53015;
    wire N__53014;
    wire N__53013;
    wire N__53012;
    wire N__53011;
    wire N__53010;
    wire N__53009;
    wire N__53008;
    wire N__53007;
    wire N__53006;
    wire N__53005;
    wire N__53004;
    wire N__53003;
    wire N__53002;
    wire N__53001;
    wire N__53000;
    wire N__52999;
    wire N__52998;
    wire N__52997;
    wire N__52996;
    wire N__52995;
    wire N__52994;
    wire N__52993;
    wire N__52992;
    wire N__52991;
    wire N__52990;
    wire N__52989;
    wire N__52988;
    wire N__52987;
    wire N__52986;
    wire N__52985;
    wire N__52984;
    wire N__52983;
    wire N__52982;
    wire N__52981;
    wire N__52980;
    wire N__52979;
    wire N__52978;
    wire N__52977;
    wire N__52976;
    wire N__52975;
    wire N__52974;
    wire N__52973;
    wire N__52972;
    wire N__52971;
    wire N__52970;
    wire N__52969;
    wire N__52968;
    wire N__52967;
    wire N__52602;
    wire N__52599;
    wire N__52596;
    wire N__52593;
    wire N__52592;
    wire N__52589;
    wire N__52586;
    wire N__52583;
    wire N__52580;
    wire N__52577;
    wire N__52574;
    wire N__52569;
    wire N__52566;
    wire N__52563;
    wire N__52560;
    wire N__52557;
    wire N__52554;
    wire N__52551;
    wire N__52548;
    wire N__52547;
    wire N__52542;
    wire N__52541;
    wire N__52540;
    wire N__52537;
    wire N__52534;
    wire N__52531;
    wire N__52524;
    wire N__52521;
    wire N__52520;
    wire N__52519;
    wire N__52516;
    wire N__52513;
    wire N__52512;
    wire N__52511;
    wire N__52508;
    wire N__52503;
    wire N__52500;
    wire N__52497;
    wire N__52488;
    wire N__52487;
    wire N__52484;
    wire N__52481;
    wire N__52476;
    wire N__52475;
    wire N__52472;
    wire N__52469;
    wire N__52464;
    wire N__52463;
    wire N__52460;
    wire N__52457;
    wire N__52454;
    wire N__52449;
    wire N__52446;
    wire N__52445;
    wire N__52444;
    wire N__52441;
    wire N__52438;
    wire N__52435;
    wire N__52430;
    wire N__52425;
    wire N__52422;
    wire N__52421;
    wire N__52420;
    wire N__52419;
    wire N__52416;
    wire N__52415;
    wire N__52414;
    wire N__52407;
    wire N__52404;
    wire N__52401;
    wire N__52398;
    wire N__52395;
    wire N__52390;
    wire N__52387;
    wire N__52384;
    wire N__52381;
    wire N__52378;
    wire N__52375;
    wire N__52372;
    wire N__52369;
    wire N__52362;
    wire N__52359;
    wire N__52356;
    wire N__52353;
    wire N__52350;
    wire N__52347;
    wire N__52344;
    wire N__52343;
    wire N__52340;
    wire N__52337;
    wire N__52334;
    wire N__52331;
    wire N__52328;
    wire N__52325;
    wire N__52320;
    wire N__52317;
    wire N__52314;
    wire N__52311;
    wire N__52308;
    wire N__52305;
    wire N__52304;
    wire N__52301;
    wire N__52298;
    wire N__52297;
    wire N__52296;
    wire N__52291;
    wire N__52288;
    wire N__52285;
    wire N__52278;
    wire N__52275;
    wire N__52272;
    wire N__52269;
    wire N__52266;
    wire N__52263;
    wire N__52260;
    wire N__52257;
    wire N__52254;
    wire N__52253;
    wire N__52250;
    wire N__52247;
    wire N__52244;
    wire N__52241;
    wire N__52236;
    wire N__52233;
    wire N__52232;
    wire N__52229;
    wire N__52226;
    wire N__52225;
    wire N__52222;
    wire N__52219;
    wire N__52216;
    wire N__52213;
    wire N__52206;
    wire N__52203;
    wire N__52200;
    wire N__52199;
    wire N__52194;
    wire N__52193;
    wire N__52190;
    wire N__52187;
    wire N__52184;
    wire N__52179;
    wire N__52176;
    wire N__52173;
    wire N__52170;
    wire N__52167;
    wire N__52164;
    wire N__52161;
    wire N__52160;
    wire N__52159;
    wire N__52158;
    wire N__52157;
    wire N__52156;
    wire N__52155;
    wire N__52154;
    wire N__52153;
    wire N__52152;
    wire N__52151;
    wire N__52150;
    wire N__52149;
    wire N__52148;
    wire N__52147;
    wire N__52146;
    wire N__52145;
    wire N__52144;
    wire N__52143;
    wire N__52142;
    wire N__52141;
    wire N__52140;
    wire N__52139;
    wire N__52138;
    wire N__52137;
    wire N__52132;
    wire N__52123;
    wire N__52122;
    wire N__52121;
    wire N__52120;
    wire N__52119;
    wire N__52118;
    wire N__52117;
    wire N__52116;
    wire N__52115;
    wire N__52114;
    wire N__52113;
    wire N__52112;
    wire N__52111;
    wire N__52110;
    wire N__52109;
    wire N__52108;
    wire N__52107;
    wire N__52106;
    wire N__52105;
    wire N__52104;
    wire N__52099;
    wire N__52096;
    wire N__52095;
    wire N__52094;
    wire N__52093;
    wire N__52092;
    wire N__52091;
    wire N__52084;
    wire N__52083;
    wire N__52082;
    wire N__52081;
    wire N__52080;
    wire N__52079;
    wire N__52078;
    wire N__52077;
    wire N__52076;
    wire N__52075;
    wire N__52074;
    wire N__52073;
    wire N__52068;
    wire N__52067;
    wire N__52066;
    wire N__52065;
    wire N__52064;
    wire N__52059;
    wire N__52054;
    wire N__52047;
    wire N__52042;
    wire N__52041;
    wire N__52036;
    wire N__52031;
    wire N__52028;
    wire N__52023;
    wire N__52020;
    wire N__52019;
    wire N__52018;
    wire N__52017;
    wire N__52016;
    wire N__52015;
    wire N__52014;
    wire N__52013;
    wire N__52012;
    wire N__52009;
    wire N__52008;
    wire N__52007;
    wire N__52006;
    wire N__52005;
    wire N__52004;
    wire N__52003;
    wire N__52002;
    wire N__52001;
    wire N__52000;
    wire N__51999;
    wire N__51998;
    wire N__51997;
    wire N__51996;
    wire N__51995;
    wire N__51994;
    wire N__51993;
    wire N__51986;
    wire N__51985;
    wire N__51984;
    wire N__51983;
    wire N__51980;
    wire N__51975;
    wire N__51974;
    wire N__51973;
    wire N__51972;
    wire N__51971;
    wire N__51970;
    wire N__51963;
    wire N__51958;
    wire N__51951;
    wire N__51948;
    wire N__51945;
    wire N__51934;
    wire N__51931;
    wire N__51924;
    wire N__51917;
    wire N__51914;
    wire N__51911;
    wire N__51910;
    wire N__51909;
    wire N__51908;
    wire N__51907;
    wire N__51906;
    wire N__51905;
    wire N__51904;
    wire N__51903;
    wire N__51902;
    wire N__51897;
    wire N__51896;
    wire N__51895;
    wire N__51894;
    wire N__51893;
    wire N__51892;
    wire N__51891;
    wire N__51890;
    wire N__51889;
    wire N__51888;
    wire N__51887;
    wire N__51886;
    wire N__51885;
    wire N__51882;
    wire N__51881;
    wire N__51880;
    wire N__51879;
    wire N__51878;
    wire N__51875;
    wire N__51868;
    wire N__51867;
    wire N__51866;
    wire N__51865;
    wire N__51864;
    wire N__51861;
    wire N__51858;
    wire N__51851;
    wire N__51848;
    wire N__51843;
    wire N__51836;
    wire N__51831;
    wire N__51826;
    wire N__51819;
    wire N__51818;
    wire N__51817;
    wire N__51816;
    wire N__51815;
    wire N__51814;
    wire N__51813;
    wire N__51812;
    wire N__51811;
    wire N__51810;
    wire N__51809;
    wire N__51808;
    wire N__51805;
    wire N__51804;
    wire N__51803;
    wire N__51802;
    wire N__51801;
    wire N__51794;
    wire N__51785;
    wire N__51778;
    wire N__51773;
    wire N__51772;
    wire N__51771;
    wire N__51770;
    wire N__51763;
    wire N__51758;
    wire N__51755;
    wire N__51752;
    wire N__51747;
    wire N__51742;
    wire N__51737;
    wire N__51730;
    wire N__51727;
    wire N__51722;
    wire N__51711;
    wire N__51704;
    wire N__51695;
    wire N__51684;
    wire N__51681;
    wire N__51678;
    wire N__51671;
    wire N__51666;
    wire N__51663;
    wire N__51656;
    wire N__51651;
    wire N__51648;
    wire N__51645;
    wire N__51638;
    wire N__51633;
    wire N__51624;
    wire N__51617;
    wire N__51610;
    wire N__51603;
    wire N__51602;
    wire N__51601;
    wire N__51600;
    wire N__51599;
    wire N__51598;
    wire N__51597;
    wire N__51596;
    wire N__51595;
    wire N__51594;
    wire N__51589;
    wire N__51582;
    wire N__51577;
    wire N__51570;
    wire N__51565;
    wire N__51556;
    wire N__51555;
    wire N__51554;
    wire N__51553;
    wire N__51552;
    wire N__51551;
    wire N__51542;
    wire N__51541;
    wire N__51540;
    wire N__51539;
    wire N__51538;
    wire N__51537;
    wire N__51530;
    wire N__51521;
    wire N__51514;
    wire N__51503;
    wire N__51502;
    wire N__51501;
    wire N__51496;
    wire N__51495;
    wire N__51494;
    wire N__51493;
    wire N__51490;
    wire N__51481;
    wire N__51480;
    wire N__51479;
    wire N__51478;
    wire N__51477;
    wire N__51472;
    wire N__51461;
    wire N__51454;
    wire N__51443;
    wire N__51434;
    wire N__51421;
    wire N__51412;
    wire N__51409;
    wire N__51406;
    wire N__51395;
    wire N__51386;
    wire N__51383;
    wire N__51380;
    wire N__51377;
    wire N__51370;
    wire N__51365;
    wire N__51362;
    wire N__51355;
    wire N__51348;
    wire N__51339;
    wire N__51334;
    wire N__51329;
    wire N__51306;
    wire N__51303;
    wire N__51300;
    wire N__51297;
    wire N__51294;
    wire N__51291;
    wire N__51288;
    wire N__51285;
    wire N__51282;
    wire N__51279;
    wire N__51276;
    wire N__51273;
    wire N__51272;
    wire N__51271;
    wire N__51270;
    wire N__51269;
    wire N__51268;
    wire N__51267;
    wire N__51266;
    wire N__51263;
    wire N__51262;
    wire N__51261;
    wire N__51260;
    wire N__51259;
    wire N__51258;
    wire N__51257;
    wire N__51254;
    wire N__51253;
    wire N__51252;
    wire N__51249;
    wire N__51248;
    wire N__51247;
    wire N__51246;
    wire N__51243;
    wire N__51242;
    wire N__51241;
    wire N__51240;
    wire N__51239;
    wire N__51236;
    wire N__51233;
    wire N__51232;
    wire N__51229;
    wire N__51226;
    wire N__51223;
    wire N__51220;
    wire N__51217;
    wire N__51216;
    wire N__51213;
    wire N__51210;
    wire N__51207;
    wire N__51204;
    wire N__51203;
    wire N__51200;
    wire N__51197;
    wire N__51194;
    wire N__51191;
    wire N__51188;
    wire N__51185;
    wire N__51182;
    wire N__51181;
    wire N__51178;
    wire N__51175;
    wire N__51172;
    wire N__51169;
    wire N__51168;
    wire N__51165;
    wire N__51164;
    wire N__51159;
    wire N__51158;
    wire N__51157;
    wire N__51156;
    wire N__51155;
    wire N__51152;
    wire N__51147;
    wire N__51140;
    wire N__51139;
    wire N__51138;
    wire N__51135;
    wire N__51134;
    wire N__51133;
    wire N__51132;
    wire N__51127;
    wire N__51122;
    wire N__51119;
    wire N__51112;
    wire N__51105;
    wire N__51102;
    wire N__51101;
    wire N__51100;
    wire N__51099;
    wire N__51096;
    wire N__51087;
    wire N__51084;
    wire N__51083;
    wire N__51082;
    wire N__51081;
    wire N__51080;
    wire N__51079;
    wire N__51078;
    wire N__51075;
    wire N__51072;
    wire N__51069;
    wire N__51066;
    wire N__51063;
    wire N__51060;
    wire N__51057;
    wire N__51054;
    wire N__51051;
    wire N__51048;
    wire N__51045;
    wire N__51042;
    wire N__51041;
    wire N__51040;
    wire N__51037;
    wire N__51034;
    wire N__51031;
    wire N__51028;
    wire N__51027;
    wire N__51026;
    wire N__51025;
    wire N__51024;
    wire N__51017;
    wire N__51010;
    wire N__51007;
    wire N__51004;
    wire N__51001;
    wire N__50994;
    wire N__50991;
    wire N__50988;
    wire N__50987;
    wire N__50986;
    wire N__50983;
    wire N__50982;
    wire N__50981;
    wire N__50978;
    wire N__50975;
    wire N__50972;
    wire N__50967;
    wire N__50956;
    wire N__50953;
    wire N__50944;
    wire N__50941;
    wire N__50938;
    wire N__50929;
    wire N__50926;
    wire N__50923;
    wire N__50920;
    wire N__50917;
    wire N__50914;
    wire N__50905;
    wire N__50898;
    wire N__50895;
    wire N__50892;
    wire N__50889;
    wire N__50886;
    wire N__50883;
    wire N__50882;
    wire N__50881;
    wire N__50874;
    wire N__50873;
    wire N__50872;
    wire N__50867;
    wire N__50860;
    wire N__50857;
    wire N__50846;
    wire N__50835;
    wire N__50828;
    wire N__50825;
    wire N__50822;
    wire N__50819;
    wire N__50814;
    wire N__50807;
    wire N__50804;
    wire N__50801;
    wire N__50796;
    wire N__50789;
    wire N__50778;
    wire N__50775;
    wire N__50772;
    wire N__50771;
    wire N__50770;
    wire N__50769;
    wire N__50766;
    wire N__50763;
    wire N__50762;
    wire N__50761;
    wire N__50758;
    wire N__50755;
    wire N__50754;
    wire N__50753;
    wire N__50750;
    wire N__50747;
    wire N__50744;
    wire N__50741;
    wire N__50740;
    wire N__50735;
    wire N__50734;
    wire N__50733;
    wire N__50732;
    wire N__50729;
    wire N__50726;
    wire N__50725;
    wire N__50724;
    wire N__50723;
    wire N__50714;
    wire N__50711;
    wire N__50710;
    wire N__50709;
    wire N__50708;
    wire N__50707;
    wire N__50704;
    wire N__50701;
    wire N__50698;
    wire N__50695;
    wire N__50694;
    wire N__50693;
    wire N__50692;
    wire N__50691;
    wire N__50688;
    wire N__50687;
    wire N__50686;
    wire N__50685;
    wire N__50682;
    wire N__50679;
    wire N__50678;
    wire N__50677;
    wire N__50676;
    wire N__50675;
    wire N__50674;
    wire N__50673;
    wire N__50672;
    wire N__50669;
    wire N__50666;
    wire N__50665;
    wire N__50664;
    wire N__50659;
    wire N__50656;
    wire N__50653;
    wire N__50650;
    wire N__50647;
    wire N__50638;
    wire N__50635;
    wire N__50632;
    wire N__50629;
    wire N__50626;
    wire N__50625;
    wire N__50622;
    wire N__50619;
    wire N__50616;
    wire N__50613;
    wire N__50608;
    wire N__50605;
    wire N__50602;
    wire N__50601;
    wire N__50600;
    wire N__50599;
    wire N__50596;
    wire N__50593;
    wire N__50592;
    wire N__50589;
    wire N__50586;
    wire N__50585;
    wire N__50584;
    wire N__50583;
    wire N__50582;
    wire N__50581;
    wire N__50580;
    wire N__50577;
    wire N__50576;
    wire N__50575;
    wire N__50574;
    wire N__50573;
    wire N__50572;
    wire N__50567;
    wire N__50564;
    wire N__50561;
    wire N__50560;
    wire N__50549;
    wire N__50542;
    wire N__50537;
    wire N__50534;
    wire N__50525;
    wire N__50518;
    wire N__50515;
    wire N__50512;
    wire N__50509;
    wire N__50504;
    wire N__50501;
    wire N__50500;
    wire N__50497;
    wire N__50494;
    wire N__50491;
    wire N__50488;
    wire N__50485;
    wire N__50482;
    wire N__50479;
    wire N__50476;
    wire N__50473;
    wire N__50470;
    wire N__50467;
    wire N__50464;
    wire N__50461;
    wire N__50458;
    wire N__50457;
    wire N__50456;
    wire N__50455;
    wire N__50454;
    wire N__50451;
    wire N__50448;
    wire N__50445;
    wire N__50442;
    wire N__50439;
    wire N__50432;
    wire N__50423;
    wire N__50422;
    wire N__50415;
    wire N__50412;
    wire N__50393;
    wire N__50386;
    wire N__50381;
    wire N__50378;
    wire N__50375;
    wire N__50372;
    wire N__50369;
    wire N__50360;
    wire N__50355;
    wire N__50352;
    wire N__50349;
    wire N__50342;
    wire N__50327;
    wire N__50316;
    wire N__50313;
    wire N__50310;
    wire N__50309;
    wire N__50308;
    wire N__50307;
    wire N__50306;
    wire N__50305;
    wire N__50302;
    wire N__50301;
    wire N__50300;
    wire N__50299;
    wire N__50296;
    wire N__50293;
    wire N__50292;
    wire N__50291;
    wire N__50288;
    wire N__50287;
    wire N__50286;
    wire N__50285;
    wire N__50284;
    wire N__50283;
    wire N__50282;
    wire N__50281;
    wire N__50278;
    wire N__50275;
    wire N__50274;
    wire N__50271;
    wire N__50268;
    wire N__50265;
    wire N__50264;
    wire N__50263;
    wire N__50262;
    wire N__50261;
    wire N__50258;
    wire N__50257;
    wire N__50256;
    wire N__50255;
    wire N__50250;
    wire N__50247;
    wire N__50244;
    wire N__50243;
    wire N__50242;
    wire N__50241;
    wire N__50240;
    wire N__50237;
    wire N__50234;
    wire N__50231;
    wire N__50230;
    wire N__50227;
    wire N__50224;
    wire N__50221;
    wire N__50218;
    wire N__50215;
    wire N__50210;
    wire N__50207;
    wire N__50200;
    wire N__50197;
    wire N__50194;
    wire N__50191;
    wire N__50188;
    wire N__50187;
    wire N__50184;
    wire N__50181;
    wire N__50180;
    wire N__50179;
    wire N__50178;
    wire N__50175;
    wire N__50174;
    wire N__50171;
    wire N__50164;
    wire N__50161;
    wire N__50158;
    wire N__50155;
    wire N__50152;
    wire N__50151;
    wire N__50144;
    wire N__50141;
    wire N__50132;
    wire N__50129;
    wire N__50124;
    wire N__50123;
    wire N__50112;
    wire N__50109;
    wire N__50108;
    wire N__50107;
    wire N__50106;
    wire N__50105;
    wire N__50100;
    wire N__50097;
    wire N__50094;
    wire N__50093;
    wire N__50092;
    wire N__50091;
    wire N__50090;
    wire N__50087;
    wire N__50084;
    wire N__50081;
    wire N__50080;
    wire N__50079;
    wire N__50078;
    wire N__50077;
    wire N__50074;
    wire N__50063;
    wire N__50060;
    wire N__50055;
    wire N__50052;
    wire N__50047;
    wire N__50044;
    wire N__50039;
    wire N__50036;
    wire N__50033;
    wire N__50030;
    wire N__50027;
    wire N__50026;
    wire N__50025;
    wire N__50024;
    wire N__50023;
    wire N__50016;
    wire N__50013;
    wire N__50010;
    wire N__50007;
    wire N__50006;
    wire N__50005;
    wire N__50004;
    wire N__50001;
    wire N__49998;
    wire N__49993;
    wire N__49990;
    wire N__49987;
    wire N__49984;
    wire N__49981;
    wire N__49974;
    wire N__49971;
    wire N__49964;
    wire N__49955;
    wire N__49952;
    wire N__49949;
    wire N__49946;
    wire N__49943;
    wire N__49940;
    wire N__49931;
    wire N__49928;
    wire N__49925;
    wire N__49922;
    wire N__49907;
    wire N__49906;
    wire N__49903;
    wire N__49896;
    wire N__49885;
    wire N__49878;
    wire N__49873;
    wire N__49870;
    wire N__49857;
    wire N__49854;
    wire N__49851;
    wire N__49848;
    wire N__49845;
    wire N__49844;
    wire N__49843;
    wire N__49842;
    wire N__49841;
    wire N__49838;
    wire N__49837;
    wire N__49836;
    wire N__49835;
    wire N__49834;
    wire N__49833;
    wire N__49830;
    wire N__49827;
    wire N__49826;
    wire N__49825;
    wire N__49824;
    wire N__49823;
    wire N__49822;
    wire N__49821;
    wire N__49820;
    wire N__49819;
    wire N__49818;
    wire N__49815;
    wire N__49812;
    wire N__49811;
    wire N__49808;
    wire N__49805;
    wire N__49802;
    wire N__49799;
    wire N__49798;
    wire N__49797;
    wire N__49796;
    wire N__49795;
    wire N__49794;
    wire N__49791;
    wire N__49790;
    wire N__49787;
    wire N__49786;
    wire N__49785;
    wire N__49784;
    wire N__49779;
    wire N__49776;
    wire N__49773;
    wire N__49770;
    wire N__49769;
    wire N__49768;
    wire N__49767;
    wire N__49766;
    wire N__49765;
    wire N__49762;
    wire N__49759;
    wire N__49756;
    wire N__49753;
    wire N__49750;
    wire N__49747;
    wire N__49744;
    wire N__49741;
    wire N__49738;
    wire N__49737;
    wire N__49736;
    wire N__49735;
    wire N__49734;
    wire N__49729;
    wire N__49726;
    wire N__49723;
    wire N__49720;
    wire N__49717;
    wire N__49714;
    wire N__49711;
    wire N__49708;
    wire N__49705;
    wire N__49704;
    wire N__49703;
    wire N__49702;
    wire N__49699;
    wire N__49696;
    wire N__49693;
    wire N__49690;
    wire N__49689;
    wire N__49686;
    wire N__49677;
    wire N__49674;
    wire N__49671;
    wire N__49668;
    wire N__49665;
    wire N__49662;
    wire N__49661;
    wire N__49652;
    wire N__49651;
    wire N__49646;
    wire N__49639;
    wire N__49636;
    wire N__49633;
    wire N__49630;
    wire N__49627;
    wire N__49626;
    wire N__49611;
    wire N__49610;
    wire N__49609;
    wire N__49608;
    wire N__49605;
    wire N__49602;
    wire N__49599;
    wire N__49596;
    wire N__49593;
    wire N__49592;
    wire N__49591;
    wire N__49590;
    wire N__49587;
    wire N__49582;
    wire N__49579;
    wire N__49576;
    wire N__49575;
    wire N__49574;
    wire N__49573;
    wire N__49572;
    wire N__49571;
    wire N__49568;
    wire N__49555;
    wire N__49552;
    wire N__49549;
    wire N__49546;
    wire N__49533;
    wire N__49530;
    wire N__49527;
    wire N__49524;
    wire N__49521;
    wire N__49518;
    wire N__49515;
    wire N__49506;
    wire N__49503;
    wire N__49500;
    wire N__49497;
    wire N__49496;
    wire N__49493;
    wire N__49486;
    wire N__49483;
    wire N__49480;
    wire N__49477;
    wire N__49474;
    wire N__49471;
    wire N__49464;
    wire N__49459;
    wire N__49454;
    wire N__49445;
    wire N__49434;
    wire N__49431;
    wire N__49416;
    wire N__49415;
    wire N__49412;
    wire N__49405;
    wire N__49400;
    wire N__49397;
    wire N__49394;
    wire N__49383;
    wire N__49380;
    wire N__49377;
    wire N__49374;
    wire N__49371;
    wire N__49368;
    wire N__49367;
    wire N__49364;
    wire N__49363;
    wire N__49362;
    wire N__49361;
    wire N__49360;
    wire N__49359;
    wire N__49358;
    wire N__49357;
    wire N__49356;
    wire N__49355;
    wire N__49354;
    wire N__49351;
    wire N__49348;
    wire N__49347;
    wire N__49346;
    wire N__49345;
    wire N__49344;
    wire N__49343;
    wire N__49340;
    wire N__49337;
    wire N__49336;
    wire N__49335;
    wire N__49334;
    wire N__49331;
    wire N__49328;
    wire N__49327;
    wire N__49326;
    wire N__49323;
    wire N__49322;
    wire N__49319;
    wire N__49316;
    wire N__49313;
    wire N__49312;
    wire N__49309;
    wire N__49308;
    wire N__49307;
    wire N__49306;
    wire N__49305;
    wire N__49302;
    wire N__49297;
    wire N__49294;
    wire N__49291;
    wire N__49288;
    wire N__49285;
    wire N__49282;
    wire N__49281;
    wire N__49276;
    wire N__49273;
    wire N__49270;
    wire N__49267;
    wire N__49264;
    wire N__49261;
    wire N__49260;
    wire N__49257;
    wire N__49254;
    wire N__49251;
    wire N__49248;
    wire N__49241;
    wire N__49238;
    wire N__49235;
    wire N__49232;
    wire N__49231;
    wire N__49230;
    wire N__49227;
    wire N__49226;
    wire N__49223;
    wire N__49222;
    wire N__49219;
    wire N__49208;
    wire N__49207;
    wire N__49202;
    wire N__49199;
    wire N__49190;
    wire N__49189;
    wire N__49188;
    wire N__49187;
    wire N__49186;
    wire N__49181;
    wire N__49178;
    wire N__49177;
    wire N__49172;
    wire N__49167;
    wire N__49166;
    wire N__49165;
    wire N__49160;
    wire N__49155;
    wire N__49152;
    wire N__49149;
    wire N__49146;
    wire N__49145;
    wire N__49144;
    wire N__49141;
    wire N__49138;
    wire N__49135;
    wire N__49132;
    wire N__49131;
    wire N__49130;
    wire N__49129;
    wire N__49126;
    wire N__49123;
    wire N__49120;
    wire N__49115;
    wire N__49112;
    wire N__49111;
    wire N__49110;
    wire N__49109;
    wire N__49106;
    wire N__49103;
    wire N__49100;
    wire N__49095;
    wire N__49092;
    wire N__49091;
    wire N__49088;
    wire N__49085;
    wire N__49082;
    wire N__49079;
    wire N__49078;
    wire N__49077;
    wire N__49076;
    wire N__49075;
    wire N__49068;
    wire N__49063;
    wire N__49060;
    wire N__49057;
    wire N__49052;
    wire N__49047;
    wire N__49044;
    wire N__49041;
    wire N__49038;
    wire N__49035;
    wire N__49028;
    wire N__49025;
    wire N__49022;
    wire N__49019;
    wire N__49016;
    wire N__49009;
    wire N__49004;
    wire N__49001;
    wire N__48998;
    wire N__48993;
    wire N__48990;
    wire N__48989;
    wire N__48988;
    wire N__48985;
    wire N__48982;
    wire N__48979;
    wire N__48976;
    wire N__48973;
    wire N__48962;
    wire N__48949;
    wire N__48930;
    wire N__48927;
    wire N__48924;
    wire N__48911;
    wire N__48910;
    wire N__48907;
    wire N__48904;
    wire N__48897;
    wire N__48894;
    wire N__48885;
    wire N__48882;
    wire N__48879;
    wire N__48876;
    wire N__48873;
    wire N__48870;
    wire N__48867;
    wire N__48866;
    wire N__48863;
    wire N__48860;
    wire N__48857;
    wire N__48854;
    wire N__48851;
    wire N__48848;
    wire N__48843;
    wire N__48842;
    wire N__48841;
    wire N__48838;
    wire N__48835;
    wire N__48834;
    wire N__48833;
    wire N__48832;
    wire N__48831;
    wire N__48830;
    wire N__48827;
    wire N__48822;
    wire N__48819;
    wire N__48818;
    wire N__48817;
    wire N__48816;
    wire N__48813;
    wire N__48812;
    wire N__48809;
    wire N__48808;
    wire N__48805;
    wire N__48802;
    wire N__48801;
    wire N__48800;
    wire N__48799;
    wire N__48798;
    wire N__48797;
    wire N__48790;
    wire N__48787;
    wire N__48786;
    wire N__48783;
    wire N__48780;
    wire N__48779;
    wire N__48778;
    wire N__48777;
    wire N__48776;
    wire N__48773;
    wire N__48770;
    wire N__48769;
    wire N__48768;
    wire N__48765;
    wire N__48762;
    wire N__48757;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48747;
    wire N__48746;
    wire N__48745;
    wire N__48744;
    wire N__48743;
    wire N__48742;
    wire N__48741;
    wire N__48740;
    wire N__48739;
    wire N__48738;
    wire N__48737;
    wire N__48736;
    wire N__48733;
    wire N__48730;
    wire N__48729;
    wire N__48728;
    wire N__48723;
    wire N__48720;
    wire N__48719;
    wire N__48718;
    wire N__48713;
    wire N__48710;
    wire N__48707;
    wire N__48706;
    wire N__48705;
    wire N__48702;
    wire N__48699;
    wire N__48694;
    wire N__48691;
    wire N__48688;
    wire N__48683;
    wire N__48678;
    wire N__48673;
    wire N__48672;
    wire N__48671;
    wire N__48670;
    wire N__48669;
    wire N__48668;
    wire N__48667;
    wire N__48664;
    wire N__48661;
    wire N__48658;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48643;
    wire N__48640;
    wire N__48637;
    wire N__48634;
    wire N__48633;
    wire N__48630;
    wire N__48627;
    wire N__48624;
    wire N__48621;
    wire N__48618;
    wire N__48613;
    wire N__48610;
    wire N__48607;
    wire N__48600;
    wire N__48599;
    wire N__48598;
    wire N__48597;
    wire N__48594;
    wire N__48593;
    wire N__48592;
    wire N__48589;
    wire N__48586;
    wire N__48583;
    wire N__48580;
    wire N__48577;
    wire N__48576;
    wire N__48575;
    wire N__48572;
    wire N__48569;
    wire N__48564;
    wire N__48561;
    wire N__48558;
    wire N__48555;
    wire N__48552;
    wire N__48549;
    wire N__48546;
    wire N__48545;
    wire N__48540;
    wire N__48531;
    wire N__48520;
    wire N__48517;
    wire N__48512;
    wire N__48507;
    wire N__48502;
    wire N__48495;
    wire N__48492;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48480;
    wire N__48477;
    wire N__48474;
    wire N__48465;
    wire N__48462;
    wire N__48459;
    wire N__48456;
    wire N__48453;
    wire N__48450;
    wire N__48447;
    wire N__48436;
    wire N__48433;
    wire N__48428;
    wire N__48425;
    wire N__48420;
    wire N__48413;
    wire N__48404;
    wire N__48401;
    wire N__48394;
    wire N__48381;
    wire N__48378;
    wire N__48367;
    wire N__48358;
    wire N__48351;
    wire N__48348;
    wire N__48345;
    wire N__48342;
    wire N__48341;
    wire N__48340;
    wire N__48339;
    wire N__48338;
    wire N__48337;
    wire N__48336;
    wire N__48333;
    wire N__48332;
    wire N__48331;
    wire N__48330;
    wire N__48329;
    wire N__48326;
    wire N__48325;
    wire N__48324;
    wire N__48321;
    wire N__48318;
    wire N__48315;
    wire N__48312;
    wire N__48311;
    wire N__48310;
    wire N__48307;
    wire N__48306;
    wire N__48305;
    wire N__48304;
    wire N__48303;
    wire N__48300;
    wire N__48297;
    wire N__48294;
    wire N__48291;
    wire N__48288;
    wire N__48285;
    wire N__48282;
    wire N__48281;
    wire N__48280;
    wire N__48279;
    wire N__48278;
    wire N__48275;
    wire N__48274;
    wire N__48273;
    wire N__48272;
    wire N__48269;
    wire N__48262;
    wire N__48259;
    wire N__48256;
    wire N__48255;
    wire N__48254;
    wire N__48251;
    wire N__48248;
    wire N__48245;
    wire N__48244;
    wire N__48241;
    wire N__48238;
    wire N__48237;
    wire N__48236;
    wire N__48235;
    wire N__48234;
    wire N__48233;
    wire N__48232;
    wire N__48231;
    wire N__48230;
    wire N__48229;
    wire N__48228;
    wire N__48227;
    wire N__48220;
    wire N__48215;
    wire N__48214;
    wire N__48213;
    wire N__48212;
    wire N__48211;
    wire N__48210;
    wire N__48205;
    wire N__48202;
    wire N__48199;
    wire N__48196;
    wire N__48193;
    wire N__48192;
    wire N__48191;
    wire N__48190;
    wire N__48189;
    wire N__48186;
    wire N__48183;
    wire N__48180;
    wire N__48177;
    wire N__48168;
    wire N__48165;
    wire N__48162;
    wire N__48161;
    wire N__48160;
    wire N__48159;
    wire N__48154;
    wire N__48153;
    wire N__48150;
    wire N__48147;
    wire N__48146;
    wire N__48143;
    wire N__48140;
    wire N__48137;
    wire N__48134;
    wire N__48131;
    wire N__48128;
    wire N__48125;
    wire N__48124;
    wire N__48121;
    wire N__48118;
    wire N__48115;
    wire N__48112;
    wire N__48109;
    wire N__48106;
    wire N__48101;
    wire N__48098;
    wire N__48095;
    wire N__48092;
    wire N__48089;
    wire N__48086;
    wire N__48075;
    wire N__48072;
    wire N__48069;
    wire N__48066;
    wire N__48063;
    wire N__48062;
    wire N__48053;
    wire N__48046;
    wire N__48043;
    wire N__48040;
    wire N__48037;
    wire N__48034;
    wire N__48031;
    wire N__48026;
    wire N__48023;
    wire N__48014;
    wire N__48007;
    wire N__48004;
    wire N__48001;
    wire N__47996;
    wire N__47989;
    wire N__47976;
    wire N__47975;
    wire N__47972;
    wire N__47963;
    wire N__47960;
    wire N__47949;
    wire N__47948;
    wire N__47943;
    wire N__47938;
    wire N__47931;
    wire N__47926;
    wire N__47923;
    wire N__47920;
    wire N__47917;
    wire N__47908;
    wire N__47905;
    wire N__47902;
    wire N__47899;
    wire N__47896;
    wire N__47887;
    wire N__47884;
    wire N__47881;
    wire N__47868;
    wire N__47865;
    wire N__47862;
    wire N__47859;
    wire N__47856;
    wire N__47853;
    wire N__47852;
    wire N__47851;
    wire N__47850;
    wire N__47849;
    wire N__47848;
    wire N__47847;
    wire N__47846;
    wire N__47845;
    wire N__47844;
    wire N__47843;
    wire N__47842;
    wire N__47841;
    wire N__47840;
    wire N__47839;
    wire N__47838;
    wire N__47837;
    wire N__47836;
    wire N__47835;
    wire N__47834;
    wire N__47833;
    wire N__47832;
    wire N__47831;
    wire N__47830;
    wire N__47829;
    wire N__47828;
    wire N__47827;
    wire N__47826;
    wire N__47825;
    wire N__47824;
    wire N__47823;
    wire N__47822;
    wire N__47821;
    wire N__47820;
    wire N__47819;
    wire N__47818;
    wire N__47817;
    wire N__47816;
    wire N__47815;
    wire N__47814;
    wire N__47813;
    wire N__47812;
    wire N__47811;
    wire N__47810;
    wire N__47809;
    wire N__47808;
    wire N__47807;
    wire N__47806;
    wire N__47805;
    wire N__47804;
    wire N__47803;
    wire N__47802;
    wire N__47801;
    wire N__47800;
    wire N__47799;
    wire N__47798;
    wire N__47797;
    wire N__47796;
    wire N__47795;
    wire N__47794;
    wire N__47793;
    wire N__47792;
    wire N__47791;
    wire N__47790;
    wire N__47789;
    wire N__47788;
    wire N__47787;
    wire N__47786;
    wire N__47785;
    wire N__47784;
    wire N__47783;
    wire N__47782;
    wire N__47781;
    wire N__47780;
    wire N__47779;
    wire N__47778;
    wire N__47777;
    wire N__47776;
    wire N__47775;
    wire N__47774;
    wire N__47773;
    wire N__47772;
    wire N__47771;
    wire N__47770;
    wire N__47769;
    wire N__47768;
    wire N__47767;
    wire N__47766;
    wire N__47765;
    wire N__47764;
    wire N__47763;
    wire N__47762;
    wire N__47761;
    wire N__47760;
    wire N__47759;
    wire N__47758;
    wire N__47757;
    wire N__47756;
    wire N__47755;
    wire N__47754;
    wire N__47753;
    wire N__47752;
    wire N__47751;
    wire N__47750;
    wire N__47749;
    wire N__47748;
    wire N__47747;
    wire N__47746;
    wire N__47745;
    wire N__47744;
    wire N__47743;
    wire N__47742;
    wire N__47741;
    wire N__47740;
    wire N__47739;
    wire N__47738;
    wire N__47737;
    wire N__47736;
    wire N__47735;
    wire N__47734;
    wire N__47733;
    wire N__47732;
    wire N__47731;
    wire N__47730;
    wire N__47729;
    wire N__47728;
    wire N__47727;
    wire N__47726;
    wire N__47725;
    wire N__47724;
    wire N__47723;
    wire N__47722;
    wire N__47721;
    wire N__47720;
    wire N__47719;
    wire N__47718;
    wire N__47717;
    wire N__47716;
    wire N__47715;
    wire N__47714;
    wire N__47713;
    wire N__47712;
    wire N__47711;
    wire N__47710;
    wire N__47709;
    wire N__47708;
    wire N__47707;
    wire N__47706;
    wire N__47705;
    wire N__47704;
    wire N__47703;
    wire N__47702;
    wire N__47397;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47384;
    wire N__47381;
    wire N__47378;
    wire N__47377;
    wire N__47376;
    wire N__47375;
    wire N__47372;
    wire N__47369;
    wire N__47366;
    wire N__47363;
    wire N__47360;
    wire N__47353;
    wire N__47350;
    wire N__47347;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47328;
    wire N__47325;
    wire N__47322;
    wire N__47319;
    wire N__47316;
    wire N__47313;
    wire N__47310;
    wire N__47307;
    wire N__47306;
    wire N__47301;
    wire N__47300;
    wire N__47297;
    wire N__47294;
    wire N__47291;
    wire N__47286;
    wire N__47283;
    wire N__47280;
    wire N__47277;
    wire N__47274;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47262;
    wire N__47259;
    wire N__47256;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47244;
    wire N__47241;
    wire N__47238;
    wire N__47235;
    wire N__47234;
    wire N__47231;
    wire N__47228;
    wire N__47225;
    wire N__47222;
    wire N__47217;
    wire N__47214;
    wire N__47211;
    wire N__47208;
    wire N__47205;
    wire N__47202;
    wire N__47199;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47187;
    wire N__47184;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47172;
    wire N__47169;
    wire N__47166;
    wire N__47163;
    wire N__47160;
    wire N__47157;
    wire N__47154;
    wire N__47151;
    wire N__47150;
    wire N__47149;
    wire N__47148;
    wire N__47147;
    wire N__47144;
    wire N__47141;
    wire N__47140;
    wire N__47139;
    wire N__47138;
    wire N__47137;
    wire N__47136;
    wire N__47135;
    wire N__47134;
    wire N__47133;
    wire N__47132;
    wire N__47131;
    wire N__47130;
    wire N__47127;
    wire N__47126;
    wire N__47123;
    wire N__47120;
    wire N__47119;
    wire N__47118;
    wire N__47117;
    wire N__47112;
    wire N__47109;
    wire N__47106;
    wire N__47103;
    wire N__47100;
    wire N__47099;
    wire N__47096;
    wire N__47093;
    wire N__47090;
    wire N__47089;
    wire N__47088;
    wire N__47085;
    wire N__47082;
    wire N__47081;
    wire N__47078;
    wire N__47075;
    wire N__47074;
    wire N__47073;
    wire N__47072;
    wire N__47071;
    wire N__47068;
    wire N__47065;
    wire N__47064;
    wire N__47063;
    wire N__47062;
    wire N__47057;
    wire N__47054;
    wire N__47053;
    wire N__47050;
    wire N__47047;
    wire N__47046;
    wire N__47045;
    wire N__47034;
    wire N__47031;
    wire N__47024;
    wire N__47021;
    wire N__47018;
    wire N__47017;
    wire N__47016;
    wire N__47013;
    wire N__47010;
    wire N__47007;
    wire N__47004;
    wire N__47001;
    wire N__46998;
    wire N__46995;
    wire N__46994;
    wire N__46993;
    wire N__46990;
    wire N__46987;
    wire N__46986;
    wire N__46985;
    wire N__46984;
    wire N__46983;
    wire N__46980;
    wire N__46977;
    wire N__46974;
    wire N__46971;
    wire N__46970;
    wire N__46967;
    wire N__46962;
    wire N__46959;
    wire N__46958;
    wire N__46957;
    wire N__46956;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46944;
    wire N__46939;
    wire N__46934;
    wire N__46931;
    wire N__46928;
    wire N__46925;
    wire N__46918;
    wire N__46913;
    wire N__46908;
    wire N__46905;
    wire N__46902;
    wire N__46899;
    wire N__46898;
    wire N__46897;
    wire N__46894;
    wire N__46891;
    wire N__46888;
    wire N__46885;
    wire N__46882;
    wire N__46881;
    wire N__46880;
    wire N__46879;
    wire N__46878;
    wire N__46877;
    wire N__46876;
    wire N__46871;
    wire N__46868;
    wire N__46865;
    wire N__46862;
    wire N__46861;
    wire N__46858;
    wire N__46853;
    wire N__46850;
    wire N__46845;
    wire N__46842;
    wire N__46835;
    wire N__46832;
    wire N__46823;
    wire N__46820;
    wire N__46811;
    wire N__46808;
    wire N__46805;
    wire N__46802;
    wire N__46795;
    wire N__46794;
    wire N__46793;
    wire N__46788;
    wire N__46785;
    wire N__46782;
    wire N__46779;
    wire N__46776;
    wire N__46773;
    wire N__46770;
    wire N__46769;
    wire N__46766;
    wire N__46759;
    wire N__46756;
    wire N__46747;
    wire N__46738;
    wire N__46733;
    wire N__46726;
    wire N__46723;
    wire N__46720;
    wire N__46717;
    wire N__46702;
    wire N__46699;
    wire N__46690;
    wire N__46687;
    wire N__46676;
    wire N__46669;
    wire N__46662;
    wire N__46659;
    wire N__46656;
    wire N__46653;
    wire N__46650;
    wire N__46647;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46635;
    wire N__46632;
    wire N__46631;
    wire N__46630;
    wire N__46629;
    wire N__46626;
    wire N__46623;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46598;
    wire N__46595;
    wire N__46590;
    wire N__46587;
    wire N__46584;
    wire N__46581;
    wire N__46578;
    wire N__46575;
    wire N__46574;
    wire N__46573;
    wire N__46570;
    wire N__46569;
    wire N__46568;
    wire N__46567;
    wire N__46566;
    wire N__46565;
    wire N__46564;
    wire N__46563;
    wire N__46560;
    wire N__46559;
    wire N__46556;
    wire N__46551;
    wire N__46538;
    wire N__46535;
    wire N__46532;
    wire N__46529;
    wire N__46528;
    wire N__46525;
    wire N__46522;
    wire N__46519;
    wire N__46514;
    wire N__46513;
    wire N__46512;
    wire N__46511;
    wire N__46508;
    wire N__46505;
    wire N__46502;
    wire N__46497;
    wire N__46490;
    wire N__46487;
    wire N__46486;
    wire N__46485;
    wire N__46482;
    wire N__46479;
    wire N__46474;
    wire N__46471;
    wire N__46468;
    wire N__46465;
    wire N__46452;
    wire N__46451;
    wire N__46450;
    wire N__46449;
    wire N__46446;
    wire N__46445;
    wire N__46442;
    wire N__46439;
    wire N__46438;
    wire N__46435;
    wire N__46432;
    wire N__46429;
    wire N__46428;
    wire N__46425;
    wire N__46422;
    wire N__46419;
    wire N__46418;
    wire N__46415;
    wire N__46414;
    wire N__46413;
    wire N__46412;
    wire N__46409;
    wire N__46406;
    wire N__46403;
    wire N__46398;
    wire N__46395;
    wire N__46392;
    wire N__46389;
    wire N__46382;
    wire N__46379;
    wire N__46376;
    wire N__46373;
    wire N__46368;
    wire N__46365;
    wire N__46362;
    wire N__46359;
    wire N__46354;
    wire N__46351;
    wire N__46348;
    wire N__46341;
    wire N__46334;
    wire N__46329;
    wire N__46328;
    wire N__46323;
    wire N__46322;
    wire N__46321;
    wire N__46320;
    wire N__46319;
    wire N__46316;
    wire N__46313;
    wire N__46308;
    wire N__46305;
    wire N__46302;
    wire N__46297;
    wire N__46296;
    wire N__46295;
    wire N__46294;
    wire N__46293;
    wire N__46292;
    wire N__46289;
    wire N__46286;
    wire N__46283;
    wire N__46272;
    wire N__46263;
    wire N__46260;
    wire N__46257;
    wire N__46254;
    wire N__46251;
    wire N__46250;
    wire N__46249;
    wire N__46248;
    wire N__46247;
    wire N__46246;
    wire N__46245;
    wire N__46244;
    wire N__46243;
    wire N__46240;
    wire N__46237;
    wire N__46234;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46217;
    wire N__46214;
    wire N__46211;
    wire N__46208;
    wire N__46207;
    wire N__46204;
    wire N__46201;
    wire N__46196;
    wire N__46193;
    wire N__46190;
    wire N__46185;
    wire N__46184;
    wire N__46181;
    wire N__46176;
    wire N__46173;
    wire N__46170;
    wire N__46165;
    wire N__46160;
    wire N__46157;
    wire N__46154;
    wire N__46151;
    wire N__46148;
    wire N__46141;
    wire N__46134;
    wire N__46133;
    wire N__46132;
    wire N__46129;
    wire N__46128;
    wire N__46125;
    wire N__46124;
    wire N__46123;
    wire N__46120;
    wire N__46119;
    wire N__46118;
    wire N__46115;
    wire N__46112;
    wire N__46105;
    wire N__46102;
    wire N__46097;
    wire N__46096;
    wire N__46093;
    wire N__46088;
    wire N__46085;
    wire N__46082;
    wire N__46079;
    wire N__46074;
    wire N__46069;
    wire N__46068;
    wire N__46067;
    wire N__46062;
    wire N__46059;
    wire N__46056;
    wire N__46053;
    wire N__46044;
    wire N__46043;
    wire N__46040;
    wire N__46037;
    wire N__46034;
    wire N__46031;
    wire N__46028;
    wire N__46025;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45990;
    wire N__45987;
    wire N__45984;
    wire N__45981;
    wire N__45978;
    wire N__45975;
    wire N__45972;
    wire N__45969;
    wire N__45966;
    wire N__45963;
    wire N__45960;
    wire N__45957;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45944;
    wire N__45943;
    wire N__45942;
    wire N__45939;
    wire N__45938;
    wire N__45935;
    wire N__45934;
    wire N__45933;
    wire N__45932;
    wire N__45931;
    wire N__45922;
    wire N__45919;
    wire N__45912;
    wire N__45911;
    wire N__45910;
    wire N__45909;
    wire N__45908;
    wire N__45905;
    wire N__45902;
    wire N__45897;
    wire N__45892;
    wire N__45891;
    wire N__45890;
    wire N__45889;
    wire N__45888;
    wire N__45887;
    wire N__45884;
    wire N__45883;
    wire N__45882;
    wire N__45881;
    wire N__45880;
    wire N__45879;
    wire N__45878;
    wire N__45877;
    wire N__45876;
    wire N__45875;
    wire N__45874;
    wire N__45873;
    wire N__45872;
    wire N__45871;
    wire N__45870;
    wire N__45869;
    wire N__45868;
    wire N__45867;
    wire N__45866;
    wire N__45865;
    wire N__45862;
    wire N__45861;
    wire N__45860;
    wire N__45859;
    wire N__45856;
    wire N__45849;
    wire N__45848;
    wire N__45847;
    wire N__45842;
    wire N__45841;
    wire N__45838;
    wire N__45829;
    wire N__45828;
    wire N__45825;
    wire N__45822;
    wire N__45817;
    wire N__45814;
    wire N__45809;
    wire N__45808;
    wire N__45807;
    wire N__45804;
    wire N__45803;
    wire N__45800;
    wire N__45799;
    wire N__45796;
    wire N__45793;
    wire N__45784;
    wire N__45783;
    wire N__45780;
    wire N__45777;
    wire N__45770;
    wire N__45765;
    wire N__45760;
    wire N__45755;
    wire N__45752;
    wire N__45751;
    wire N__45750;
    wire N__45747;
    wire N__45746;
    wire N__45741;
    wire N__45738;
    wire N__45737;
    wire N__45736;
    wire N__45735;
    wire N__45734;
    wire N__45731;
    wire N__45730;
    wire N__45729;
    wire N__45728;
    wire N__45723;
    wire N__45718;
    wire N__45717;
    wire N__45716;
    wire N__45713;
    wire N__45712;
    wire N__45711;
    wire N__45710;
    wire N__45709;
    wire N__45706;
    wire N__45701;
    wire N__45698;
    wire N__45695;
    wire N__45690;
    wire N__45687;
    wire N__45684;
    wire N__45681;
    wire N__45676;
    wire N__45667;
    wire N__45664;
    wire N__45661;
    wire N__45656;
    wire N__45651;
    wire N__45648;
    wire N__45645;
    wire N__45640;
    wire N__45639;
    wire N__45636;
    wire N__45629;
    wire N__45624;
    wire N__45621;
    wire N__45618;
    wire N__45611;
    wire N__45606;
    wire N__45603;
    wire N__45596;
    wire N__45591;
    wire N__45582;
    wire N__45567;
    wire N__45564;
    wire N__45557;
    wire N__45534;
    wire N__45533;
    wire N__45530;
    wire N__45529;
    wire N__45528;
    wire N__45527;
    wire N__45526;
    wire N__45525;
    wire N__45524;
    wire N__45523;
    wire N__45522;
    wire N__45521;
    wire N__45520;
    wire N__45519;
    wire N__45518;
    wire N__45515;
    wire N__45512;
    wire N__45507;
    wire N__45502;
    wire N__45501;
    wire N__45496;
    wire N__45495;
    wire N__45494;
    wire N__45493;
    wire N__45492;
    wire N__45491;
    wire N__45490;
    wire N__45487;
    wire N__45482;
    wire N__45481;
    wire N__45480;
    wire N__45477;
    wire N__45472;
    wire N__45465;
    wire N__45462;
    wire N__45459;
    wire N__45458;
    wire N__45457;
    wire N__45454;
    wire N__45449;
    wire N__45444;
    wire N__45441;
    wire N__45440;
    wire N__45439;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45425;
    wire N__45424;
    wire N__45423;
    wire N__45422;
    wire N__45421;
    wire N__45416;
    wire N__45415;
    wire N__45414;
    wire N__45411;
    wire N__45406;
    wire N__45401;
    wire N__45396;
    wire N__45393;
    wire N__45390;
    wire N__45387;
    wire N__45384;
    wire N__45381;
    wire N__45374;
    wire N__45373;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45361;
    wire N__45358;
    wire N__45353;
    wire N__45348;
    wire N__45341;
    wire N__45334;
    wire N__45329;
    wire N__45324;
    wire N__45303;
    wire N__45300;
    wire N__45297;
    wire N__45294;
    wire N__45291;
    wire N__45288;
    wire N__45285;
    wire N__45282;
    wire N__45279;
    wire N__45276;
    wire N__45273;
    wire N__45270;
    wire N__45267;
    wire N__45264;
    wire N__45261;
    wire N__45258;
    wire N__45255;
    wire N__45252;
    wire N__45249;
    wire N__45246;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45234;
    wire N__45231;
    wire N__45228;
    wire N__45225;
    wire N__45222;
    wire N__45219;
    wire N__45216;
    wire N__45213;
    wire N__45210;
    wire N__45207;
    wire N__45204;
    wire N__45201;
    wire N__45198;
    wire N__45195;
    wire N__45192;
    wire N__45189;
    wire N__45186;
    wire N__45183;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45171;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45153;
    wire N__45150;
    wire N__45147;
    wire N__45144;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45132;
    wire N__45129;
    wire N__45126;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45093;
    wire N__45090;
    wire N__45087;
    wire N__45084;
    wire N__45081;
    wire N__45078;
    wire N__45075;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45042;
    wire N__45039;
    wire N__45036;
    wire N__45033;
    wire N__45030;
    wire N__45027;
    wire N__45024;
    wire N__45021;
    wire N__45018;
    wire N__45015;
    wire N__45012;
    wire N__45009;
    wire N__45006;
    wire N__45003;
    wire N__45000;
    wire N__44997;
    wire N__44994;
    wire N__44993;
    wire N__44990;
    wire N__44987;
    wire N__44984;
    wire N__44981;
    wire N__44976;
    wire N__44973;
    wire N__44970;
    wire N__44967;
    wire N__44964;
    wire N__44961;
    wire N__44960;
    wire N__44959;
    wire N__44958;
    wire N__44957;
    wire N__44954;
    wire N__44953;
    wire N__44952;
    wire N__44949;
    wire N__44946;
    wire N__44943;
    wire N__44940;
    wire N__44935;
    wire N__44932;
    wire N__44931;
    wire N__44926;
    wire N__44923;
    wire N__44920;
    wire N__44915;
    wire N__44912;
    wire N__44909;
    wire N__44906;
    wire N__44901;
    wire N__44898;
    wire N__44897;
    wire N__44896;
    wire N__44893;
    wire N__44890;
    wire N__44885;
    wire N__44880;
    wire N__44871;
    wire N__44870;
    wire N__44869;
    wire N__44868;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44855;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44839;
    wire N__44836;
    wire N__44833;
    wire N__44832;
    wire N__44831;
    wire N__44828;
    wire N__44825;
    wire N__44822;
    wire N__44817;
    wire N__44808;
    wire N__44807;
    wire N__44804;
    wire N__44801;
    wire N__44798;
    wire N__44797;
    wire N__44794;
    wire N__44791;
    wire N__44788;
    wire N__44785;
    wire N__44782;
    wire N__44779;
    wire N__44778;
    wire N__44775;
    wire N__44770;
    wire N__44767;
    wire N__44762;
    wire N__44759;
    wire N__44754;
    wire N__44751;
    wire N__44750;
    wire N__44749;
    wire N__44746;
    wire N__44745;
    wire N__44742;
    wire N__44741;
    wire N__44738;
    wire N__44735;
    wire N__44732;
    wire N__44731;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44723;
    wire N__44722;
    wire N__44719;
    wire N__44718;
    wire N__44717;
    wire N__44716;
    wire N__44711;
    wire N__44706;
    wire N__44701;
    wire N__44698;
    wire N__44695;
    wire N__44694;
    wire N__44693;
    wire N__44690;
    wire N__44687;
    wire N__44682;
    wire N__44679;
    wire N__44674;
    wire N__44669;
    wire N__44664;
    wire N__44649;
    wire N__44646;
    wire N__44645;
    wire N__44644;
    wire N__44641;
    wire N__44638;
    wire N__44637;
    wire N__44636;
    wire N__44633;
    wire N__44628;
    wire N__44625;
    wire N__44622;
    wire N__44617;
    wire N__44614;
    wire N__44613;
    wire N__44610;
    wire N__44605;
    wire N__44602;
    wire N__44595;
    wire N__44594;
    wire N__44593;
    wire N__44592;
    wire N__44589;
    wire N__44588;
    wire N__44587;
    wire N__44586;
    wire N__44583;
    wire N__44580;
    wire N__44577;
    wire N__44572;
    wire N__44571;
    wire N__44568;
    wire N__44565;
    wire N__44560;
    wire N__44555;
    wire N__44554;
    wire N__44553;
    wire N__44550;
    wire N__44549;
    wire N__44546;
    wire N__44543;
    wire N__44540;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44528;
    wire N__44525;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44511;
    wire N__44508;
    wire N__44503;
    wire N__44500;
    wire N__44497;
    wire N__44492;
    wire N__44481;
    wire N__44478;
    wire N__44475;
    wire N__44472;
    wire N__44471;
    wire N__44470;
    wire N__44469;
    wire N__44466;
    wire N__44463;
    wire N__44460;
    wire N__44459;
    wire N__44456;
    wire N__44453;
    wire N__44446;
    wire N__44445;
    wire N__44444;
    wire N__44443;
    wire N__44440;
    wire N__44437;
    wire N__44434;
    wire N__44431;
    wire N__44430;
    wire N__44425;
    wire N__44422;
    wire N__44415;
    wire N__44412;
    wire N__44411;
    wire N__44410;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44390;
    wire N__44387;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44331;
    wire N__44328;
    wire N__44325;
    wire N__44322;
    wire N__44319;
    wire N__44316;
    wire N__44313;
    wire N__44310;
    wire N__44307;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44271;
    wire N__44268;
    wire N__44265;
    wire N__44262;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44229;
    wire N__44226;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44211;
    wire N__44208;
    wire N__44205;
    wire N__44202;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44190;
    wire N__44187;
    wire N__44184;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44166;
    wire N__44163;
    wire N__44160;
    wire N__44157;
    wire N__44154;
    wire N__44151;
    wire N__44148;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44126;
    wire N__44123;
    wire N__44122;
    wire N__44119;
    wire N__44116;
    wire N__44113;
    wire N__44110;
    wire N__44105;
    wire N__44102;
    wire N__44099;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44085;
    wire N__44082;
    wire N__44079;
    wire N__44076;
    wire N__44073;
    wire N__44070;
    wire N__44067;
    wire N__44064;
    wire N__44061;
    wire N__44058;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44043;
    wire N__44040;
    wire N__44037;
    wire N__44034;
    wire N__44031;
    wire N__44030;
    wire N__44029;
    wire N__44026;
    wire N__44023;
    wire N__44020;
    wire N__44017;
    wire N__44014;
    wire N__44011;
    wire N__44008;
    wire N__44003;
    wire N__43998;
    wire N__43995;
    wire N__43992;
    wire N__43989;
    wire N__43986;
    wire N__43983;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43971;
    wire N__43968;
    wire N__43965;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43953;
    wire N__43950;
    wire N__43947;
    wire N__43944;
    wire N__43941;
    wire N__43938;
    wire N__43935;
    wire N__43932;
    wire N__43929;
    wire N__43926;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43914;
    wire N__43911;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43868;
    wire N__43863;
    wire N__43862;
    wire N__43861;
    wire N__43860;
    wire N__43857;
    wire N__43856;
    wire N__43855;
    wire N__43848;
    wire N__43847;
    wire N__43846;
    wire N__43845;
    wire N__43844;
    wire N__43843;
    wire N__43840;
    wire N__43837;
    wire N__43834;
    wire N__43833;
    wire N__43832;
    wire N__43829;
    wire N__43824;
    wire N__43817;
    wire N__43812;
    wire N__43809;
    wire N__43806;
    wire N__43803;
    wire N__43800;
    wire N__43797;
    wire N__43792;
    wire N__43779;
    wire N__43776;
    wire N__43775;
    wire N__43772;
    wire N__43771;
    wire N__43768;
    wire N__43765;
    wire N__43762;
    wire N__43759;
    wire N__43754;
    wire N__43751;
    wire N__43748;
    wire N__43745;
    wire N__43740;
    wire N__43737;
    wire N__43734;
    wire N__43731;
    wire N__43728;
    wire N__43725;
    wire N__43722;
    wire N__43719;
    wire N__43716;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43695;
    wire N__43692;
    wire N__43689;
    wire N__43688;
    wire N__43687;
    wire N__43686;
    wire N__43683;
    wire N__43682;
    wire N__43679;
    wire N__43678;
    wire N__43675;
    wire N__43674;
    wire N__43673;
    wire N__43672;
    wire N__43671;
    wire N__43670;
    wire N__43669;
    wire N__43668;
    wire N__43667;
    wire N__43666;
    wire N__43665;
    wire N__43662;
    wire N__43659;
    wire N__43654;
    wire N__43647;
    wire N__43644;
    wire N__43641;
    wire N__43638;
    wire N__43637;
    wire N__43636;
    wire N__43635;
    wire N__43634;
    wire N__43633;
    wire N__43630;
    wire N__43629;
    wire N__43628;
    wire N__43625;
    wire N__43624;
    wire N__43623;
    wire N__43622;
    wire N__43621;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43611;
    wire N__43608;
    wire N__43607;
    wire N__43606;
    wire N__43603;
    wire N__43596;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43581;
    wire N__43580;
    wire N__43579;
    wire N__43578;
    wire N__43577;
    wire N__43576;
    wire N__43575;
    wire N__43572;
    wire N__43569;
    wire N__43566;
    wire N__43565;
    wire N__43564;
    wire N__43559;
    wire N__43556;
    wire N__43551;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43543;
    wire N__43542;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43528;
    wire N__43521;
    wire N__43520;
    wire N__43519;
    wire N__43518;
    wire N__43517;
    wire N__43516;
    wire N__43515;
    wire N__43514;
    wire N__43513;
    wire N__43508;
    wire N__43503;
    wire N__43502;
    wire N__43501;
    wire N__43500;
    wire N__43495;
    wire N__43492;
    wire N__43489;
    wire N__43480;
    wire N__43479;
    wire N__43476;
    wire N__43473;
    wire N__43468;
    wire N__43465;
    wire N__43462;
    wire N__43455;
    wire N__43452;
    wire N__43451;
    wire N__43450;
    wire N__43449;
    wire N__43448;
    wire N__43441;
    wire N__43434;
    wire N__43429;
    wire N__43426;
    wire N__43417;
    wire N__43408;
    wire N__43403;
    wire N__43396;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43376;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43356;
    wire N__43353;
    wire N__43344;
    wire N__43337;
    wire N__43334;
    wire N__43311;
    wire N__43308;
    wire N__43305;
    wire N__43302;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43287;
    wire N__43284;
    wire N__43283;
    wire N__43282;
    wire N__43281;
    wire N__43278;
    wire N__43273;
    wire N__43270;
    wire N__43269;
    wire N__43266;
    wire N__43261;
    wire N__43260;
    wire N__43257;
    wire N__43256;
    wire N__43255;
    wire N__43254;
    wire N__43249;
    wire N__43246;
    wire N__43243;
    wire N__43238;
    wire N__43235;
    wire N__43230;
    wire N__43227;
    wire N__43226;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43216;
    wire N__43213;
    wire N__43208;
    wire N__43205;
    wire N__43200;
    wire N__43191;
    wire N__43190;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43179;
    wire N__43178;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43168;
    wire N__43161;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43149;
    wire N__43146;
    wire N__43145;
    wire N__43144;
    wire N__43143;
    wire N__43142;
    wire N__43141;
    wire N__43140;
    wire N__43139;
    wire N__43138;
    wire N__43135;
    wire N__43130;
    wire N__43127;
    wire N__43120;
    wire N__43115;
    wire N__43108;
    wire N__43095;
    wire N__43092;
    wire N__43089;
    wire N__43086;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43078;
    wire N__43075;
    wire N__43072;
    wire N__43071;
    wire N__43068;
    wire N__43063;
    wire N__43060;
    wire N__43057;
    wire N__43054;
    wire N__43051;
    wire N__43048;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43032;
    wire N__43029;
    wire N__43026;
    wire N__43023;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43011;
    wire N__43008;
    wire N__43005;
    wire N__43002;
    wire N__42999;
    wire N__42996;
    wire N__42993;
    wire N__42992;
    wire N__42989;
    wire N__42986;
    wire N__42985;
    wire N__42984;
    wire N__42979;
    wire N__42978;
    wire N__42977;
    wire N__42974;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42961;
    wire N__42960;
    wire N__42957;
    wire N__42954;
    wire N__42951;
    wire N__42948;
    wire N__42945;
    wire N__42942;
    wire N__42939;
    wire N__42936;
    wire N__42933;
    wire N__42922;
    wire N__42919;
    wire N__42916;
    wire N__42913;
    wire N__42906;
    wire N__42903;
    wire N__42900;
    wire N__42897;
    wire N__42894;
    wire N__42891;
    wire N__42888;
    wire N__42885;
    wire N__42882;
    wire N__42879;
    wire N__42876;
    wire N__42873;
    wire N__42870;
    wire N__42867;
    wire N__42864;
    wire N__42861;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42834;
    wire N__42831;
    wire N__42828;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42816;
    wire N__42813;
    wire N__42810;
    wire N__42807;
    wire N__42804;
    wire N__42801;
    wire N__42798;
    wire N__42795;
    wire N__42792;
    wire N__42789;
    wire N__42786;
    wire N__42783;
    wire N__42780;
    wire N__42777;
    wire N__42774;
    wire N__42771;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42759;
    wire N__42756;
    wire N__42753;
    wire N__42750;
    wire N__42747;
    wire N__42744;
    wire N__42741;
    wire N__42738;
    wire N__42735;
    wire N__42732;
    wire N__42729;
    wire N__42726;
    wire N__42723;
    wire N__42720;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42708;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42696;
    wire N__42693;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42657;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42641;
    wire N__42640;
    wire N__42639;
    wire N__42638;
    wire N__42635;
    wire N__42632;
    wire N__42631;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42623;
    wire N__42620;
    wire N__42615;
    wire N__42614;
    wire N__42611;
    wire N__42610;
    wire N__42607;
    wire N__42604;
    wire N__42601;
    wire N__42598;
    wire N__42595;
    wire N__42592;
    wire N__42589;
    wire N__42586;
    wire N__42583;
    wire N__42576;
    wire N__42569;
    wire N__42566;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42533;
    wire N__42532;
    wire N__42531;
    wire N__42530;
    wire N__42529;
    wire N__42528;
    wire N__42527;
    wire N__42526;
    wire N__42525;
    wire N__42524;
    wire N__42523;
    wire N__42522;
    wire N__42519;
    wire N__42518;
    wire N__42517;
    wire N__42514;
    wire N__42511;
    wire N__42508;
    wire N__42505;
    wire N__42500;
    wire N__42497;
    wire N__42492;
    wire N__42489;
    wire N__42484;
    wire N__42483;
    wire N__42480;
    wire N__42479;
    wire N__42476;
    wire N__42473;
    wire N__42470;
    wire N__42467;
    wire N__42464;
    wire N__42461;
    wire N__42458;
    wire N__42451;
    wire N__42448;
    wire N__42447;
    wire N__42444;
    wire N__42441;
    wire N__42438;
    wire N__42429;
    wire N__42426;
    wire N__42417;
    wire N__42414;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42383;
    wire N__42382;
    wire N__42381;
    wire N__42380;
    wire N__42379;
    wire N__42378;
    wire N__42377;
    wire N__42376;
    wire N__42375;
    wire N__42374;
    wire N__42373;
    wire N__42370;
    wire N__42367;
    wire N__42366;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42351;
    wire N__42348;
    wire N__42345;
    wire N__42338;
    wire N__42333;
    wire N__42330;
    wire N__42325;
    wire N__42322;
    wire N__42315;
    wire N__42308;
    wire N__42305;
    wire N__42302;
    wire N__42299;
    wire N__42298;
    wire N__42295;
    wire N__42292;
    wire N__42289;
    wire N__42286;
    wire N__42283;
    wire N__42280;
    wire N__42277;
    wire N__42274;
    wire N__42269;
    wire N__42266;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42243;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42233;
    wire N__42232;
    wire N__42231;
    wire N__42230;
    wire N__42229;
    wire N__42228;
    wire N__42227;
    wire N__42226;
    wire N__42225;
    wire N__42224;
    wire N__42223;
    wire N__42222;
    wire N__42221;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42174;
    wire N__42171;
    wire N__42168;
    wire N__42165;
    wire N__42162;
    wire N__42159;
    wire N__42156;
    wire N__42153;
    wire N__42150;
    wire N__42147;
    wire N__42144;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42132;
    wire N__42129;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42117;
    wire N__42114;
    wire N__42113;
    wire N__42108;
    wire N__42105;
    wire N__42102;
    wire N__42099;
    wire N__42096;
    wire N__42093;
    wire N__42090;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42077;
    wire N__42074;
    wire N__42071;
    wire N__42066;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42051;
    wire N__42048;
    wire N__42047;
    wire N__42042;
    wire N__42039;
    wire N__42036;
    wire N__42033;
    wire N__42032;
    wire N__42031;
    wire N__42028;
    wire N__42025;
    wire N__42022;
    wire N__42015;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__42003;
    wire N__42000;
    wire N__41997;
    wire N__41994;
    wire N__41991;
    wire N__41988;
    wire N__41985;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41970;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41922;
    wire N__41919;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41898;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41871;
    wire N__41868;
    wire N__41867;
    wire N__41866;
    wire N__41863;
    wire N__41860;
    wire N__41857;
    wire N__41854;
    wire N__41851;
    wire N__41848;
    wire N__41845;
    wire N__41842;
    wire N__41839;
    wire N__41832;
    wire N__41829;
    wire N__41826;
    wire N__41823;
    wire N__41820;
    wire N__41817;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41805;
    wire N__41802;
    wire N__41799;
    wire N__41796;
    wire N__41793;
    wire N__41790;
    wire N__41787;
    wire N__41784;
    wire N__41781;
    wire N__41778;
    wire N__41777;
    wire N__41776;
    wire N__41773;
    wire N__41772;
    wire N__41769;
    wire N__41766;
    wire N__41763;
    wire N__41760;
    wire N__41757;
    wire N__41754;
    wire N__41751;
    wire N__41748;
    wire N__41745;
    wire N__41736;
    wire N__41733;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41723;
    wire N__41720;
    wire N__41717;
    wire N__41716;
    wire N__41713;
    wire N__41710;
    wire N__41707;
    wire N__41702;
    wire N__41699;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41676;
    wire N__41673;
    wire N__41670;
    wire N__41667;
    wire N__41664;
    wire N__41661;
    wire N__41658;
    wire N__41655;
    wire N__41652;
    wire N__41649;
    wire N__41646;
    wire N__41643;
    wire N__41640;
    wire N__41637;
    wire N__41634;
    wire N__41631;
    wire N__41628;
    wire N__41625;
    wire N__41622;
    wire N__41619;
    wire N__41616;
    wire N__41613;
    wire N__41610;
    wire N__41607;
    wire N__41604;
    wire N__41601;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41589;
    wire N__41586;
    wire N__41583;
    wire N__41580;
    wire N__41577;
    wire N__41574;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41562;
    wire N__41559;
    wire N__41556;
    wire N__41553;
    wire N__41550;
    wire N__41547;
    wire N__41544;
    wire N__41541;
    wire N__41538;
    wire N__41535;
    wire N__41532;
    wire N__41529;
    wire N__41526;
    wire N__41523;
    wire N__41520;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41508;
    wire N__41505;
    wire N__41502;
    wire N__41499;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41478;
    wire N__41475;
    wire N__41472;
    wire N__41469;
    wire N__41466;
    wire N__41463;
    wire N__41460;
    wire N__41457;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41439;
    wire N__41436;
    wire N__41433;
    wire N__41430;
    wire N__41427;
    wire N__41424;
    wire N__41421;
    wire N__41418;
    wire N__41415;
    wire N__41412;
    wire N__41409;
    wire N__41406;
    wire N__41403;
    wire N__41400;
    wire N__41397;
    wire N__41394;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41382;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41355;
    wire N__41352;
    wire N__41349;
    wire N__41346;
    wire N__41343;
    wire N__41340;
    wire N__41337;
    wire N__41334;
    wire N__41331;
    wire N__41328;
    wire N__41325;
    wire N__41322;
    wire N__41319;
    wire N__41316;
    wire N__41313;
    wire N__41310;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41283;
    wire N__41280;
    wire N__41277;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41247;
    wire N__41244;
    wire N__41241;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41229;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41217;
    wire N__41214;
    wire N__41211;
    wire N__41208;
    wire N__41205;
    wire N__41202;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41187;
    wire N__41184;
    wire N__41181;
    wire N__41178;
    wire N__41175;
    wire N__41172;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41157;
    wire N__41154;
    wire N__41151;
    wire N__41148;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41121;
    wire N__41118;
    wire N__41115;
    wire N__41112;
    wire N__41109;
    wire N__41106;
    wire N__41103;
    wire N__41100;
    wire N__41097;
    wire N__41094;
    wire N__41091;
    wire N__41088;
    wire N__41085;
    wire N__41082;
    wire N__41079;
    wire N__41076;
    wire N__41073;
    wire N__41070;
    wire N__41067;
    wire N__41064;
    wire N__41061;
    wire N__41058;
    wire N__41055;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41043;
    wire N__41040;
    wire N__41037;
    wire N__41034;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41016;
    wire N__41013;
    wire N__41010;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__40998;
    wire N__40995;
    wire N__40992;
    wire N__40989;
    wire N__40986;
    wire N__40983;
    wire N__40980;
    wire N__40977;
    wire N__40974;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40959;
    wire N__40956;
    wire N__40953;
    wire N__40950;
    wire N__40947;
    wire N__40944;
    wire N__40941;
    wire N__40938;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40926;
    wire N__40923;
    wire N__40920;
    wire N__40917;
    wire N__40914;
    wire N__40911;
    wire N__40908;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40893;
    wire N__40890;
    wire N__40887;
    wire N__40884;
    wire N__40881;
    wire N__40878;
    wire N__40875;
    wire N__40872;
    wire N__40869;
    wire N__40866;
    wire N__40863;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40845;
    wire N__40842;
    wire N__40839;
    wire N__40836;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40815;
    wire N__40812;
    wire N__40809;
    wire N__40806;
    wire N__40803;
    wire N__40800;
    wire N__40797;
    wire N__40794;
    wire N__40791;
    wire N__40788;
    wire N__40785;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40767;
    wire N__40764;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40752;
    wire N__40749;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40737;
    wire N__40734;
    wire N__40731;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40716;
    wire N__40713;
    wire N__40710;
    wire N__40707;
    wire N__40704;
    wire N__40701;
    wire N__40698;
    wire N__40695;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40683;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40665;
    wire N__40662;
    wire N__40659;
    wire N__40656;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40638;
    wire N__40637;
    wire N__40636;
    wire N__40635;
    wire N__40634;
    wire N__40633;
    wire N__40630;
    wire N__40619;
    wire N__40614;
    wire N__40613;
    wire N__40612;
    wire N__40611;
    wire N__40610;
    wire N__40609;
    wire N__40608;
    wire N__40605;
    wire N__40604;
    wire N__40603;
    wire N__40600;
    wire N__40587;
    wire N__40586;
    wire N__40585;
    wire N__40584;
    wire N__40583;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40575;
    wire N__40572;
    wire N__40569;
    wire N__40556;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40542;
    wire N__40541;
    wire N__40540;
    wire N__40539;
    wire N__40538;
    wire N__40535;
    wire N__40534;
    wire N__40533;
    wire N__40532;
    wire N__40531;
    wire N__40526;
    wire N__40523;
    wire N__40520;
    wire N__40519;
    wire N__40518;
    wire N__40517;
    wire N__40516;
    wire N__40513;
    wire N__40512;
    wire N__40511;
    wire N__40508;
    wire N__40505;
    wire N__40502;
    wire N__40499;
    wire N__40496;
    wire N__40495;
    wire N__40490;
    wire N__40485;
    wire N__40482;
    wire N__40479;
    wire N__40472;
    wire N__40465;
    wire N__40462;
    wire N__40459;
    wire N__40454;
    wire N__40449;
    wire N__40444;
    wire N__40441;
    wire N__40422;
    wire N__40419;
    wire N__40418;
    wire N__40417;
    wire N__40416;
    wire N__40413;
    wire N__40412;
    wire N__40409;
    wire N__40408;
    wire N__40407;
    wire N__40406;
    wire N__40403;
    wire N__40402;
    wire N__40401;
    wire N__40400;
    wire N__40399;
    wire N__40398;
    wire N__40397;
    wire N__40396;
    wire N__40395;
    wire N__40392;
    wire N__40379;
    wire N__40376;
    wire N__40367;
    wire N__40360;
    wire N__40359;
    wire N__40356;
    wire N__40355;
    wire N__40352;
    wire N__40349;
    wire N__40348;
    wire N__40347;
    wire N__40340;
    wire N__40337;
    wire N__40336;
    wire N__40335;
    wire N__40334;
    wire N__40333;
    wire N__40330;
    wire N__40329;
    wire N__40328;
    wire N__40327;
    wire N__40326;
    wire N__40325;
    wire N__40324;
    wire N__40323;
    wire N__40320;
    wire N__40315;
    wire N__40310;
    wire N__40307;
    wire N__40306;
    wire N__40305;
    wire N__40304;
    wire N__40301;
    wire N__40296;
    wire N__40291;
    wire N__40288;
    wire N__40283;
    wire N__40278;
    wire N__40269;
    wire N__40264;
    wire N__40261;
    wire N__40254;
    wire N__40251;
    wire N__40230;
    wire N__40227;
    wire N__40224;
    wire N__40221;
    wire N__40218;
    wire N__40215;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40173;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40158;
    wire N__40155;
    wire N__40152;
    wire N__40149;
    wire N__40146;
    wire N__40143;
    wire N__40140;
    wire N__40137;
    wire N__40134;
    wire N__40131;
    wire N__40128;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40098;
    wire N__40095;
    wire N__40092;
    wire N__40089;
    wire N__40088;
    wire N__40085;
    wire N__40082;
    wire N__40079;
    wire N__40076;
    wire N__40073;
    wire N__40068;
    wire N__40065;
    wire N__40062;
    wire N__40059;
    wire N__40056;
    wire N__40053;
    wire N__40050;
    wire N__40047;
    wire N__40044;
    wire N__40041;
    wire N__40038;
    wire N__40035;
    wire N__40032;
    wire N__40029;
    wire N__40026;
    wire N__40023;
    wire N__40020;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40005;
    wire N__40002;
    wire N__39999;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39978;
    wire N__39975;
    wire N__39972;
    wire N__39971;
    wire N__39968;
    wire N__39967;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39955;
    wire N__39954;
    wire N__39951;
    wire N__39948;
    wire N__39945;
    wire N__39942;
    wire N__39939;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39879;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39858;
    wire N__39855;
    wire N__39852;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39840;
    wire N__39837;
    wire N__39834;
    wire N__39831;
    wire N__39828;
    wire N__39825;
    wire N__39824;
    wire N__39821;
    wire N__39818;
    wire N__39817;
    wire N__39814;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39802;
    wire N__39799;
    wire N__39794;
    wire N__39791;
    wire N__39786;
    wire N__39783;
    wire N__39780;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39759;
    wire N__39756;
    wire N__39753;
    wire N__39750;
    wire N__39747;
    wire N__39744;
    wire N__39741;
    wire N__39738;
    wire N__39735;
    wire N__39732;
    wire N__39729;
    wire N__39726;
    wire N__39723;
    wire N__39720;
    wire N__39717;
    wire N__39714;
    wire N__39711;
    wire N__39708;
    wire N__39705;
    wire N__39702;
    wire N__39699;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39687;
    wire N__39684;
    wire N__39681;
    wire N__39678;
    wire N__39675;
    wire N__39672;
    wire N__39669;
    wire N__39666;
    wire N__39663;
    wire N__39660;
    wire N__39657;
    wire N__39654;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39636;
    wire N__39635;
    wire N__39632;
    wire N__39631;
    wire N__39628;
    wire N__39627;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39610;
    wire N__39607;
    wire N__39604;
    wire N__39597;
    wire N__39594;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39576;
    wire N__39573;
    wire N__39570;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39552;
    wire N__39549;
    wire N__39546;
    wire N__39543;
    wire N__39540;
    wire N__39537;
    wire N__39534;
    wire N__39531;
    wire N__39528;
    wire N__39525;
    wire N__39522;
    wire N__39519;
    wire N__39516;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39495;
    wire N__39492;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39477;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39453;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39438;
    wire N__39435;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39408;
    wire N__39405;
    wire N__39402;
    wire N__39399;
    wire N__39396;
    wire N__39393;
    wire N__39390;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39354;
    wire N__39351;
    wire N__39348;
    wire N__39345;
    wire N__39342;
    wire N__39341;
    wire N__39338;
    wire N__39335;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39321;
    wire N__39320;
    wire N__39315;
    wire N__39312;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39296;
    wire N__39293;
    wire N__39290;
    wire N__39287;
    wire N__39284;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39264;
    wire N__39263;
    wire N__39260;
    wire N__39257;
    wire N__39252;
    wire N__39249;
    wire N__39246;
    wire N__39243;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39207;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39135;
    wire N__39132;
    wire N__39129;
    wire N__39126;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39090;
    wire N__39087;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39075;
    wire N__39072;
    wire N__39069;
    wire N__39066;
    wire N__39063;
    wire N__39060;
    wire N__39057;
    wire N__39054;
    wire N__39051;
    wire N__39048;
    wire N__39045;
    wire N__39042;
    wire N__39039;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39024;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39012;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38964;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38910;
    wire N__38907;
    wire N__38904;
    wire N__38901;
    wire N__38898;
    wire N__38895;
    wire N__38892;
    wire N__38889;
    wire N__38886;
    wire N__38883;
    wire N__38880;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38778;
    wire N__38775;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38724;
    wire N__38721;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38594;
    wire N__38591;
    wire N__38588;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38576;
    wire N__38573;
    wire N__38570;
    wire N__38565;
    wire N__38564;
    wire N__38563;
    wire N__38558;
    wire N__38555;
    wire N__38554;
    wire N__38553;
    wire N__38552;
    wire N__38549;
    wire N__38546;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38528;
    wire N__38527;
    wire N__38526;
    wire N__38525;
    wire N__38522;
    wire N__38519;
    wire N__38512;
    wire N__38509;
    wire N__38506;
    wire N__38503;
    wire N__38496;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38481;
    wire N__38478;
    wire N__38475;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38454;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38442;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38397;
    wire N__38394;
    wire N__38391;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38361;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38343;
    wire N__38340;
    wire N__38337;
    wire N__38334;
    wire N__38331;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38295;
    wire N__38292;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38282;
    wire N__38279;
    wire N__38276;
    wire N__38273;
    wire N__38268;
    wire N__38267;
    wire N__38264;
    wire N__38261;
    wire N__38258;
    wire N__38253;
    wire N__38250;
    wire N__38247;
    wire N__38244;
    wire N__38241;
    wire N__38238;
    wire N__38235;
    wire N__38232;
    wire N__38229;
    wire N__38228;
    wire N__38227;
    wire N__38226;
    wire N__38225;
    wire N__38222;
    wire N__38213;
    wire N__38210;
    wire N__38207;
    wire N__38206;
    wire N__38205;
    wire N__38204;
    wire N__38203;
    wire N__38200;
    wire N__38197;
    wire N__38188;
    wire N__38185;
    wire N__38178;
    wire N__38175;
    wire N__38172;
    wire N__38169;
    wire N__38166;
    wire N__38163;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38148;
    wire N__38145;
    wire N__38142;
    wire N__38139;
    wire N__38136;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38121;
    wire N__38118;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38106;
    wire N__38103;
    wire N__38100;
    wire N__38097;
    wire N__38094;
    wire N__38091;
    wire N__38088;
    wire N__38085;
    wire N__38082;
    wire N__38081;
    wire N__38080;
    wire N__38079;
    wire N__38078;
    wire N__38077;
    wire N__38076;
    wire N__38075;
    wire N__38074;
    wire N__38073;
    wire N__38072;
    wire N__38071;
    wire N__38070;
    wire N__38069;
    wire N__38068;
    wire N__38065;
    wire N__38062;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38034;
    wire N__38033;
    wire N__38030;
    wire N__38027;
    wire N__38024;
    wire N__38021;
    wire N__38020;
    wire N__38019;
    wire N__38018;
    wire N__38009;
    wire N__38000;
    wire N__37991;
    wire N__37982;
    wire N__37977;
    wire N__37972;
    wire N__37971;
    wire N__37970;
    wire N__37969;
    wire N__37968;
    wire N__37967;
    wire N__37966;
    wire N__37965;
    wire N__37964;
    wire N__37959;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37945;
    wire N__37944;
    wire N__37941;
    wire N__37940;
    wire N__37937;
    wire N__37936;
    wire N__37933;
    wire N__37932;
    wire N__37931;
    wire N__37930;
    wire N__37929;
    wire N__37928;
    wire N__37925;
    wire N__37924;
    wire N__37921;
    wire N__37920;
    wire N__37917;
    wire N__37916;
    wire N__37913;
    wire N__37912;
    wire N__37911;
    wire N__37910;
    wire N__37909;
    wire N__37908;
    wire N__37907;
    wire N__37904;
    wire N__37903;
    wire N__37898;
    wire N__37895;
    wire N__37878;
    wire N__37875;
    wire N__37874;
    wire N__37873;
    wire N__37870;
    wire N__37869;
    wire N__37866;
    wire N__37865;
    wire N__37862;
    wire N__37845;
    wire N__37842;
    wire N__37841;
    wire N__37838;
    wire N__37837;
    wire N__37834;
    wire N__37833;
    wire N__37830;
    wire N__37829;
    wire N__37828;
    wire N__37825;
    wire N__37824;
    wire N__37821;
    wire N__37818;
    wire N__37811;
    wire N__37794;
    wire N__37791;
    wire N__37774;
    wire N__37767;
    wire N__37762;
    wire N__37757;
    wire N__37752;
    wire N__37749;
    wire N__37746;
    wire N__37743;
    wire N__37738;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37704;
    wire N__37701;
    wire N__37698;
    wire N__37695;
    wire N__37692;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37677;
    wire N__37674;
    wire N__37671;
    wire N__37668;
    wire N__37665;
    wire N__37662;
    wire N__37659;
    wire N__37656;
    wire N__37653;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37635;
    wire N__37632;
    wire N__37629;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37581;
    wire N__37578;
    wire N__37575;
    wire N__37572;
    wire N__37569;
    wire N__37566;
    wire N__37563;
    wire N__37560;
    wire N__37557;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37539;
    wire N__37536;
    wire N__37533;
    wire N__37530;
    wire N__37527;
    wire N__37524;
    wire N__37521;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37493;
    wire N__37492;
    wire N__37491;
    wire N__37490;
    wire N__37489;
    wire N__37476;
    wire N__37473;
    wire N__37470;
    wire N__37467;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37452;
    wire N__37449;
    wire N__37446;
    wire N__37443;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37410;
    wire N__37407;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37386;
    wire N__37383;
    wire N__37380;
    wire N__37377;
    wire N__37374;
    wire N__37371;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37353;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37332;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37305;
    wire N__37302;
    wire N__37299;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37251;
    wire N__37248;
    wire N__37245;
    wire N__37244;
    wire N__37241;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37228;
    wire N__37221;
    wire N__37220;
    wire N__37215;
    wire N__37212;
    wire N__37209;
    wire N__37208;
    wire N__37207;
    wire N__37204;
    wire N__37201;
    wire N__37198;
    wire N__37191;
    wire N__37188;
    wire N__37187;
    wire N__37186;
    wire N__37185;
    wire N__37182;
    wire N__37177;
    wire N__37174;
    wire N__37171;
    wire N__37164;
    wire N__37163;
    wire N__37162;
    wire N__37157;
    wire N__37154;
    wire N__37153;
    wire N__37148;
    wire N__37145;
    wire N__37140;
    wire N__37139;
    wire N__37138;
    wire N__37135;
    wire N__37132;
    wire N__37129;
    wire N__37122;
    wire N__37119;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37107;
    wire N__37104;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37092;
    wire N__37089;
    wire N__37088;
    wire N__37087;
    wire N__37084;
    wire N__37083;
    wire N__37080;
    wire N__37079;
    wire N__37076;
    wire N__37075;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37062;
    wire N__37059;
    wire N__37058;
    wire N__37055;
    wire N__37054;
    wire N__37053;
    wire N__37050;
    wire N__37047;
    wire N__37044;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37016;
    wire N__37009;
    wire N__37006;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36984;
    wire N__36981;
    wire N__36978;
    wire N__36975;
    wire N__36974;
    wire N__36973;
    wire N__36972;
    wire N__36969;
    wire N__36964;
    wire N__36961;
    wire N__36960;
    wire N__36959;
    wire N__36958;
    wire N__36957;
    wire N__36956;
    wire N__36955;
    wire N__36952;
    wire N__36949;
    wire N__36946;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36934;
    wire N__36931;
    wire N__36928;
    wire N__36925;
    wire N__36922;
    wire N__36917;
    wire N__36914;
    wire N__36911;
    wire N__36908;
    wire N__36901;
    wire N__36888;
    wire N__36885;
    wire N__36884;
    wire N__36883;
    wire N__36882;
    wire N__36879;
    wire N__36878;
    wire N__36877;
    wire N__36874;
    wire N__36873;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36860;
    wire N__36859;
    wire N__36856;
    wire N__36855;
    wire N__36852;
    wire N__36849;
    wire N__36848;
    wire N__36845;
    wire N__36844;
    wire N__36841;
    wire N__36840;
    wire N__36837;
    wire N__36832;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36819;
    wire N__36814;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36806;
    wire N__36805;
    wire N__36804;
    wire N__36801;
    wire N__36798;
    wire N__36795;
    wire N__36786;
    wire N__36783;
    wire N__36782;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36768;
    wire N__36763;
    wire N__36760;
    wire N__36753;
    wire N__36748;
    wire N__36745;
    wire N__36742;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36711;
    wire N__36708;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36693;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36681;
    wire N__36678;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36666;
    wire N__36663;
    wire N__36660;
    wire N__36659;
    wire N__36656;
    wire N__36655;
    wire N__36654;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36637;
    wire N__36634;
    wire N__36633;
    wire N__36630;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36620;
    wire N__36617;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36607;
    wire N__36604;
    wire N__36599;
    wire N__36596;
    wire N__36593;
    wire N__36590;
    wire N__36573;
    wire N__36570;
    wire N__36569;
    wire N__36566;
    wire N__36563;
    wire N__36558;
    wire N__36555;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36545;
    wire N__36542;
    wire N__36541;
    wire N__36538;
    wire N__36535;
    wire N__36532;
    wire N__36531;
    wire N__36530;
    wire N__36529;
    wire N__36526;
    wire N__36525;
    wire N__36522;
    wire N__36521;
    wire N__36518;
    wire N__36517;
    wire N__36514;
    wire N__36511;
    wire N__36508;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36498;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36472;
    wire N__36463;
    wire N__36458;
    wire N__36455;
    wire N__36444;
    wire N__36443;
    wire N__36442;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36431;
    wire N__36430;
    wire N__36427;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36406;
    wire N__36405;
    wire N__36402;
    wire N__36397;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36376;
    wire N__36373;
    wire N__36366;
    wire N__36361;
    wire N__36348;
    wire N__36347;
    wire N__36346;
    wire N__36345;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36333;
    wire N__36332;
    wire N__36329;
    wire N__36328;
    wire N__36327;
    wire N__36324;
    wire N__36323;
    wire N__36320;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36310;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36290;
    wire N__36287;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36271;
    wire N__36268;
    wire N__36255;
    wire N__36254;
    wire N__36253;
    wire N__36252;
    wire N__36251;
    wire N__36248;
    wire N__36247;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36232;
    wire N__36231;
    wire N__36230;
    wire N__36229;
    wire N__36228;
    wire N__36225;
    wire N__36220;
    wire N__36217;
    wire N__36214;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36191;
    wire N__36184;
    wire N__36171;
    wire N__36170;
    wire N__36169;
    wire N__36166;
    wire N__36163;
    wire N__36162;
    wire N__36159;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36148;
    wire N__36147;
    wire N__36146;
    wire N__36141;
    wire N__36138;
    wire N__36137;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36116;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36081;
    wire N__36080;
    wire N__36079;
    wire N__36076;
    wire N__36073;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36065;
    wire N__36064;
    wire N__36063;
    wire N__36060;
    wire N__36057;
    wire N__36054;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36029;
    wire N__36026;
    wire N__36023;
    wire N__36018;
    wire N__36013;
    wire N__36000;
    wire N__35997;
    wire N__35996;
    wire N__35995;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35981;
    wire N__35980;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35964;
    wire N__35961;
    wire N__35960;
    wire N__35957;
    wire N__35952;
    wire N__35951;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35932;
    wire N__35929;
    wire N__35926;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35912;
    wire N__35909;
    wire N__35906;
    wire N__35889;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35881;
    wire N__35878;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35870;
    wire N__35867;
    wire N__35864;
    wire N__35861;
    wire N__35858;
    wire N__35857;
    wire N__35854;
    wire N__35851;
    wire N__35850;
    wire N__35849;
    wire N__35846;
    wire N__35843;
    wire N__35842;
    wire N__35839;
    wire N__35836;
    wire N__35833;
    wire N__35830;
    wire N__35827;
    wire N__35824;
    wire N__35819;
    wire N__35816;
    wire N__35811;
    wire N__35808;
    wire N__35793;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35775;
    wire N__35772;
    wire N__35769;
    wire N__35768;
    wire N__35767;
    wire N__35764;
    wire N__35763;
    wire N__35762;
    wire N__35761;
    wire N__35758;
    wire N__35755;
    wire N__35752;
    wire N__35749;
    wire N__35746;
    wire N__35743;
    wire N__35740;
    wire N__35739;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35713;
    wire N__35708;
    wire N__35705;
    wire N__35698;
    wire N__35695;
    wire N__35682;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35669;
    wire N__35664;
    wire N__35661;
    wire N__35658;
    wire N__35655;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35647;
    wire N__35646;
    wire N__35643;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35633;
    wire N__35632;
    wire N__35631;
    wire N__35628;
    wire N__35627;
    wire N__35624;
    wire N__35621;
    wire N__35618;
    wire N__35617;
    wire N__35614;
    wire N__35609;
    wire N__35606;
    wire N__35603;
    wire N__35598;
    wire N__35595;
    wire N__35592;
    wire N__35589;
    wire N__35586;
    wire N__35571;
    wire N__35568;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35550;
    wire N__35547;
    wire N__35544;
    wire N__35541;
    wire N__35540;
    wire N__35537;
    wire N__35536;
    wire N__35533;
    wire N__35532;
    wire N__35529;
    wire N__35526;
    wire N__35523;
    wire N__35522;
    wire N__35521;
    wire N__35520;
    wire N__35517;
    wire N__35516;
    wire N__35511;
    wire N__35508;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35496;
    wire N__35493;
    wire N__35488;
    wire N__35485;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35463;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35436;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35418;
    wire N__35415;
    wire N__35414;
    wire N__35411;
    wire N__35410;
    wire N__35409;
    wire N__35406;
    wire N__35403;
    wire N__35400;
    wire N__35397;
    wire N__35396;
    wire N__35393;
    wire N__35388;
    wire N__35385;
    wire N__35384;
    wire N__35381;
    wire N__35380;
    wire N__35379;
    wire N__35376;
    wire N__35373;
    wire N__35370;
    wire N__35369;
    wire N__35366;
    wire N__35361;
    wire N__35358;
    wire N__35353;
    wire N__35350;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35328;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35316;
    wire N__35315;
    wire N__35312;
    wire N__35311;
    wire N__35310;
    wire N__35307;
    wire N__35306;
    wire N__35303;
    wire N__35302;
    wire N__35299;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35284;
    wire N__35281;
    wire N__35278;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35250;
    wire N__35235;
    wire N__35232;
    wire N__35231;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35219;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35204;
    wire N__35203;
    wire N__35202;
    wire N__35199;
    wire N__35196;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35188;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35165;
    wire N__35164;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35141;
    wire N__35136;
    wire N__35133;
    wire N__35128;
    wire N__35115;
    wire N__35112;
    wire N__35111;
    wire N__35108;
    wire N__35105;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35075;
    wire N__35072;
    wire N__35069;
    wire N__35064;
    wire N__35063;
    wire N__35062;
    wire N__35059;
    wire N__35058;
    wire N__35055;
    wire N__35052;
    wire N__35051;
    wire N__35050;
    wire N__35047;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35035;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35024;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__35003;
    wire N__35000;
    wire N__34997;
    wire N__34990;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34968;
    wire N__34965;
    wire N__34964;
    wire N__34961;
    wire N__34958;
    wire N__34957;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34949;
    wire N__34946;
    wire N__34943;
    wire N__34942;
    wire N__34941;
    wire N__34936;
    wire N__34933;
    wire N__34930;
    wire N__34929;
    wire N__34926;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34866;
    wire N__34863;
    wire N__34860;
    wire N__34857;
    wire N__34856;
    wire N__34853;
    wire N__34852;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34835;
    wire N__34834;
    wire N__34833;
    wire N__34828;
    wire N__34827;
    wire N__34824;
    wire N__34821;
    wire N__34818;
    wire N__34817;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34805;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34727;
    wire N__34726;
    wire N__34723;
    wire N__34720;
    wire N__34717;
    wire N__34714;
    wire N__34711;
    wire N__34710;
    wire N__34707;
    wire N__34706;
    wire N__34701;
    wire N__34700;
    wire N__34699;
    wire N__34696;
    wire N__34695;
    wire N__34692;
    wire N__34691;
    wire N__34688;
    wire N__34685;
    wire N__34682;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34629;
    wire N__34626;
    wire N__34623;
    wire N__34620;
    wire N__34619;
    wire N__34616;
    wire N__34613;
    wire N__34612;
    wire N__34609;
    wire N__34606;
    wire N__34605;
    wire N__34602;
    wire N__34601;
    wire N__34598;
    wire N__34595;
    wire N__34594;
    wire N__34591;
    wire N__34588;
    wire N__34585;
    wire N__34582;
    wire N__34579;
    wire N__34576;
    wire N__34575;
    wire N__34574;
    wire N__34571;
    wire N__34568;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34549;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34514;
    wire N__34511;
    wire N__34508;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34493;
    wire N__34490;
    wire N__34489;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34479;
    wire N__34476;
    wire N__34475;
    wire N__34472;
    wire N__34469;
    wire N__34466;
    wire N__34463;
    wire N__34460;
    wire N__34455;
    wire N__34454;
    wire N__34453;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34445;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34425;
    wire N__34422;
    wire N__34419;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34397;
    wire N__34394;
    wire N__34391;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34365;
    wire N__34364;
    wire N__34361;
    wire N__34358;
    wire N__34355;
    wire N__34350;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34319;
    wire N__34316;
    wire N__34313;
    wire N__34308;
    wire N__34305;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34290;
    wire N__34287;
    wire N__34284;
    wire N__34281;
    wire N__34278;
    wire N__34275;
    wire N__34274;
    wire N__34271;
    wire N__34268;
    wire N__34265;
    wire N__34260;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34250;
    wire N__34245;
    wire N__34244;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34230;
    wire N__34227;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34217;
    wire N__34214;
    wire N__34211;
    wire N__34208;
    wire N__34207;
    wire N__34202;
    wire N__34201;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34182;
    wire N__34179;
    wire N__34174;
    wire N__34161;
    wire N__34158;
    wire N__34155;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34101;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34074;
    wire N__34071;
    wire N__34068;
    wire N__34065;
    wire N__34062;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33947;
    wire N__33942;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33903;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33891;
    wire N__33890;
    wire N__33887;
    wire N__33884;
    wire N__33879;
    wire N__33876;
    wire N__33873;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33861;
    wire N__33858;
    wire N__33855;
    wire N__33852;
    wire N__33849;
    wire N__33848;
    wire N__33843;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33833;
    wire N__33830;
    wire N__33827;
    wire N__33822;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33779;
    wire N__33774;
    wire N__33771;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33753;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33723;
    wire N__33720;
    wire N__33717;
    wire N__33714;
    wire N__33711;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33699;
    wire N__33696;
    wire N__33693;
    wire N__33690;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33678;
    wire N__33675;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33657;
    wire N__33654;
    wire N__33651;
    wire N__33648;
    wire N__33645;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33609;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33566;
    wire N__33565;
    wire N__33564;
    wire N__33563;
    wire N__33562;
    wire N__33561;
    wire N__33560;
    wire N__33559;
    wire N__33558;
    wire N__33557;
    wire N__33556;
    wire N__33555;
    wire N__33554;
    wire N__33553;
    wire N__33552;
    wire N__33551;
    wire N__33550;
    wire N__33549;
    wire N__33548;
    wire N__33547;
    wire N__33546;
    wire N__33545;
    wire N__33544;
    wire N__33543;
    wire N__33542;
    wire N__33541;
    wire N__33532;
    wire N__33523;
    wire N__33514;
    wire N__33505;
    wire N__33504;
    wire N__33503;
    wire N__33494;
    wire N__33485;
    wire N__33484;
    wire N__33479;
    wire N__33476;
    wire N__33475;
    wire N__33470;
    wire N__33465;
    wire N__33460;
    wire N__33459;
    wire N__33458;
    wire N__33457;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33446;
    wire N__33445;
    wire N__33444;
    wire N__33443;
    wire N__33438;
    wire N__33435;
    wire N__33434;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33416;
    wire N__33409;
    wire N__33400;
    wire N__33395;
    wire N__33392;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33380;
    wire N__33375;
    wire N__33370;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33339;
    wire N__33330;
    wire N__33327;
    wire N__33324;
    wire N__33321;
    wire N__33320;
    wire N__33317;
    wire N__33314;
    wire N__33311;
    wire N__33306;
    wire N__33305;
    wire N__33304;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33287;
    wire N__33286;
    wire N__33285;
    wire N__33278;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33259;
    wire N__33256;
    wire N__33251;
    wire N__33248;
    wire N__33245;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33230;
    wire N__33225;
    wire N__33224;
    wire N__33223;
    wire N__33222;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33214;
    wire N__33213;
    wire N__33206;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33194;
    wire N__33191;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33177;
    wire N__33172;
    wire N__33169;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33150;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33129;
    wire N__33126;
    wire N__33123;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33050;
    wire N__33047;
    wire N__33044;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33029;
    wire N__33026;
    wire N__33023;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33009;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32987;
    wire N__32984;
    wire N__32981;
    wire N__32976;
    wire N__32973;
    wire N__32970;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32942;
    wire N__32939;
    wire N__32936;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32897;
    wire N__32894;
    wire N__32891;
    wire N__32886;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32862;
    wire N__32859;
    wire N__32856;
    wire N__32853;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32834;
    wire N__32831;
    wire N__32828;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32816;
    wire N__32813;
    wire N__32810;
    wire N__32805;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32795;
    wire N__32792;
    wire N__32789;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32772;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32736;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32691;
    wire N__32690;
    wire N__32689;
    wire N__32688;
    wire N__32687;
    wire N__32686;
    wire N__32685;
    wire N__32684;
    wire N__32683;
    wire N__32682;
    wire N__32681;
    wire N__32680;
    wire N__32679;
    wire N__32678;
    wire N__32677;
    wire N__32676;
    wire N__32675;
    wire N__32672;
    wire N__32665;
    wire N__32658;
    wire N__32649;
    wire N__32640;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32634;
    wire N__32633;
    wire N__32632;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32624;
    wire N__32623;
    wire N__32614;
    wire N__32611;
    wire N__32604;
    wire N__32599;
    wire N__32596;
    wire N__32595;
    wire N__32594;
    wire N__32591;
    wire N__32590;
    wire N__32587;
    wire N__32584;
    wire N__32583;
    wire N__32580;
    wire N__32569;
    wire N__32566;
    wire N__32563;
    wire N__32562;
    wire N__32559;
    wire N__32558;
    wire N__32555;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32547;
    wire N__32546;
    wire N__32543;
    wire N__32540;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32516;
    wire N__32515;
    wire N__32510;
    wire N__32507;
    wire N__32506;
    wire N__32505;
    wire N__32504;
    wire N__32503;
    wire N__32502;
    wire N__32501;
    wire N__32500;
    wire N__32499;
    wire N__32498;
    wire N__32497;
    wire N__32496;
    wire N__32495;
    wire N__32494;
    wire N__32493;
    wire N__32490;
    wire N__32487;
    wire N__32484;
    wire N__32479;
    wire N__32476;
    wire N__32471;
    wire N__32470;
    wire N__32469;
    wire N__32468;
    wire N__32467;
    wire N__32466;
    wire N__32463;
    wire N__32456;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32444;
    wire N__32441;
    wire N__32434;
    wire N__32423;
    wire N__32414;
    wire N__32413;
    wire N__32410;
    wire N__32407;
    wire N__32404;
    wire N__32399;
    wire N__32398;
    wire N__32391;
    wire N__32386;
    wire N__32383;
    wire N__32380;
    wire N__32377;
    wire N__32372;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32354;
    wire N__32353;
    wire N__32352;
    wire N__32351;
    wire N__32350;
    wire N__32347;
    wire N__32340;
    wire N__32337;
    wire N__32332;
    wire N__32327;
    wire N__32326;
    wire N__32323;
    wire N__32318;
    wire N__32309;
    wire N__32302;
    wire N__32299;
    wire N__32296;
    wire N__32293;
    wire N__32290;
    wire N__32287;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32254;
    wire N__32251;
    wire N__32246;
    wire N__32239;
    wire N__32236;
    wire N__32229;
    wire N__32228;
    wire N__32227;
    wire N__32226;
    wire N__32225;
    wire N__32224;
    wire N__32223;
    wire N__32222;
    wire N__32221;
    wire N__32220;
    wire N__32219;
    wire N__32218;
    wire N__32217;
    wire N__32216;
    wire N__32215;
    wire N__32214;
    wire N__32213;
    wire N__32212;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32198;
    wire N__32197;
    wire N__32196;
    wire N__32187;
    wire N__32186;
    wire N__32185;
    wire N__32184;
    wire N__32183;
    wire N__32182;
    wire N__32181;
    wire N__32180;
    wire N__32179;
    wire N__32178;
    wire N__32177;
    wire N__32176;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32165;
    wire N__32164;
    wire N__32163;
    wire N__32160;
    wire N__32159;
    wire N__32154;
    wire N__32153;
    wire N__32152;
    wire N__32151;
    wire N__32148;
    wire N__32141;
    wire N__32138;
    wire N__32123;
    wire N__32120;
    wire N__32103;
    wire N__32102;
    wire N__32099;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32077;
    wire N__32072;
    wire N__32069;
    wire N__32068;
    wire N__32067;
    wire N__32066;
    wire N__32063;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32042;
    wire N__32037;
    wire N__32032;
    wire N__32023;
    wire N__32016;
    wire N__32009;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31993;
    wire N__31980;
    wire N__31977;
    wire N__31974;
    wire N__31973;
    wire N__31970;
    wire N__31969;
    wire N__31968;
    wire N__31967;
    wire N__31966;
    wire N__31965;
    wire N__31964;
    wire N__31963;
    wire N__31962;
    wire N__31961;
    wire N__31960;
    wire N__31959;
    wire N__31958;
    wire N__31957;
    wire N__31956;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31948;
    wire N__31947;
    wire N__31946;
    wire N__31945;
    wire N__31944;
    wire N__31943;
    wire N__31942;
    wire N__31941;
    wire N__31940;
    wire N__31939;
    wire N__31938;
    wire N__31937;
    wire N__31936;
    wire N__31935;
    wire N__31934;
    wire N__31927;
    wire N__31922;
    wire N__31917;
    wire N__31916;
    wire N__31915;
    wire N__31914;
    wire N__31913;
    wire N__31912;
    wire N__31911;
    wire N__31910;
    wire N__31897;
    wire N__31892;
    wire N__31889;
    wire N__31886;
    wire N__31885;
    wire N__31884;
    wire N__31883;
    wire N__31882;
    wire N__31873;
    wire N__31866;
    wire N__31849;
    wire N__31848;
    wire N__31847;
    wire N__31840;
    wire N__31835;
    wire N__31824;
    wire N__31817;
    wire N__31814;
    wire N__31805;
    wire N__31798;
    wire N__31793;
    wire N__31788;
    wire N__31773;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31724;
    wire N__31721;
    wire N__31718;
    wire N__31713;
    wire N__31712;
    wire N__31711;
    wire N__31710;
    wire N__31709;
    wire N__31708;
    wire N__31707;
    wire N__31698;
    wire N__31697;
    wire N__31696;
    wire N__31695;
    wire N__31694;
    wire N__31693;
    wire N__31686;
    wire N__31685;
    wire N__31684;
    wire N__31683;
    wire N__31680;
    wire N__31671;
    wire N__31670;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31645;
    wire N__31642;
    wire N__31629;
    wire N__31626;
    wire N__31623;
    wire N__31620;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31590;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31485;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31434;
    wire N__31431;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31391;
    wire N__31390;
    wire N__31389;
    wire N__31388;
    wire N__31387;
    wire N__31380;
    wire N__31379;
    wire N__31376;
    wire N__31373;
    wire N__31370;
    wire N__31367;
    wire N__31364;
    wire N__31363;
    wire N__31360;
    wire N__31351;
    wire N__31350;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31326;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31305;
    wire N__31302;
    wire N__31301;
    wire N__31300;
    wire N__31299;
    wire N__31298;
    wire N__31297;
    wire N__31294;
    wire N__31293;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31280;
    wire N__31273;
    wire N__31270;
    wire N__31263;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31247;
    wire N__31242;
    wire N__31237;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31106;
    wire N__31105;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31094;
    wire N__31091;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31081;
    wire N__31078;
    wire N__31075;
    wire N__31074;
    wire N__31073;
    wire N__31072;
    wire N__31071;
    wire N__31070;
    wire N__31067;
    wire N__31064;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31048;
    wire N__31045;
    wire N__31040;
    wire N__31037;
    wire N__31020;
    wire N__31017;
    wire N__31016;
    wire N__31013;
    wire N__31010;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30992;
    wire N__30991;
    wire N__30988;
    wire N__30985;
    wire N__30982;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30947;
    wire N__30946;
    wire N__30943;
    wire N__30938;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30926;
    wire N__30923;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30911;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30897;
    wire N__30896;
    wire N__30893;
    wire N__30890;
    wire N__30887;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30873;
    wire N__30872;
    wire N__30871;
    wire N__30870;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30783;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30771;
    wire N__30770;
    wire N__30767;
    wire N__30764;
    wire N__30759;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30747;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30735;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30723;
    wire N__30722;
    wire N__30719;
    wire N__30716;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30704;
    wire N__30703;
    wire N__30702;
    wire N__30701;
    wire N__30700;
    wire N__30699;
    wire N__30698;
    wire N__30697;
    wire N__30678;
    wire N__30675;
    wire N__30672;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30603;
    wire N__30600;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30558;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30539;
    wire N__30536;
    wire N__30533;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30507;
    wire N__30504;
    wire N__30503;
    wire N__30500;
    wire N__30497;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30470;
    wire N__30467;
    wire N__30464;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30431;
    wire N__30428;
    wire N__30425;
    wire N__30420;
    wire N__30417;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30369;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30357;
    wire N__30354;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30339;
    wire N__30338;
    wire N__30335;
    wire N__30332;
    wire N__30327;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30306;
    wire N__30303;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30279;
    wire N__30276;
    wire N__30273;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30263;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30253;
    wire N__30248;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30096;
    wire N__30093;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30033;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30009;
    wire N__30006;
    wire N__30003;
    wire N__30000;
    wire N__29997;
    wire N__29994;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29943;
    wire N__29940;
    wire N__29939;
    wire N__29938;
    wire N__29937;
    wire N__29934;
    wire N__29933;
    wire N__29926;
    wire N__29925;
    wire N__29924;
    wire N__29923;
    wire N__29922;
    wire N__29921;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29898;
    wire N__29889;
    wire N__29886;
    wire N__29883;
    wire N__29880;
    wire N__29877;
    wire N__29874;
    wire N__29871;
    wire N__29870;
    wire N__29869;
    wire N__29868;
    wire N__29865;
    wire N__29864;
    wire N__29861;
    wire N__29860;
    wire N__29857;
    wire N__29856;
    wire N__29853;
    wire N__29852;
    wire N__29851;
    wire N__29838;
    wire N__29833;
    wire N__29830;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29751;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29699;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29376;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29346;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29192;
    wire N__29191;
    wire N__29190;
    wire N__29189;
    wire N__29188;
    wire N__29185;
    wire N__29180;
    wire N__29177;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29162;
    wire N__29159;
    wire N__29148;
    wire N__29145;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29133;
    wire N__29130;
    wire N__29129;
    wire N__29128;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29106;
    wire N__29105;
    wire N__29104;
    wire N__29103;
    wire N__29102;
    wire N__29101;
    wire N__29100;
    wire N__29099;
    wire N__29098;
    wire N__29097;
    wire N__29096;
    wire N__29095;
    wire N__29094;
    wire N__29093;
    wire N__29090;
    wire N__29085;
    wire N__29084;
    wire N__29073;
    wire N__29064;
    wire N__29061;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29051;
    wire N__29048;
    wire N__29045;
    wire N__29042;
    wire N__29041;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29024;
    wire N__29019;
    wire N__29014;
    wire N__29011;
    wire N__29006;
    wire N__29003;
    wire N__29000;
    wire N__28989;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28977;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28875;
    wire N__28872;
    wire N__28869;
    wire N__28866;
    wire N__28863;
    wire N__28860;
    wire N__28857;
    wire N__28854;
    wire N__28851;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28841;
    wire N__28838;
    wire N__28837;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28812;
    wire N__28809;
    wire N__28806;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28794;
    wire N__28793;
    wire N__28792;
    wire N__28789;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28704;
    wire N__28701;
    wire N__28698;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28674;
    wire N__28673;
    wire N__28670;
    wire N__28667;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28650;
    wire N__28647;
    wire N__28644;
    wire N__28641;
    wire N__28638;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28626;
    wire N__28623;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28499;
    wire N__28496;
    wire N__28493;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28451;
    wire N__28448;
    wire N__28445;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28404;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28353;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28242;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28109;
    wire N__28106;
    wire N__28103;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28067;
    wire N__28064;
    wire N__28061;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28034;
    wire N__28031;
    wire N__28028;
    wire N__28025;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27980;
    wire N__27979;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27966;
    wire N__27963;
    wire N__27960;
    wire N__27957;
    wire N__27956;
    wire N__27953;
    wire N__27948;
    wire N__27945;
    wire N__27942;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27912;
    wire N__27911;
    wire N__27908;
    wire N__27907;
    wire N__27904;
    wire N__27901;
    wire N__27898;
    wire N__27897;
    wire N__27894;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27882;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27865;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27807;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27777;
    wire N__27776;
    wire N__27773;
    wire N__27770;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27750;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27705;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27635;
    wire N__27632;
    wire N__27629;
    wire N__27626;
    wire N__27621;
    wire N__27618;
    wire N__27617;
    wire N__27616;
    wire N__27615;
    wire N__27612;
    wire N__27607;
    wire N__27606;
    wire N__27603;
    wire N__27602;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27583;
    wire N__27576;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27546;
    wire N__27543;
    wire N__27542;
    wire N__27541;
    wire N__27540;
    wire N__27537;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27527;
    wire N__27524;
    wire N__27521;
    wire N__27518;
    wire N__27515;
    wire N__27512;
    wire N__27505;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27491;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27470;
    wire N__27467;
    wire N__27464;
    wire N__27461;
    wire N__27456;
    wire N__27453;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27443;
    wire N__27438;
    wire N__27437;
    wire N__27434;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27396;
    wire N__27393;
    wire N__27392;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27378;
    wire N__27375;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27363;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27341;
    wire N__27336;
    wire N__27333;
    wire N__27332;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27314;
    wire N__27313;
    wire N__27312;
    wire N__27311;
    wire N__27306;
    wire N__27303;
    wire N__27298;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27045;
    wire N__27042;
    wire N__27041;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27002;
    wire N__27001;
    wire N__27000;
    wire N__26995;
    wire N__26994;
    wire N__26989;
    wire N__26986;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26966;
    wire N__26963;
    wire N__26958;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26852;
    wire N__26849;
    wire N__26846;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26828;
    wire N__26827;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26815;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26652;
    wire N__26649;
    wire N__26646;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26615;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26582;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26565;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26547;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26529;
    wire N__26528;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26516;
    wire N__26511;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26493;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26478;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26442;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26424;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26406;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26388;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26370;
    wire N__26367;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26349;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26331;
    wire N__26330;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26313;
    wire N__26310;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26299;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26287;
    wire N__26284;
    wire N__26281;
    wire N__26274;
    wire N__26271;
    wire N__26268;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26243;
    wire N__26242;
    wire N__26241;
    wire N__26240;
    wire N__26239;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26208;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26187;
    wire N__26184;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26169;
    wire N__26168;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26151;
    wire N__26150;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26120;
    wire N__26117;
    wire N__26116;
    wire N__26115;
    wire N__26112;
    wire N__26111;
    wire N__26108;
    wire N__26099;
    wire N__26094;
    wire N__26091;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26081;
    wire N__26080;
    wire N__26077;
    wire N__26076;
    wire N__26071;
    wire N__26066;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26042;
    wire N__26039;
    wire N__26038;
    wire N__26037;
    wire N__26036;
    wire N__26035;
    wire N__26026;
    wire N__26021;
    wire N__26016;
    wire N__26015;
    wire N__26014;
    wire N__26013;
    wire N__26012;
    wire N__26005;
    wire N__26000;
    wire N__25995;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25968;
    wire N__25965;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25932;
    wire N__25929;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25917;
    wire N__25914;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25902;
    wire N__25899;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25887;
    wire N__25884;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25869;
    wire N__25866;
    wire N__25865;
    wire N__25864;
    wire N__25863;
    wire N__25862;
    wire N__25861;
    wire N__25860;
    wire N__25859;
    wire N__25848;
    wire N__25841;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25829;
    wire N__25826;
    wire N__25823;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25796;
    wire N__25795;
    wire N__25792;
    wire N__25789;
    wire N__25786;
    wire N__25779;
    wire N__25778;
    wire N__25775;
    wire N__25774;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25761;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25710;
    wire N__25707;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25674;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25662;
    wire N__25661;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25647;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25635;
    wire N__25634;
    wire N__25631;
    wire N__25628;
    wire N__25623;
    wire N__25620;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25608;
    wire N__25605;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25590;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25578;
    wire N__25575;
    wire N__25574;
    wire N__25573;
    wire N__25570;
    wire N__25567;
    wire N__25564;
    wire N__25557;
    wire N__25556;
    wire N__25553;
    wire N__25552;
    wire N__25549;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25533;
    wire N__25532;
    wire N__25529;
    wire N__25526;
    wire N__25521;
    wire N__25518;
    wire N__25517;
    wire N__25516;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25488;
    wire N__25485;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25332;
    wire N__25329;
    wire N__25326;
    wire N__25323;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25311;
    wire N__25308;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25224;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25212;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25197;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25076;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25066;
    wire N__25061;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25022;
    wire N__25019;
    wire N__25016;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24954;
    wire N__24951;
    wire N__24948;
    wire N__24945;
    wire N__24944;
    wire N__24943;
    wire N__24942;
    wire N__24941;
    wire N__24940;
    wire N__24939;
    wire N__24938;
    wire N__24935;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24911;
    wire N__24910;
    wire N__24909;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24890;
    wire N__24879;
    wire N__24878;
    wire N__24875;
    wire N__24874;
    wire N__24871;
    wire N__24866;
    wire N__24859;
    wire N__24852;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24824;
    wire N__24823;
    wire N__24822;
    wire N__24819;
    wire N__24818;
    wire N__24817;
    wire N__24816;
    wire N__24811;
    wire N__24808;
    wire N__24805;
    wire N__24800;
    wire N__24799;
    wire N__24798;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24790;
    wire N__24787;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24768;
    wire N__24765;
    wire N__24758;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24719;
    wire N__24718;
    wire N__24715;
    wire N__24714;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24703;
    wire N__24700;
    wire N__24699;
    wire N__24698;
    wire N__24695;
    wire N__24694;
    wire N__24691;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24669;
    wire N__24664;
    wire N__24651;
    wire N__24648;
    wire N__24647;
    wire N__24646;
    wire N__24645;
    wire N__24642;
    wire N__24637;
    wire N__24634;
    wire N__24627;
    wire N__24626;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24614;
    wire N__24613;
    wire N__24612;
    wire N__24611;
    wire N__24610;
    wire N__24603;
    wire N__24602;
    wire N__24599;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24525;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24509;
    wire N__24508;
    wire N__24507;
    wire N__24506;
    wire N__24503;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24491;
    wire N__24490;
    wire N__24489;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24477;
    wire N__24470;
    wire N__24469;
    wire N__24468;
    wire N__24467;
    wire N__24466;
    wire N__24465;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24451;
    wire N__24438;
    wire N__24429;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24380;
    wire N__24379;
    wire N__24378;
    wire N__24377;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24365;
    wire N__24362;
    wire N__24361;
    wire N__24358;
    wire N__24357;
    wire N__24352;
    wire N__24347;
    wire N__24344;
    wire N__24339;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24314;
    wire N__24311;
    wire N__24310;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24277;
    wire N__24274;
    wire N__24273;
    wire N__24272;
    wire N__24265;
    wire N__24260;
    wire N__24259;
    wire N__24258;
    wire N__24257;
    wire N__24252;
    wire N__24247;
    wire N__24244;
    wire N__24241;
    wire N__24236;
    wire N__24231;
    wire N__24230;
    wire N__24229;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24204;
    wire N__24203;
    wire N__24202;
    wire N__24201;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24189;
    wire N__24186;
    wire N__24177;
    wire N__24176;
    wire N__24173;
    wire N__24168;
    wire N__24165;
    wire N__24164;
    wire N__24163;
    wire N__24160;
    wire N__24155;
    wire N__24152;
    wire N__24147;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24065;
    wire N__24060;
    wire N__24059;
    wire N__24058;
    wire N__24057;
    wire N__24056;
    wire N__24053;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24041;
    wire N__24040;
    wire N__24033;
    wire N__24028;
    wire N__24025;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23987;
    wire N__23984;
    wire N__23979;
    wire N__23978;
    wire N__23973;
    wire N__23972;
    wire N__23971;
    wire N__23970;
    wire N__23967;
    wire N__23966;
    wire N__23965;
    wire N__23964;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23948;
    wire N__23945;
    wire N__23940;
    wire N__23935;
    wire N__23932;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23910;
    wire N__23907;
    wire N__23906;
    wire N__23903;
    wire N__23902;
    wire N__23901;
    wire N__23900;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23892;
    wire N__23887;
    wire N__23884;
    wire N__23879;
    wire N__23878;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23864;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23848;
    wire N__23845;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23829;
    wire N__23826;
    wire N__23823;
    wire N__23820;
    wire N__23819;
    wire N__23818;
    wire N__23811;
    wire N__23808;
    wire N__23807;
    wire N__23802;
    wire N__23799;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23789;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23763;
    wire N__23760;
    wire N__23757;
    wire N__23756;
    wire N__23751;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23739;
    wire N__23736;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23728;
    wire N__23727;
    wire N__23726;
    wire N__23721;
    wire N__23718;
    wire N__23717;
    wire N__23712;
    wire N__23709;
    wire N__23704;
    wire N__23697;
    wire N__23694;
    wire N__23693;
    wire N__23692;
    wire N__23689;
    wire N__23688;
    wire N__23683;
    wire N__23682;
    wire N__23679;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23642;
    wire N__23641;
    wire N__23636;
    wire N__23633;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23507;
    wire N__23502;
    wire N__23499;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23487;
    wire N__23484;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23472;
    wire N__23469;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23457;
    wire N__23454;
    wire N__23451;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23430;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23355;
    wire N__23352;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23340;
    wire N__23337;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23325;
    wire N__23322;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23307;
    wire N__23304;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23292;
    wire N__23289;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23277;
    wire N__23274;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23262;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23246;
    wire N__23245;
    wire N__23244;
    wire N__23243;
    wire N__23242;
    wire N__23241;
    wire N__23240;
    wire N__23231;
    wire N__23230;
    wire N__23229;
    wire N__23228;
    wire N__23227;
    wire N__23226;
    wire N__23225;
    wire N__23224;
    wire N__23223;
    wire N__23222;
    wire N__23221;
    wire N__23220;
    wire N__23219;
    wire N__23218;
    wire N__23217;
    wire N__23216;
    wire N__23215;
    wire N__23206;
    wire N__23203;
    wire N__23194;
    wire N__23185;
    wire N__23176;
    wire N__23167;
    wire N__23154;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23136;
    wire N__23133;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23121;
    wire N__23118;
    wire N__23115;
    wire N__23112;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23085;
    wire N__23082;
    wire N__23079;
    wire N__23076;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22989;
    wire N__22986;
    wire N__22983;
    wire N__22980;
    wire N__22977;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22640;
    wire N__22639;
    wire N__22638;
    wire N__22637;
    wire N__22636;
    wire N__22631;
    wire N__22630;
    wire N__22629;
    wire N__22628;
    wire N__22627;
    wire N__22624;
    wire N__22619;
    wire N__22618;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22606;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22590;
    wire N__22587;
    wire N__22576;
    wire N__22569;
    wire N__22566;
    wire N__22563;
    wire N__22560;
    wire N__22557;
    wire N__22556;
    wire N__22555;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22532;
    wire N__22531;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22494;
    wire N__22493;
    wire N__22492;
    wire N__22487;
    wire N__22484;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22469;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22379;
    wire N__22378;
    wire N__22377;
    wire N__22376;
    wire N__22375;
    wire N__22374;
    wire N__22373;
    wire N__22364;
    wire N__22355;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22289;
    wire N__22284;
    wire N__22281;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22170;
    wire N__22167;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22022;
    wire N__22019;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22007;
    wire N__22004;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21965;
    wire N__21964;
    wire N__21961;
    wire N__21956;
    wire N__21951;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21701;
    wire N__21700;
    wire N__21697;
    wire N__21696;
    wire N__21695;
    wire N__21694;
    wire N__21693;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21662;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21641;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21624;
    wire N__21623;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21606;
    wire N__21605;
    wire N__21602;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21585;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21573;
    wire N__21570;
    wire N__21569;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21540;
    wire N__21537;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21525;
    wire N__21524;
    wire N__21521;
    wire N__21520;
    wire N__21517;
    wire N__21512;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21489;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21470;
    wire N__21465;
    wire N__21462;
    wire N__21461;
    wire N__21460;
    wire N__21459;
    wire N__21458;
    wire N__21457;
    wire N__21456;
    wire N__21455;
    wire N__21444;
    wire N__21437;
    wire N__21432;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21422;
    wire N__21417;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21409;
    wire N__21408;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21314;
    wire N__21309;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21299;
    wire N__21298;
    wire N__21297;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21278;
    wire N__21275;
    wire N__21272;
    wire N__21265;
    wire N__21262;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21219;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21207;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21192;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21180;
    wire N__21177;
    wire N__21176;
    wire N__21173;
    wire N__21172;
    wire N__21169;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21110;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21086;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21029;
    wire N__21028;
    wire N__21027;
    wire N__21026;
    wire N__21023;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21007;
    wire N__21000;
    wire N__20999;
    wire N__20996;
    wire N__20995;
    wire N__20994;
    wire N__20987;
    wire N__20986;
    wire N__20985;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20864;
    wire N__20863;
    wire N__20860;
    wire N__20857;
    wire N__20854;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20840;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20813;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20796;
    wire N__20793;
    wire N__20792;
    wire N__20791;
    wire N__20790;
    wire N__20789;
    wire N__20788;
    wire N__20787;
    wire N__20786;
    wire N__20779;
    wire N__20774;
    wire N__20767;
    wire N__20760;
    wire N__20757;
    wire N__20756;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20736;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20702;
    wire N__20701;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20627;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20613;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20559;
    wire N__20556;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20544;
    wire N__20541;
    wire N__20538;
    wire N__20535;
    wire N__20532;
    wire N__20529;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire clk_c;
    wire \pll128M2_inst.pll_clk64_0 ;
    wire \pll128M2_inst.pll_clk128 ;
    wire VCCG0;
    wire button_mode_c;
    wire button_mode_ibuf_RNIN5KZ0Z7;
    wire DAC_cs_c;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1 ;
    wire \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i ;
    wire \spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i_cascade_ ;
    wire bfn_2_11_0_;
    wire sRAM_pointer_read_cry_0;
    wire sRAM_pointer_read_cry_1;
    wire sRAM_pointer_read_cry_2;
    wire sRAM_pointer_read_cry_3;
    wire sRAM_pointer_read_cry_4;
    wire sRAM_pointer_read_cry_5;
    wire sRAM_pointer_read_cry_6;
    wire sRAM_pointer_read_cry_7;
    wire bfn_2_12_0_;
    wire sRAM_pointer_read_cry_8;
    wire sRAM_pointer_read_cry_9;
    wire sRAM_pointer_read_cry_10;
    wire sRAM_pointer_read_cry_11;
    wire sRAM_pointer_read_cry_12;
    wire sRAM_pointer_read_cry_13;
    wire sRAM_pointer_read_cry_14;
    wire sRAM_pointer_read_cry_15;
    wire bfn_2_13_0_;
    wire sRAM_pointer_read_cry_16;
    wire sRAM_pointer_read_cry_17;
    wire N_28_g;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_s_0 ;
    wire bfn_3_3_0_;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_s_1 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2 ;
    wire bfn_3_4_0_;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0 ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1 ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4 ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3 ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4 ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO ;
    wire bfn_3_5_0_;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0 ;
    wire DAC_mosi_c;
    wire \spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4 ;
    wire DAC_sclk_c;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6 ;
    wire \spi_master_inst.o_sclk_RNIH6AC ;
    wire \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO ;
    wire bfn_5_5_0_;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_0 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_1 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_2 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_3 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_4 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_5 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_i_cry_6 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4 ;
    wire \spi_master_inst.sclk_gen_u0.N_1666_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4 ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0 ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.N_48_cascade_ ;
    wire \spi_master_inst.ss_start_i ;
    wire sEEPonPoff_i_0;
    wire bfn_5_10_0_;
    wire sEEPonPoff_i_1;
    wire un4_spoff_cry_0;
    wire sEEPonPoff_i_2;
    wire un4_spoff_cry_1;
    wire sEEPonPoff_i_3;
    wire un4_spoff_cry_2;
    wire sEEPonPoff_i_4;
    wire un4_spoff_cry_3;
    wire sEEPonPoff_i_5;
    wire un4_spoff_cry_4;
    wire sEEPonPoff_i_6;
    wire un4_spoff_cry_5;
    wire sEEPonPoff_i_7;
    wire un4_spoff_cry_6;
    wire un4_spoff_cry_7;
    wire bfn_5_11_0_;
    wire un4_spoff_cry_8;
    wire un4_spoff_cry_9;
    wire un4_spoff_cry_10;
    wire un4_spoff_cry_11;
    wire un4_spoff_cry_12;
    wire un4_spoff_cry_13;
    wire un4_spoff_cry_14;
    wire un4_spoff_cry_15;
    wire bfn_5_12_0_;
    wire un4_spoff_cry_16;
    wire un4_spoff_cry_17;
    wire un4_spoff_cry_18;
    wire un4_spoff_cry_19;
    wire un4_spoff_cry_20;
    wire un4_spoff_cry_21;
    wire un4_spoff_cry_22;
    wire un4_spoff_cry_23;
    wire bfn_5_13_0_;
    wire \spi_master_inst.spi_data_path_u1.N_1423 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1 ;
    wire \spi_master_inst.spi_data_path_u1.N_1416 ;
    wire \spi_master_inst.spi_data_path_u1.N_1415 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14_cascade_ ;
    wire \spi_master_inst.spi_data_path_u1.N_1419 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_ ;
    wire \spi_master_inst.spi_data_path_u1.N_1422 ;
    wire \spi_master_inst.sclk_gen_u0.N_1520 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_start_i_i ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15_cascade_ ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ;
    wire \spi_master_inst.spi_data_path_u1.N_1412 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1 ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2 ;
    wire \spi_master_inst.sclk_gen_u0.N_1666 ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0 ;
    wire \spi_master_inst.sclk_gen_u0.N_1515_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.N_36_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.N_48 ;
    wire \spi_master_inst.sclk_gen_u0.N_5_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.delay_count_start_iZ0 ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1 ;
    wire sEEPonPoffZ0Z_0;
    wire sEEPonPoffZ0Z_1;
    wire sEEPonPoffZ0Z_2;
    wire sEEPonPoffZ0Z_3;
    wire sEEPonPoffZ0Z_4;
    wire sEEPonPoffZ0Z_5;
    wire sEEPonPoffZ0Z_6;
    wire sEEPonPoffZ0Z_7;
    wire sEEPonZ0Z_0;
    wire sEEPon_i_0;
    wire bfn_6_11_0_;
    wire sEEPonZ0Z_1;
    wire sEEPon_i_1;
    wire un7_spon_cry_0;
    wire sEEPonZ0Z_2;
    wire sEEPon_i_2;
    wire un7_spon_cry_1;
    wire sEEPonZ0Z_3;
    wire sEEPon_i_3;
    wire un7_spon_cry_2;
    wire sEEPonZ0Z_4;
    wire sEEPon_i_4;
    wire un7_spon_cry_3;
    wire sEEPonZ0Z_5;
    wire sEEPon_i_5;
    wire un7_spon_cry_4;
    wire sEEPonZ0Z_6;
    wire sEEPon_i_6;
    wire un7_spon_cry_5;
    wire sEEPonZ0Z_7;
    wire sEEPon_i_7;
    wire un7_spon_cry_6;
    wire un7_spon_cry_7;
    wire bfn_6_12_0_;
    wire un7_spon_cry_8;
    wire un7_spon_cry_9;
    wire un7_spon_cry_10;
    wire un7_spon_cry_11;
    wire un7_spon_cry_12;
    wire un7_spon_cry_13;
    wire un7_spon_cry_14;
    wire un7_spon_cry_15;
    wire bfn_6_13_0_;
    wire un7_spon_cry_16;
    wire un7_spon_cry_17;
    wire un7_spon_cry_18;
    wire un7_spon_cry_19;
    wire un7_spon_cry_20;
    wire un7_spon_cry_21;
    wire un7_spon_cry_22;
    wire un7_spon_cry_23;
    wire bfn_6_14_0_;
    wire pon_obuf_RNOZ0;
    wire g1_0_5;
    wire g1;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1 ;
    wire sEESingleContZ0;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3 ;
    wire \spi_master_inst.sclk_gen_u0.N_1515 ;
    wire sEESingleCont_1_sqmuxa;
    wire un3_trig_0_2;
    wire un3_trig_0_1;
    wire g1_3_cascade_;
    wire sEETrigInternal_prev_RNISEUGZ0_cascade_;
    wire sTrigInternal_RNIOMLDZ0Z1_cascade_;
    wire sTrigInternal_RNIOMLDZ0Z1;
    wire sTrigInternal_RNOZ0Z_0_cascade_;
    wire un3_trig_0;
    wire un3_trig_0_4;
    wire un1_reset_rpi_inv_2_i_o3_8;
    wire un1_reset_rpi_inv_2_i_o3_18_cascade_;
    wire un3_trig_0_5;
    wire un1_reset_rpi_inv_2_i_o3_13;
    wire g0_2_0_3;
    wire sbuttonModeStatus_0_sqmuxa_22_cascade_;
    wire sbuttonModeStatusZ0;
    wire g1_0_0_3;
    wire un1_reset_rpi_inv_2_i_o3_16;
    wire g0_2_0_4;
    wire g2_0_4;
    wire g2_0_3;
    wire g1_0_1_1_cascade_;
    wire g1_0_4;
    wire op_gt_op_gt_un13_striginternallto23_13;
    wire op_gt_op_gt_un13_striginternal_0_cascade_;
    wire op_gt_op_gt_un13_striginternallto23_11_cascade_;
    wire op_gt_op_gt_un13_striginternallto23_16;
    wire sTrigInternalZ0;
    wire op_gt_op_gt_un13_striginternal_0;
    wire LED_ACQ_obuf_RNOZ0;
    wire op_gt_op_gt_un13_striginternallto23_18;
    wire bfn_7_16_0_;
    wire sCounterRAM_cry_0;
    wire sCounterRAM_cry_1;
    wire sCounterRAM_cry_2;
    wire sCounterRAM_cry_3;
    wire sCounterRAM_cry_4;
    wire sCounterRAM_cry_5;
    wire un1_spi_data_miso_0_sqmuxa_1_i_0_N_3_0;
    wire sCounterRAM_cry_6;
    wire sSPI_MSB0LSB1_RNIO3VPZ0Z1;
    wire sbuttonModeStatus_0_sqmuxa_16;
    wire sbuttonModeStatus_0_sqmuxa_14;
    wire sbuttonModeStatus_0_sqmuxa_15;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10 ;
    wire \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12 ;
    wire \spi_master_inst.sclk_gen_u0.N_150_0 ;
    wire \spi_master_inst.sclk_gen_u0.N_36 ;
    wire \spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0 ;
    wire \spi_master_inst.sclk_gen_u0.div_clk_iZ0 ;
    wire \spi_master_inst.sclk_gen_u0.delay_clk_iZ0 ;
    wire g0_2_0_2;
    wire g1_1;
    wire g2_0_2_cascade_;
    wire g1_0_3;
    wire g0_2_0_1;
    wire g2_0_1_cascade_;
    wire g1_2;
    wire g1_0_0_1;
    wire g1_0_2;
    wire g0_2_0_0;
    wire g2_0_0_cascade_;
    wire g1_0_0_0;
    wire g1_0_1;
    wire g0_2_0;
    wire g1_4;
    wire g2_0_cascade_;
    wire sEEPeriodZ0Z_0;
    wire sEEPeriod_i_0;
    wire bfn_8_10_0_;
    wire sEEPeriodZ0Z_1;
    wire sEEPeriod_i_1;
    wire un4_speriod_cry_0;
    wire sEEPeriodZ0Z_2;
    wire sEEPeriod_i_2;
    wire un4_speriod_cry_1;
    wire sEEPeriodZ0Z_3;
    wire sEEPeriod_i_3;
    wire un4_speriod_cry_2;
    wire sEEPeriodZ0Z_4;
    wire sEEPeriod_i_4;
    wire un4_speriod_cry_3;
    wire sEEPeriodZ0Z_5;
    wire sEEPeriod_i_5;
    wire un4_speriod_cry_4;
    wire sEEPeriodZ0Z_6;
    wire sEEPeriod_i_6;
    wire un4_speriod_cry_5;
    wire sEEPeriodZ0Z_7;
    wire sEEPeriod_i_7;
    wire un4_speriod_cry_6;
    wire un4_speriod_cry_7;
    wire sEEPeriod_i_8;
    wire bfn_8_11_0_;
    wire sEEPeriod_i_9;
    wire un4_speriod_cry_8;
    wire sEEPeriod_i_10;
    wire un4_speriod_cry_9;
    wire sEEPeriod_i_11;
    wire un4_speriod_cry_10;
    wire sEEPeriod_i_12;
    wire un4_speriod_cry_11;
    wire sEEPeriod_i_13;
    wire un4_speriod_cry_12;
    wire sEEPeriod_i_14;
    wire un4_speriod_cry_13;
    wire sEEPeriod_i_15;
    wire un4_speriod_cry_14;
    wire un4_speriod_cry_15;
    wire sEEPeriodZ0Z_16;
    wire sEEPeriod_i_16;
    wire bfn_8_12_0_;
    wire sEEPeriodZ0Z_17;
    wire sEEPeriod_i_17;
    wire un4_speriod_cry_16;
    wire sEEPeriodZ0Z_18;
    wire sEEPeriod_i_18;
    wire un4_speriod_cry_17;
    wire sEEPeriodZ0Z_19;
    wire sEEPeriod_i_19;
    wire un4_speriod_cry_18;
    wire sEEPeriodZ0Z_20;
    wire sEEPeriod_i_20;
    wire un4_speriod_cry_19;
    wire sEEPeriodZ0Z_21;
    wire sEEPeriod_i_21;
    wire un4_speriod_cry_20;
    wire sEEPeriodZ0Z_22;
    wire sEEPeriod_i_22;
    wire un4_speriod_cry_21;
    wire sEEPeriodZ0Z_23;
    wire sEEPeriod_i_23;
    wire un4_speriod_cry_22;
    wire un4_speriod_cry_23;
    wire bfn_8_13_0_;
    wire un1_reset_rpi_inv_2_i_o3_15;
    wire un1_reset_rpi_inv_2_i_o3_11;
    wire sbuttonModeStatus_0_sqmuxa_17;
    wire bfn_8_14_0_;
    wire sCounter_cry_0;
    wire sCounter_cry_1;
    wire sCounter_cry_2;
    wire sCounter_cry_3;
    wire sCounter_cry_4;
    wire sCounter_cry_5;
    wire sCounter_cry_6;
    wire sCounter_cry_7;
    wire bfn_8_15_0_;
    wire sCounter_cry_8;
    wire sCounter_cry_9;
    wire sCounter_cry_10;
    wire sCounter_cry_11;
    wire sCounter_cry_12;
    wire sCounter_cry_13;
    wire sCounter_cry_14;
    wire sCounter_cry_15;
    wire bfn_8_16_0_;
    wire sCounter_cry_16;
    wire sCounter_cry_17;
    wire sCounter_cry_18;
    wire sCounter_cry_19;
    wire sCounter_cry_20;
    wire sCounter_cry_21;
    wire LED_ACQ_c_i;
    wire sCounter_cry_22;
    wire bfn_8_17_0_;
    wire un1_button_debounce_counter_cry_1;
    wire un1_button_debounce_counter_cry_2;
    wire un1_button_debounce_counter_cry_3;
    wire un1_button_debounce_counter_cry_4;
    wire button_debounce_counterZ0Z_6;
    wire un1_button_debounce_counter_cry_5;
    wire button_debounce_counterZ0Z_7;
    wire un1_button_debounce_counter_cry_6;
    wire button_debounce_counterZ0Z_8;
    wire un1_button_debounce_counter_cry_7;
    wire un1_button_debounce_counter_cry_8;
    wire button_debounce_counterZ0Z_9;
    wire bfn_8_18_0_;
    wire button_debounce_counterZ0Z_10;
    wire un1_button_debounce_counter_cry_9;
    wire button_debounce_counterZ0Z_11;
    wire un1_button_debounce_counter_cry_10;
    wire button_debounce_counterZ0Z_12;
    wire un1_button_debounce_counter_cry_11;
    wire button_debounce_counterZ0Z_13;
    wire un1_button_debounce_counter_cry_12;
    wire button_debounce_counterZ0Z_14;
    wire un1_button_debounce_counter_cry_13;
    wire button_debounce_counterZ0Z_15;
    wire un1_button_debounce_counter_cry_14;
    wire button_debounce_counterZ0Z_16;
    wire un1_button_debounce_counter_cry_15;
    wire un1_button_debounce_counter_cry_16;
    wire button_debounce_counterZ0Z_17;
    wire bfn_8_19_0_;
    wire button_debounce_counterZ0Z_18;
    wire un1_button_debounce_counter_cry_17;
    wire button_debounce_counterZ0Z_19;
    wire un1_button_debounce_counter_cry_18;
    wire button_debounce_counterZ0Z_20;
    wire un1_button_debounce_counter_cry_19;
    wire un1_button_debounce_counter_cry_20;
    wire un1_button_debounce_counter_cry_21;
    wire un1_button_debounce_counter_cry_22;
    wire un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO;
    wire un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO;
    wire bfn_8_20_0_;
    wire button_debounce_counterZ0Z_23;
    wire bfn_9_3_0_;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0 ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1 ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2 ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3 ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4 ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO ;
    wire \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11 ;
    wire \spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10 ;
    wire \spi_master_inst.sclk_gen_u0.N_158_7 ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ;
    wire \spi_master_inst.sclk_gen_u0.N_158_7_cascade_ ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ;
    wire \spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0 ;
    wire \spi_master_inst.sclk_gen_u0.falling_count_start_iZ0 ;
    wire un3_trig_0_0;
    wire un3_trig_0_0_cascade_;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2 ;
    wire \spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2 ;
    wire trig_ext_c;
    wire trig_rpi_c;
    wire trig_ft_c;
    wire un8_trig_prev_0_c5_a0_0_0_cascade_;
    wire un8_trig_prev_0_c4_a0_1_cascade_;
    wire sEETrigCounterZ0Z_5;
    wire sEETrigCounterZ0Z_6;
    wire sEETrigCounterZ0Z_7;
    wire un8_trig_prev_0_c7_a0_1_cascade_;
    wire un8_trig_prev_0_c4_a0_1;
    wire sEETrigCounterZ0Z_4;
    wire un8_trig_prev_0_c5_a0_0;
    wire sTrigCounter_i_0;
    wire bfn_9_8_0_;
    wire sTrigCounter_i_1;
    wire un10_trig_prev_cry_0;
    wire sTrigCounter_i_2;
    wire un10_trig_prev_cry_1;
    wire sTrigCounter_i_3;
    wire un10_trig_prev_cry_2;
    wire un10_trig_prev_4;
    wire sTrigCounter_i_4;
    wire un10_trig_prev_cry_3;
    wire un10_trig_prev_5;
    wire sTrigCounter_i_5;
    wire un10_trig_prev_cry_4;
    wire un10_trig_prev_6;
    wire sTrigCounter_i_6;
    wire un10_trig_prev_cry_5;
    wire un10_trig_prev_7;
    wire sTrigCounter_i_7;
    wire un10_trig_prev_cry_6;
    wire un10_trig_prev_cry_7;
    wire bfn_9_9_0_;
    wire sAddress_RNI9IH12_1Z0Z_1;
    wire trig_prevZ0;
    wire un3_trig_0_3;
    wire g1_0_0_2;
    wire g1_0_0;
    wire g1_0;
    wire sPeriod_prevZ0;
    wire LED_MODE_c;
    wire sTrigCounterZ0Z_4;
    wire sTrigCounterZ0Z_3;
    wire un1_sTrigCounter_ac0_0_0_cascade_;
    wire un1_reset_rpi_inv_2_i_o3_0_0;
    wire un1_sTrigCounter_ac0_0_2_0_cascade_;
    wire un10_trig_prev_cry_7_THRU_CO;
    wire sTrigCounterZ0Z_5;
    wire un1_sTrigCounter_ac0_0_2;
    wire un1_sTrigCounter_ac0_3_out_cascade_;
    wire sTrigCounterZ0Z_2;
    wire g1_0_1_0;
    wire g1_3_0;
    wire sEEPeriodZ0Z_10;
    wire sEEPeriodZ0Z_11;
    wire sEEPeriodZ0Z_12;
    wire sEEPeriodZ0Z_13;
    wire sEEPeriodZ0Z_14;
    wire sEEPeriodZ0Z_15;
    wire sEEPeriodZ0Z_8;
    wire sEEPeriodZ0Z_9;
    wire op_gt_op_gt_un13_striginternallto23_12;
    wire un1_reset_rpi_inv_2_i_o3_12;
    wire op_gt_op_gt_un13_striginternallto23_15;
    wire sEETrigInternal_prevZ0;
    wire N_5_0;
    wire un4_speriod_cry_23_THRU_CO;
    wire un1_reset_rpi_inv_2_i_1_1_0_cascade_;
    wire un1_reset_rpi_inv_2_i_1_cascade_;
    wire un1_sTrigCounter_ac0_0_4;
    wire sTrigCounterZ0Z_6;
    wire un1_sTrigCounter_axbxc7_m7_0_a2_2;
    wire un1_reset_rpi_inv_2_i_1;
    wire N_123;
    wire sTrigCounterZ0Z_7;
    wire bfn_9_13_0_;
    wire un1_spoff_cry_0;
    wire un1_spoff_cry_1;
    wire un1_spoff_cry_2;
    wire un1_spoff_cry_3;
    wire un1_spoff_cry_4;
    wire un1_spoff_cry_5;
    wire un1_spoff_cry_6;
    wire un1_spoff_cry_7;
    wire bfn_9_14_0_;
    wire un1_spoff_cry_8;
    wire un1_spoff_cry_9;
    wire un1_spoff_cry_10;
    wire un1_spoff_cry_11;
    wire un1_spoff_cry_12;
    wire un1_spoff_cry_13;
    wire un1_spoff_cry_14;
    wire un1_spoff_cry_15;
    wire sCounter_i_16;
    wire bfn_9_15_0_;
    wire sCounter_i_17;
    wire un1_spoff_cry_16;
    wire sCounter_i_18;
    wire un1_spoff_cry_17;
    wire sCounter_i_19;
    wire un1_spoff_cry_18;
    wire sCounter_i_20;
    wire un1_spoff_cry_19;
    wire sCounter_i_21;
    wire un1_spoff_cry_20;
    wire sCounter_i_22;
    wire un1_spoff_cry_21;
    wire sCounter_i_23;
    wire un1_spoff_cry_22;
    wire un1_spoff_cry_23;
    wire un4_spoff_cry_23_THRU_CO;
    wire bfn_9_16_0_;
    wire N_1612_i;
    wire sCounterRAMZ0Z_6;
    wire sCounterRAMZ0Z_3;
    wire button_debounce_counterZ0Z_21;
    wire button_debounce_counterZ0Z_22;
    wire sbuttonModeStatus_0_sqmuxa_0;
    wire sbuttonModeStatus_0_sqmuxa_18;
    wire button_debounce_counterZ0Z_4;
    wire button_debounce_counterZ0Z_3;
    wire button_debounce_counterZ0Z_5;
    wire button_debounce_counterZ0Z_2;
    wire sbuttonModeStatus_0_sqmuxa_13;
    wire sEEDelayACQ_i_0;
    wire bfn_9_17_0_;
    wire sEEDelayACQ_i_1;
    wire un4_sacqtime_cry_0;
    wire sEEDelayACQ_i_2;
    wire un4_sacqtime_cry_1;
    wire sEEDelayACQ_i_3;
    wire un4_sacqtime_cry_2;
    wire sEEDelayACQ_i_4;
    wire un4_sacqtime_cry_3;
    wire sEEDelayACQ_i_5;
    wire un4_sacqtime_cry_4;
    wire sEEDelayACQ_i_6;
    wire un4_sacqtime_cry_5;
    wire sEEDelayACQ_i_7;
    wire un4_sacqtime_cry_6;
    wire un4_sacqtime_cry_7;
    wire sEEDelayACQ_i_8;
    wire bfn_9_18_0_;
    wire sEEDelayACQ_i_9;
    wire un4_sacqtime_cry_8;
    wire sEEDelayACQ_i_10;
    wire un4_sacqtime_cry_9;
    wire sEEDelayACQ_i_11;
    wire un4_sacqtime_cry_10;
    wire sEEDelayACQ_i_12;
    wire un4_sacqtime_cry_11;
    wire sEEDelayACQ_i_13;
    wire un4_sacqtime_cry_12;
    wire sEEDelayACQ_i_14;
    wire un4_sacqtime_cry_13;
    wire sEEDelayACQ_i_15;
    wire un4_sacqtime_cry_14;
    wire un4_sacqtime_cry_15;
    wire bfn_9_19_0_;
    wire un4_sacqtime_cry_16;
    wire un4_sacqtime_cry_17;
    wire un4_sacqtime_cry_18;
    wire un4_sacqtime_cry_19;
    wire op_gt_op_gt_un13_striginternallto23_8;
    wire un4_sacqtime_cry_20;
    wire un4_sacqtime_cry_21;
    wire un4_sacqtime_cry_22;
    wire un4_sacqtime_cry_23;
    wire bfn_9_20_0_;
    wire LED3_c_0;
    wire bfn_10_2_0_;
    wire \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0 ;
    wire \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1 ;
    wire \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2 ;
    wire \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3 ;
    wire \spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4 ;
    wire \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_i6_3_cascade_ ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2 ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_ ;
    wire \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_5 ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3 ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1 ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0 ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4 ;
    wire \spi_slave_inst.un23_i_ssn_3_cascade_ ;
    wire \spi_slave_inst.un23_i_ssn ;
    wire \spi_slave_inst.un23_i_ssn_cascade_ ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa ;
    wire \spi_slave_inst.un23_i_ssn_3 ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5 ;
    wire \spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_6 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_1 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_2 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_11 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_12 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_3 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_14 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_15 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0 ;
    wire bfn_10_6_0_;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5 ;
    wire \spi_master_inst.sclk_gen_u0.falling_count_start_i_i ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7 ;
    wire \spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i ;
    wire sEETrigCounterZ0Z_3;
    wire un10_trig_prev_3;
    wire sEETrigCounterZ0Z_2;
    wire un10_trig_prev_2;
    wire un10_trig_prev_0;
    wire sEETrigCounterZ0Z_0;
    wire sEETrigCounterZ0Z_1;
    wire un10_trig_prev_1;
    wire \spi_slave_inst.rx_done_reg3_iZ0 ;
    wire \spi_slave_inst.rx_ready_i_RNOZ0Z_0_cascade_ ;
    wire \spi_slave_inst.un4_tx_done_reg2_i_cascade_ ;
    wire button_debounce_counterZ0Z_0;
    wire button_debounce_counterZ0Z_1;
    wire N_3089_g;
    wire spi_mosi_ready_prevZ0Z2;
    wire spi_mosi_ready_prevZ0;
    wire spi_mosi_ready_prevZ0Z3;
    wire spi_mosi_ready_prev3_RNILKERZ0_cascade_;
    wire \spi_slave_inst.tx_ready_iZ0 ;
    wire sCounter_i_0;
    wire bfn_10_14_0_;
    wire sCounter_i_1;
    wire un1_sacqtime_cry_0;
    wire sCounter_i_2;
    wire un1_sacqtime_cry_1;
    wire sCounter_i_3;
    wire un1_sacqtime_cry_2;
    wire sCounter_i_4;
    wire un1_sacqtime_cry_3;
    wire sCounter_i_5;
    wire un1_sacqtime_cry_4;
    wire sCounter_i_6;
    wire un1_sacqtime_cry_5;
    wire sCounter_i_7;
    wire un1_sacqtime_cry_6;
    wire un1_sacqtime_cry_7;
    wire sCounter_i_8;
    wire bfn_10_15_0_;
    wire sCounter_i_9;
    wire un1_sacqtime_cry_8;
    wire sCounter_i_10;
    wire un1_sacqtime_cry_9;
    wire sCounter_i_11;
    wire un1_sacqtime_cry_10;
    wire sCounter_i_12;
    wire un1_sacqtime_cry_11;
    wire sCounter_i_13;
    wire un1_sacqtime_cry_12;
    wire sCounter_i_14;
    wire un1_sacqtime_cry_13;
    wire sCounter_i_15;
    wire un1_sacqtime_cry_14;
    wire un1_sacqtime_cry_15;
    wire un1_sacqtime_cry_16_sf;
    wire bfn_10_16_0_;
    wire un1_sacqtime_cry_17_sf;
    wire un1_sacqtime_cry_16;
    wire un1_sacqtime_cry_18_sf;
    wire un1_sacqtime_cry_17;
    wire un1_sacqtime_cry_19_sf;
    wire un1_sacqtime_cry_18;
    wire un1_sacqtime_cry_20_sf;
    wire un1_sacqtime_cry_19;
    wire un1_sacqtime_cry_21_sf;
    wire un1_sacqtime_cry_20;
    wire un1_sacqtime_cry_22_sf;
    wire un1_sacqtime_cry_21;
    wire un1_sacqtime_cry_23_sf;
    wire un1_sacqtime_cry_22;
    wire un1_sacqtime_cry_23;
    wire bfn_10_17_0_;
    wire RAM_DATA_cl_10Z0Z_15;
    wire N_106;
    wire N_26;
    wire N_76_i;
    wire N_71_cascade_;
    wire sEEDelayACQZ0Z_0;
    wire sEEDelayACQZ0Z_1;
    wire sEEDelayACQZ0Z_2;
    wire sEEDelayACQZ0Z_3;
    wire sEEDelayACQZ0Z_4;
    wire sEEDelayACQZ0Z_5;
    wire sEEDelayACQZ0Z_6;
    wire sEEDelayACQZ0Z_7;
    wire sEEDelayACQZ0Z_10;
    wire sEEDelayACQZ0Z_11;
    wire sEEDelayACQZ0Z_12;
    wire sEEDelayACQZ0Z_13;
    wire sEEDelayACQZ0Z_14;
    wire sEEDelayACQZ0Z_15;
    wire sEEDelayACQZ0Z_8;
    wire sEEDelayACQZ0Z_9;
    wire sAddress_RNIA6242Z0Z_0;
    wire N_99_cascade_;
    wire RAM_DATA_cl_12Z0Z_15;
    wire N_94_cascade_;
    wire RAM_DATA_cl_11Z0Z_15;
    wire N_104_cascade_;
    wire RAM_DATA_cl_14Z0Z_15;
    wire sDAC_dataZ0Z_2;
    wire \spi_slave_inst.rx_data_count_neg_sclk_i6 ;
    wire \INVspi_slave_inst.rx_done_neg_sclk_iC_net ;
    wire \spi_slave_inst.rx_done_neg_sclk_iZ0 ;
    wire \spi_slave_inst.rx_done_pos_sclk_iZ0 ;
    wire \spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0 ;
    wire \spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0 ;
    wire \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0 ;
    wire \spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0 ;
    wire \spi_master_inst.sclk_gen_u0.spi_start_iZ0 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_4 ;
    wire \spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3_cascade_ ;
    wire \spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0 ;
    wire \spi_slave_inst.N_1394 ;
    wire \spi_slave_inst.N_1397_cascade_ ;
    wire \spi_slave_inst.tx_done_reg1_iZ0 ;
    wire \spi_slave_inst.tx_done_reg2_iZ0 ;
    wire \spi_slave_inst.tx_done_reg3_iZ0 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_0 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_3 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_7 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_5 ;
    wire \spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_1 ;
    wire \spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_2 ;
    wire \spi_slave_inst.txdata_reg_iZ0Z_6 ;
    wire N_206;
    wire N_206_cascade_;
    wire sAddress_RNIA6242_1Z0Z_0;
    wire spi_mosi_ready64_prevZ0Z2;
    wire spi_mosi_ready64_prevZ0;
    wire spi_mosi_ready64_prevZ0Z3;
    wire spi_mosi_ready;
    wire spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_;
    wire LED3_c_i;
    wire \spi_slave_inst.data_in_reg_iZ0Z_0 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_1 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_2 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_3 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_4 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_5 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_6 ;
    wire \spi_slave_inst.data_in_reg_iZ0Z_7 ;
    wire \spi_slave_inst.un4_i_wr ;
    wire RAM_DATA_in_6;
    wire RAM_DATA_in_14;
    wire spi_data_misoZ0Z_6;
    wire RAM_DATA_in_7;
    wire RAM_DATA_in_15;
    wire spi_data_misoZ0Z_7;
    wire RAM_nWE_0_i;
    wire sADC_clk_prevZ0;
    wire ADC_clk_c;
    wire N_127;
    wire N_1470_i;
    wire N_86;
    wire sRead_dataZ0;
    wire sCounterRAMZ0Z_5;
    wire sCounterRAMZ0Z_4;
    wire sCounterRAMZ0Z_7;
    wire sCounterRAMZ0Z_0;
    wire sCounterRAMZ0Z_2;
    wire sCounterRAMZ0Z_1;
    wire spi_data_miso_0_sqmuxa_2_i_o2_5_cascade_;
    wire spi_data_miso_0_sqmuxa_2_i_o2_4;
    wire N_75_cascade_;
    wire sSPI_MSB0LSBZ0Z1;
    wire spi_mosi_ready_prev3_RNILKERZ0;
    wire N_88;
    wire N_88_cascade_;
    wire N_28;
    wire N_93_cascade_;
    wire RAM_DATA_cl_9Z0Z_15;
    wire N_98_cascade_;
    wire RAM_DATA_clZ0Z_15;
    wire N_96_cascade_;
    wire RAM_DATA_cl_8Z0Z_15;
    wire sRAM_pointer_readZ0Z_14;
    wire RAM_ADD_c_14;
    wire sRAM_pointer_readZ0Z_15;
    wire RAM_ADD_c_15;
    wire sRAM_pointer_readZ0Z_16;
    wire RAM_ADD_c_16;
    wire sRAM_pointer_readZ0Z_17;
    wire RAM_ADD_c_17;
    wire sRAM_pointer_readZ0Z_18;
    wire RAM_ADD_c_18;
    wire sRAM_pointer_readZ0Z_2;
    wire RAM_ADD_c_2;
    wire sRAM_pointer_readZ0Z_3;
    wire RAM_ADD_c_3;
    wire sRAM_pointer_readZ0Z_4;
    wire RAM_ADD_c_4;
    wire sRAM_pointer_readZ0Z_5;
    wire RAM_ADD_c_5;
    wire sRAM_pointer_readZ0Z_6;
    wire RAM_ADD_c_6;
    wire sRAM_pointer_readZ0Z_7;
    wire RAM_ADD_c_7;
    wire sRAM_pointer_readZ0Z_8;
    wire RAM_ADD_c_8;
    wire sRAM_pointer_readZ0Z_9;
    wire RAM_ADD_c_9;
    wire N_102;
    wire RAM_DATA_cl_15Z0Z_15;
    wire spi_sclk_ft_c;
    wire spi_sclk;
    wire \spi_slave_inst.rx_done_reg1_iZ0 ;
    wire \spi_slave_inst.rx_done_reg2_iZ0 ;
    wire \spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_10 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_13 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_4 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_5 ;
    wire sDAC_dataZ0Z_0;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_0 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_7 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_8 ;
    wire \spi_master_inst.spi_data_path_u1.data_inZ0Z_9 ;
    wire \spi_master_inst.spi_data_path_u1.tx_ready_iZ0 ;
    wire un1_spointer11_5_0_2_cascade_;
    wire sAddress_RNIA6242_0Z0Z_2;
    wire sDAC_mem_23_1_sqmuxa;
    wire N_275_cascade_;
    wire N_360_cascade_;
    wire N_269;
    wire N_132;
    wire sAddress_RNIA6242_0Z0Z_0;
    wire un1_spointer11_7_0_tz;
    wire un1_spointer11_7_0_tz_cascade_;
    wire sAddress_RNID9242Z0Z_3;
    wire \spi_slave_inst.un1_spointer11_2_0_a2_0_6_4 ;
    wire \spi_slave_inst.un1_spointer11_2_0_a2_0_6_5_cascade_ ;
    wire un1_spointer11_2_0;
    wire N_285_cascade_;
    wire sPointerZ0Z_0;
    wire N_116_cascade_;
    wire N_159;
    wire N_117_cascade_;
    wire spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1;
    wire sEETrigInternalZ0;
    wire sEEPoffZ0Z_0;
    wire sEEPoffZ0Z_1;
    wire sEEPoffZ0Z_2;
    wire sEEPoffZ0Z_3;
    wire sEEPoffZ0Z_4;
    wire sEEPoffZ0Z_5;
    wire sEEPoffZ0Z_6;
    wire sEEPoffZ0Z_7;
    wire sEEPoffZ0Z_10;
    wire sEEPoffZ0Z_11;
    wire sEEPoffZ0Z_12;
    wire sEEPoffZ0Z_13;
    wire sEEPoffZ0Z_14;
    wire sEEPoffZ0Z_15;
    wire sEEPoffZ0Z_8;
    wire sEEPoffZ0Z_9;
    wire sAddress_RNIA6242_1Z0Z_2;
    wire bfn_12_15_0_;
    wire sCounterADC_cry_0;
    wire sCounterADC_cry_1;
    wire sCounterADC_cry_2;
    wire sCounterADC_cry_3;
    wire sCounterADC_cry_4;
    wire sCounterADC_cry_5;
    wire sCounterADC_cry_6;
    wire RAM_DATA_in_8;
    wire RAM_DATA_in_0;
    wire spi_data_misoZ0Z_0;
    wire RAM_DATA_in_9;
    wire RAM_DATA_in_1;
    wire spi_data_misoZ0Z_1;
    wire RAM_DATA_in_10;
    wire RAM_DATA_in_2;
    wire spi_data_misoZ0Z_2;
    wire RAM_DATA_in_11;
    wire RAM_DATA_in_3;
    wire spi_data_misoZ0Z_3;
    wire RAM_DATA_in_12;
    wire RAM_DATA_in_4;
    wire spi_data_misoZ0Z_4;
    wire un4_sacqtime_cry_23_c_RNITTSZ0Z3;
    wire RAM_DATA_in_5;
    wire N_75;
    wire RAM_DATA_in_13;
    wire spi_data_misoZ0Z_5;
    wire N_6;
    wire sRAM_pointer_readZ0Z_0;
    wire RAM_ADD_c_0;
    wire reset_rpi_ibuf_RNI7JCVZ0;
    wire sRAM_ADD_0_sqmuxa_i_0;
    wire sRAM_pointer_readZ0Z_1;
    wire RAM_ADD_c_1;
    wire sRAM_pointer_readZ0Z_10;
    wire RAM_ADD_c_10;
    wire sRAM_pointer_readZ0Z_11;
    wire RAM_ADD_c_11;
    wire sRAM_pointer_readZ0Z_12;
    wire RAM_ADD_c_12;
    wire sRAM_pointer_readZ0Z_13;
    wire RAM_ADD_c_13;
    wire N_67_i;
    wire ADC3_c;
    wire RAM_DATA_1Z0Z_3;
    wire ADC0_c;
    wire RAM_DATA_1Z0Z_0;
    wire ADC5_c;
    wire RAM_DATA_1Z0Z_5;
    wire ADC1_c;
    wire RAM_DATA_1Z0Z_1;
    wire ADC7_c;
    wire RAM_DATA_1Z0Z_8;
    wire ADC8_c;
    wire RAM_DATA_1Z0Z_9;
    wire RAM_DATA_1Z0Z_15;
    wire RAM_DATA_1Z0Z_7;
    wire RAM_DATA_cl_1Z0Z_15;
    wire N_100;
    wire RAM_DATA_cl_13Z0Z_15;
    wire N_97;
    wire RAM_DATA_cl_2Z0Z_15;
    wire N_101;
    wire N_103;
    wire RAM_DATA_cl_3Z0Z_15;
    wire spi_mosi_ft_c;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6 ;
    wire \spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7 ;
    wire spi_sclk_g;
    wire \spi_slave_inst.spi_cs_iZ0 ;
    wire sDAC_mem_23Z0Z_2;
    wire sDAC_mem_22Z0Z_2;
    wire sDAC_mem_23Z0Z_3;
    wire sDAC_mem_22Z0Z_3;
    wire sDAC_mem_23Z0Z_4;
    wire sDAC_mem_22Z0Z_4;
    wire N_291_cascade_;
    wire sEEPonPoff_1_sqmuxa;
    wire sAddressZ0Z_6;
    wire sAddressZ0Z_7;
    wire sEEPonPoff_1_sqmuxa_0_a2_1;
    wire sEEPon_1_sqmuxa;
    wire N_291;
    wire sDAC_mem_33_1_sqmuxa;
    wire sDAC_mem_17_1_sqmuxa;
    wire sDAC_mem_32_1_sqmuxa;
    wire N_141;
    wire sEETrigCounter_1_sqmuxa;
    wire N_1480_cascade_;
    wire un1_spointer11_5_0_2;
    wire sAddress_RNIA6242_2Z0Z_2;
    wire N_280_cascade_;
    wire sDAC_mem_19_1_sqmuxa;
    wire sDAC_mem_19Z0Z_4;
    wire sDAC_mem_18Z0Z_4;
    wire sDAC_mem_19Z0Z_5;
    wire sDAC_mem_18Z0Z_5;
    wire sDAC_mem_19Z0Z_6;
    wire sDAC_mem_18Z0Z_6;
    wire sAddress_RNIA6242Z0Z_2;
    wire ADC4_c;
    wire RAM_DATA_1Z0Z_4;
    wire ADC6_c;
    wire RAM_DATA_1Z0Z_6;
    wire ADC9_c;
    wire RAM_DATA_1Z0Z_10;
    wire top_tour1_c;
    wire RAM_DATA_1Z0Z_11;
    wire top_tour2_c;
    wire RAM_DATA_1Z0Z_12;
    wire sTrigCounterZ0Z_0;
    wire RAM_DATA_1Z0Z_13;
    wire sTrigCounterZ0Z_1;
    wire RAM_DATA_1Z0Z_14;
    wire ADC2_c;
    wire RAM_DATA_1Z0Z_2;
    wire N_31_i;
    wire N_107_cascade_;
    wire RAM_DATA_cl_5Z0Z_15;
    wire N_108_cascade_;
    wire RAM_DATA_cl_6Z0Z_15;
    wire LED3_c;
    wire un4_sacqtime_cry_23_THRU_CO;
    wire N_95_cascade_;
    wire un1_sacqtime_cry_23_THRU_CO;
    wire RAM_DATA_cl_7Z0Z_15;
    wire RAM_DATA_cl_4Z0Z_15;
    wire N_71;
    wire N_105;
    wire sRAM_pointer_writeZ0Z_0;
    wire bfn_13_18_0_;
    wire sRAM_pointer_writeZ0Z_1;
    wire sRAM_pointer_write_cry_0;
    wire sRAM_pointer_writeZ0Z_2;
    wire sRAM_pointer_write_cry_1;
    wire sRAM_pointer_writeZ0Z_3;
    wire sRAM_pointer_write_cry_2;
    wire sRAM_pointer_writeZ0Z_4;
    wire sRAM_pointer_write_cry_3;
    wire sRAM_pointer_writeZ0Z_5;
    wire sRAM_pointer_write_cry_4;
    wire sRAM_pointer_writeZ0Z_6;
    wire sRAM_pointer_write_cry_5;
    wire sRAM_pointer_writeZ0Z_7;
    wire sRAM_pointer_write_cry_6;
    wire sRAM_pointer_write_cry_7;
    wire sRAM_pointer_writeZ0Z_8;
    wire bfn_13_19_0_;
    wire sRAM_pointer_writeZ0Z_9;
    wire sRAM_pointer_write_cry_8;
    wire sRAM_pointer_writeZ0Z_10;
    wire sRAM_pointer_write_cry_9;
    wire sRAM_pointer_writeZ0Z_11;
    wire sRAM_pointer_write_cry_10;
    wire sRAM_pointer_writeZ0Z_12;
    wire sRAM_pointer_write_cry_11;
    wire sRAM_pointer_writeZ0Z_13;
    wire sRAM_pointer_write_cry_12;
    wire sRAM_pointer_writeZ0Z_14;
    wire sRAM_pointer_write_cry_13;
    wire sRAM_pointer_writeZ0Z_15;
    wire sRAM_pointer_write_cry_14;
    wire sRAM_pointer_write_cry_15;
    wire sRAM_pointer_writeZ0Z_16;
    wire bfn_13_20_0_;
    wire sRAM_pointer_writeZ0Z_17;
    wire sRAM_pointer_write_cry_16;
    wire sEEPointerResetZ0;
    wire sRAM_pointer_write_cry_17;
    wire sRAM_pointer_writeZ0Z_18;
    wire N_26_g;
    wire spi_cs_ft_c;
    wire \spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_ ;
    wire \spi_slave_inst.spi_csZ0 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_ ;
    wire \spi_slave_inst.tx_done_neg_sclk_iZ0 ;
    wire \INVspi_slave_inst.tx_done_neg_sclk_iC_net ;
    wire spi_miso_flash_c;
    wire spi_miso_rpi_c;
    wire sDAC_data_2_13_bm_1_3_cascade_;
    wire sDAC_mem_6Z0Z_0;
    wire sDAC_mem_38Z0Z_1;
    wire sDAC_data_2_13_bm_1_4_cascade_;
    wire sDAC_mem_6Z0Z_1;
    wire sDAC_mem_6Z0Z_2;
    wire sDAC_data_2_13_bm_1_5_cascade_;
    wire sDAC_data_2_13_am_1_5_cascade_;
    wire sDAC_mem_4Z0Z_2;
    wire sDAC_data_2_13_am_1_6_cascade_;
    wire sDAC_mem_4Z0Z_3;
    wire sDAC_mem_4Z0Z_4;
    wire sDAC_data_2_13_am_1_7_cascade_;
    wire sDAC_mem_2Z0Z_0;
    wire sDAC_data_2_6_bm_1_3_cascade_;
    wire sDAC_mem_3Z0Z_0;
    wire sDAC_data_RNO_17Z0Z_5_cascade_;
    wire sDAC_data_2_20_am_1_5_cascade_;
    wire sDAC_data_RNO_7Z0Z_5_cascade_;
    wire sDAC_data_RNO_8Z0Z_5;
    wire sDAC_data_RNO_21Z0Z_5;
    wire sDAC_data_RNO_10Z0Z_5_cascade_;
    wire sDAC_data_2_32_ns_1_5;
    wire sDAC_data_RNO_5Z0Z_5;
    wire sDAC_data_2_14_ns_1_5_cascade_;
    wire sDAC_data_RNO_4Z0Z_5;
    wire sDAC_data_RNO_2Z0Z_5;
    wire sDAC_data_RNO_1Z0Z_5_cascade_;
    wire sDAC_data_2_41_ns_1_5;
    wire sDAC_data_2_5_cascade_;
    wire sDAC_dataZ0Z_5;
    wire sDAC_mem_2Z0Z_2;
    wire sDAC_data_2_6_bm_1_5_cascade_;
    wire sDAC_mem_3Z0Z_2;
    wire sDAC_data_RNO_15Z0Z_5;
    wire sDAC_data_2_20_am_1_7_cascade_;
    wire sDAC_data_RNO_17Z0Z_7_cascade_;
    wire sDAC_data_RNO_8Z0Z_7_cascade_;
    wire sDAC_data_RNO_7Z0Z_7;
    wire sDAC_mem_33Z0Z_5;
    wire sDAC_data_RNO_27Z0Z_8_cascade_;
    wire sDAC_mem_32Z0Z_5;
    wire sDAC_data_RNO_26Z0Z_8;
    wire sDAC_mem_1Z0Z_5;
    wire sDAC_mem_33Z0Z_6;
    wire sDAC_data_RNO_26Z0Z_9_cascade_;
    wire sDAC_mem_32Z0Z_6;
    wire sDAC_data_RNO_27Z0Z_9;
    wire sDAC_mem_1Z0Z_6;
    wire sDAC_mem_2Z0Z_6;
    wire sDAC_data_2_6_bm_1_9_cascade_;
    wire sDAC_mem_3Z0Z_6;
    wire sDAC_mem_33Z0Z_1;
    wire sDAC_data_RNO_26Z0Z_4_cascade_;
    wire sDAC_mem_1Z0Z_1;
    wire sDAC_mem_32Z0Z_1;
    wire sDAC_data_RNO_27Z0Z_4;
    wire sDAC_mem_33Z0Z_2;
    wire sDAC_data_RNO_26Z0Z_5_cascade_;
    wire sDAC_data_RNO_14Z0Z_5;
    wire sDAC_mem_32Z0Z_2;
    wire sDAC_mem_1Z0Z_2;
    wire sDAC_data_RNO_27Z0Z_5;
    wire op_le_op_le_un15_sdacdynlt4_cascade_;
    wire un17_sdacdyn_0;
    wire sDAC_mem_10Z0Z_7;
    wire sDAC_mem_19Z0Z_7;
    wire sDAC_mem_18Z0Z_7;
    wire sDAC_mem_19Z0Z_0;
    wire sDAC_mem_18Z0Z_0;
    wire sDAC_mem_19Z0Z_1;
    wire sDAC_mem_18Z0Z_1;
    wire sDAC_mem_19Z0Z_2;
    wire sDAC_data_RNO_30Z0Z_5;
    wire sDAC_mem_18Z0Z_2;
    wire sDAC_mem_18_1_sqmuxa;
    wire sDAC_data_RNO_18Z0Z_5_cascade_;
    wire sDAC_data_RNO_19Z0Z_5;
    wire sDAC_data_2_24_ns_1_5;
    wire sDAC_data_RNO_18Z0Z_6_cascade_;
    wire sDAC_data_RNO_19Z0Z_6;
    wire sDAC_mem_12Z0Z_2;
    wire sDAC_mem_12Z0Z_3;
    wire sDAC_mem_31_1_sqmuxa;
    wire sCounterADCZ0Z_3;
    wire sCounterADCZ0Z_2;
    wire sEEADC_freqZ0Z_2;
    wire sEEADC_freqZ0Z_3;
    wire sCounterADCZ0Z_5;
    wire sCounterADCZ0Z_4;
    wire sEEADC_freqZ0Z_4;
    wire sEEADC_freqZ0Z_5;
    wire sCounterADCZ0Z_6;
    wire sCounterADCZ0Z_7;
    wire un7_spon_0;
    wire sEEACQZ0Z_0;
    wire sEEACQ_i_0;
    wire bfn_14_16_0_;
    wire sEEACQZ0Z_1;
    wire un7_spon_1;
    wire sEEACQ_i_1;
    wire un5_sdacdyn_cry_0;
    wire un7_spon_2;
    wire sEEACQZ0Z_2;
    wire sEEACQ_i_2;
    wire un5_sdacdyn_cry_1;
    wire un7_spon_3;
    wire sEEACQZ0Z_3;
    wire sEEACQ_i_3;
    wire un5_sdacdyn_cry_2;
    wire sEEACQZ0Z_4;
    wire sEEACQ_i_4;
    wire un5_sdacdyn_cry_3;
    wire un7_spon_5;
    wire sEEACQZ0Z_5;
    wire sEEACQ_i_5;
    wire un5_sdacdyn_cry_4;
    wire un7_spon_6;
    wire sEEACQZ0Z_6;
    wire sEEACQ_i_6;
    wire un5_sdacdyn_cry_5;
    wire un7_spon_7;
    wire sEEACQZ0Z_7;
    wire sEEACQ_i_7;
    wire un5_sdacdyn_cry_6;
    wire un5_sdacdyn_cry_7;
    wire un7_spon_8;
    wire sEEACQZ0Z_8;
    wire sEEACQ_i_8;
    wire bfn_14_17_0_;
    wire un7_spon_9;
    wire sEEACQZ0Z_9;
    wire sEEACQ_i_9;
    wire un5_sdacdyn_cry_8;
    wire un7_spon_10;
    wire sEEACQZ0Z_10;
    wire sEEACQ_i_10;
    wire un5_sdacdyn_cry_9;
    wire un7_spon_11;
    wire sEEACQZ0Z_11;
    wire sEEACQ_i_11;
    wire un5_sdacdyn_cry_10;
    wire sEEACQZ0Z_12;
    wire un7_spon_12;
    wire sEEACQ_i_12;
    wire un5_sdacdyn_cry_11;
    wire un7_spon_13;
    wire sEEACQZ0Z_13;
    wire sEEACQ_i_13;
    wire un5_sdacdyn_cry_12;
    wire un7_spon_14;
    wire sEEACQZ0Z_14;
    wire sEEACQ_i_14;
    wire un5_sdacdyn_cry_13;
    wire un7_spon_15;
    wire sEEACQZ0Z_15;
    wire sEEACQ_i_15;
    wire un5_sdacdyn_cry_14;
    wire un5_sdacdyn_cry_15;
    wire un7_spon_16;
    wire bfn_14_18_0_;
    wire un7_spon_17;
    wire un5_sdacdyn_cry_16;
    wire un7_spon_18;
    wire un5_sdacdyn_cry_17;
    wire un7_spon_19;
    wire un5_sdacdyn_cry_18;
    wire un7_spon_20;
    wire un5_sdacdyn_cry_19;
    wire un7_spon_21;
    wire un5_sdacdyn_cry_20;
    wire un7_spon_22;
    wire un5_sdacdyn_cry_21;
    wire un7_spon_23;
    wire un5_sdacdyn_cry_22;
    wire un5_sdacdyn_cry_23;
    wire un17_sdacdyn_1;
    wire N_1479;
    wire un7_spon_4;
    wire bfn_14_19_0_;
    wire sDAC_mem_24Z0Z_3;
    wire sDAC_mem_24Z0Z_6;
    wire sDAC_mem_17Z0Z_2;
    wire sDAC_data_RNO_29Z0Z_5;
    wire sDAC_mem_16Z0Z_2;
    wire sDAC_mem_pointerZ0Z_6;
    wire sDAC_mem_pointerZ0Z_7;
    wire \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0 ;
    wire bfn_15_2_0_;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1 ;
    wire \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_i6 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2 ;
    wire \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3 ;
    wire \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4 ;
    wire \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3 ;
    wire \spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4 ;
    wire \spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5 ;
    wire \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ;
    wire sDAC_mem_34Z0Z_0;
    wire sDAC_mem_34Z0Z_2;
    wire sDAC_mem_34Z0Z_6;
    wire sDAC_mem_7Z0Z_0;
    wire sDAC_mem_7Z0Z_1;
    wire sDAC_mem_7Z0Z_2;
    wire sDAC_mem_5Z0Z_2;
    wire sDAC_mem_5Z0Z_3;
    wire sDAC_mem_5Z0Z_4;
    wire sDAC_mem_2_1_sqmuxa;
    wire sDAC_mem_5_1_sqmuxa;
    wire sDAC_mem_7_1_sqmuxa;
    wire N_279;
    wire N_279_cascade_;
    wire sDAC_data_RNO_21Z0Z_7;
    wire sDAC_data_2_14_ns_1_7_cascade_;
    wire sDAC_data_RNO_4Z0Z_7;
    wire sDAC_data_RNO_10Z0Z_7;
    wire sDAC_data_RNO_2Z0Z_7;
    wire sDAC_data_2_41_ns_1_7_cascade_;
    wire sDAC_data_RNO_1Z0Z_7;
    wire sDAC_data_2_7_cascade_;
    wire sDAC_dataZ0Z_7;
    wire sDAC_data_RNO_17Z0Z_9_cascade_;
    wire sDAC_data_RNO_8Z0Z_9_cascade_;
    wire sDAC_data_2_20_am_1_9_cascade_;
    wire sDAC_data_RNO_7Z0Z_9;
    wire sDAC_mem_17Z0Z_4;
    wire sDAC_mem_16Z0Z_4;
    wire sDAC_mem_17Z0Z_5;
    wire sDAC_mem_16Z0Z_5;
    wire sDAC_mem_17Z0Z_6;
    wire sDAC_mem_16Z0Z_6;
    wire bfn_15_10_0_;
    wire sDAC_mem_pointer_0_cry_1;
    wire sDAC_mem_pointer_0_cry_2;
    wire sDAC_mem_pointer_0_cry_3;
    wire sDAC_mem_pointer_0_cry_4;
    wire sDAC_data_RNO_23Z0Z_9_cascade_;
    wire sDAC_data_RNO_17Z0Z_10;
    wire sDAC_data_2_24_ns_1_10;
    wire sDAC_data_RNO_8Z0Z_10_cascade_;
    wire sDAC_data_2_20_am_1_10_cascade_;
    wire sDAC_data_RNO_7Z0Z_10;
    wire sDAC_mem_28Z0Z_6;
    wire sDAC_dataZ0Z_1;
    wire sDAC_dataZ0Z_11;
    wire sDAC_dataZ0Z_12;
    wire CONSTANT_ONE_NET;
    wire sDAC_dataZ0Z_13;
    wire sDAC_dataZ0Z_14;
    wire GNDG0;
    wire sDAC_dataZ0Z_15;
    wire sDAC_data_RNO_31Z0Z_8_cascade_;
    wire sDAC_data_2_39_ns_1_8_cascade_;
    wire sDAC_data_RNO_32Z0Z_8;
    wire sDAC_data_RNO_23Z0Z_8;
    wire sDAC_mem_31Z0Z_5;
    wire sDAC_data_RNO_24Z0Z_8;
    wire sDAC_mem_24Z0Z_5;
    wire sDAC_data_RNO_31Z0Z_9;
    wire sDAC_data_RNO_32Z0Z_9;
    wire sDAC_data_2_39_ns_1_9;
    wire sDAC_mem_26Z0Z_0;
    wire sDAC_mem_26Z0Z_5;
    wire sDAC_mem_26Z0Z_6;
    wire sDAC_data_RNO_18Z0Z_9_cascade_;
    wire sDAC_data_RNO_19Z0Z_9;
    wire sDAC_data_2_24_ns_1_9;
    wire sCounterADCZ0Z_1;
    wire sCounterADCZ0Z_0;
    wire un11_sacqtime_NE_3;
    wire un11_sacqtime_NE_2;
    wire un11_sacqtime_NE_0_0_cascade_;
    wire un11_sacqtime_NE_1;
    wire un11_sacqtime_NE_0;
    wire sDAC_mem_31Z0Z_6;
    wire sDAC_data_RNO_24Z0Z_9;
    wire sDAC_mem_29Z0Z_5;
    wire sDAC_mem_29Z0Z_6;
    wire sDAC_mem_29_1_sqmuxa;
    wire sDAC_mem_29Z0Z_3;
    wire sDAC_data_RNO_23Z0Z_6;
    wire sDAC_mem_24Z0Z_4;
    wire sDAC_data_RNO_31Z0Z_7_cascade_;
    wire sDAC_data_2_39_ns_1_7_cascade_;
    wire sDAC_data_RNO_11Z0Z_7;
    wire sDAC_mem_28Z0Z_3;
    wire sDAC_mem_26Z0Z_4;
    wire sDAC_data_RNO_32Z0Z_7;
    wire sDAC_mem_31Z0Z_3;
    wire sDAC_data_RNO_24Z0Z_6;
    wire sDAC_data_RNO_31Z0Z_5_cascade_;
    wire sDAC_data_2_39_ns_1_5_cascade_;
    wire sDAC_data_RNO_11Z0Z_5;
    wire sDAC_mem_26Z0Z_2;
    wire sDAC_data_RNO_32Z0Z_5;
    wire sDAC_mem_29Z0Z_2;
    wire sDAC_data_RNO_23Z0Z_5;
    wire sDAC_mem_31Z0Z_2;
    wire sDAC_data_RNO_24Z0Z_5;
    wire sDAC_mem_24Z0Z_2;
    wire sDAC_data_RNO_31Z0Z_6;
    wire sDAC_data_2_39_ns_1_6;
    wire sDAC_mem_29Z0Z_4;
    wire sDAC_data_RNO_23Z0Z_7;
    wire sDAC_mem_26Z0Z_3;
    wire sDAC_data_RNO_32Z0Z_6;
    wire sDAC_mem_24Z0Z_0;
    wire sDAC_mem_17Z0Z_3;
    wire \spi_slave_inst.spi_miso ;
    wire spi_select_c;
    wire spi_miso_ft_c;
    wire sDAC_mem_36Z0Z_2;
    wire sDAC_mem_36Z0Z_3;
    wire sDAC_mem_36Z0Z_4;
    wire sDAC_mem_37Z0Z_2;
    wire sDAC_mem_37Z0Z_3;
    wire sDAC_mem_37Z0Z_4;
    wire sDAC_mem_8Z0Z_2;
    wire sDAC_mem_8Z0Z_4;
    wire sDAC_mem_8Z0Z_6;
    wire sDAC_mem_8Z0Z_7;
    wire sDAC_mem_8_1_sqmuxa;
    wire sDAC_data_RNO_20Z0Z_7;
    wire sDAC_mem_20Z0Z_4;
    wire sDAC_mem_20Z0Z_5;
    wire sDAC_mem_20Z0Z_6;
    wire sDAC_mem_23Z0Z_7;
    wire sDAC_mem_22Z0Z_7;
    wire sDAC_mem_23Z0Z_0;
    wire sDAC_mem_22Z0Z_0;
    wire sDAC_data_2_13_bm_1_7_cascade_;
    wire sDAC_mem_7Z0Z_4;
    wire sDAC_data_RNO_5Z0Z_7;
    wire sDAC_data_RNO_30Z0Z_7;
    wire sDAC_data_RNO_29Z0Z_7;
    wire sDAC_data_2_32_ns_1_7;
    wire sDAC_mem_34Z0Z_4;
    wire sDAC_mem_2Z0Z_4;
    wire sDAC_mem_3Z0Z_4;
    wire sDAC_data_2_6_bm_1_7_cascade_;
    wire sDAC_data_RNO_15Z0Z_7;
    wire sDAC_mem_36Z0Z_5;
    wire sDAC_mem_37Z0Z_5;
    wire sDAC_data_2_13_am_1_8_cascade_;
    wire sDAC_mem_5Z0Z_5;
    wire sDAC_mem_4Z0Z_5;
    wire sDAC_mem_36Z0Z_6;
    wire sDAC_mem_37Z0Z_6;
    wire sDAC_data_2_13_am_1_9_cascade_;
    wire sDAC_mem_5Z0Z_6;
    wire sDAC_mem_4Z0Z_6;
    wire sDAC_mem_6Z0Z_7;
    wire sDAC_data_2_13_bm_1_10_cascade_;
    wire sDAC_mem_7Z0Z_7;
    wire sDAC_data_RNO_4Z0Z_9;
    wire sDAC_data_RNO_2Z0Z_9;
    wire sDAC_data_RNO_1Z0Z_9_cascade_;
    wire sDAC_data_2_9_cascade_;
    wire sDAC_dataZ0Z_9;
    wire sDAC_data_RNO_15Z0Z_9;
    wire sDAC_data_RNO_14Z0Z_9;
    wire sDAC_data_2_14_ns_1_9;
    wire sDAC_data_RNO_29Z0Z_9;
    wire sDAC_data_RNO_30Z0Z_9;
    wire sDAC_data_2_32_ns_1_9_cascade_;
    wire sDAC_data_RNO_20Z0Z_9;
    wire sDAC_data_RNO_10Z0Z_9_cascade_;
    wire sDAC_data_RNO_11Z0Z_9;
    wire sDAC_data_2_41_ns_1_9;
    wire sDAC_mem_2Z0Z_5;
    wire sDAC_mem_34Z0Z_5;
    wire sDAC_data_2_6_bm_1_8_cascade_;
    wire sDAC_mem_3Z0Z_5;
    wire sDAC_mem_33Z0Z_7;
    wire sDAC_data_RNO_26Z0Z_10_cascade_;
    wire sDAC_mem_1Z0Z_7;
    wire sDAC_mem_32Z0Z_7;
    wire sDAC_data_RNO_27Z0Z_10;
    wire sDAC_mem_1Z0Z_0;
    wire sDAC_mem_32Z0Z_0;
    wire sDAC_mem_33Z0Z_0;
    wire sDAC_data_RNO_26Z0Z_3_cascade_;
    wire sDAC_data_RNO_27Z0Z_3;
    wire sDAC_data_RNO_21Z0Z_10;
    wire sDAC_data_RNO_30Z0Z_10;
    wire sDAC_data_2_32_ns_1_10;
    wire sDAC_data_RNO_14Z0Z_10;
    wire sDAC_data_RNO_5Z0Z_10;
    wire sDAC_data_2_14_ns_1_10_cascade_;
    wire sDAC_data_RNO_10Z0Z_10;
    wire sDAC_data_RNO_2Z0Z_10;
    wire sDAC_data_2_41_ns_1_10_cascade_;
    wire sDAC_data_RNO_1Z0Z_10;
    wire sDAC_data_2_10_cascade_;
    wire sDAC_dataZ0Z_10;
    wire sDAC_mem_36Z0Z_7;
    wire sDAC_mem_37Z0Z_7;
    wire sDAC_data_2_13_am_1_10_cascade_;
    wire sDAC_mem_5Z0Z_7;
    wire sDAC_data_RNO_4Z0Z_10;
    wire sDAC_mem_4Z0Z_7;
    wire sDAC_mem_36Z0Z_0;
    wire sDAC_mem_37Z0Z_0;
    wire sDAC_data_2_13_am_1_3_cascade_;
    wire sDAC_mem_5Z0Z_0;
    wire sDAC_mem_4Z0Z_0;
    wire sDAC_mem_4_1_sqmuxa;
    wire sDAC_mem_36Z0Z_1;
    wire sDAC_mem_4Z0Z_1;
    wire sDAC_mem_37Z0Z_1;
    wire sDAC_data_2_13_am_1_4_cascade_;
    wire sDAC_mem_5Z0Z_1;
    wire sDAC_data_RNO_20Z0Z_10;
    wire sDAC_mem_26_1_sqmuxa;
    wire N_142_cascade_;
    wire sDAC_mem_30Z0Z_2;
    wire sDAC_mem_30Z0Z_3;
    wire sDAC_mem_30Z0Z_5;
    wire sDAC_mem_30Z0Z_6;
    wire sDAC_mem_30_1_sqmuxa;
    wire sDAC_mem_23Z0Z_5;
    wire sDAC_mem_22Z0Z_5;
    wire sDAC_mem_23Z0Z_6;
    wire sDAC_data_RNO_21Z0Z_9;
    wire sDAC_mem_22Z0Z_6;
    wire sDAC_mem_22_1_sqmuxa;
    wire sDAC_mem_29Z0Z_1;
    wire sDAC_mem_30Z0Z_1;
    wire sDAC_mem_31Z0Z_1;
    wire sDAC_mem_31Z0Z_4;
    wire sDAC_mem_30Z0Z_4;
    wire sDAC_data_RNO_24Z0Z_7;
    wire sDAC_data_RNO_31Z0Z_10_cascade_;
    wire sDAC_data_2_39_ns_1_10_cascade_;
    wire sDAC_data_RNO_11Z0Z_10;
    wire sDAC_mem_26Z0Z_7;
    wire sDAC_data_RNO_32Z0Z_10;
    wire sDAC_mem_29Z0Z_7;
    wire sDAC_data_RNO_23Z0Z_10;
    wire sDAC_mem_31Z0Z_7;
    wire sDAC_mem_30Z0Z_7;
    wire sDAC_data_RNO_24Z0Z_10;
    wire sDAC_mem_24Z0Z_7;
    wire sDAC_mem_24_1_sqmuxa;
    wire sDAC_data_RNO_32Z0Z_3;
    wire sDAC_data_RNO_31Z0Z_3;
    wire sDAC_mem_25Z0Z_4;
    wire sDAC_mem_25Z0Z_7;
    wire sDAC_mem_25Z0Z_2;
    wire sDAC_mem_25Z0Z_5;
    wire sDAC_mem_25Z0Z_0;
    wire sDAC_mem_25Z0Z_6;
    wire sDAC_mem_25Z0Z_3;
    wire sDAC_mem_34_1_sqmuxa;
    wire sDAC_mem_39Z0Z_0;
    wire sDAC_mem_39Z0Z_1;
    wire sDAC_mem_39Z0Z_2;
    wire sDAC_mem_39Z0Z_4;
    wire sDAC_mem_39Z0Z_7;
    wire sDAC_mem_37_1_sqmuxa;
    wire sDAC_mem_39_1_sqmuxa;
    wire sDAC_mem_36_1_sqmuxa;
    wire N_288;
    wire sAddressZ0Z_3;
    wire N_288_cascade_;
    wire sAddressZ0Z_0;
    wire sDAC_mem_35Z0Z_0;
    wire sDAC_mem_35Z0Z_2;
    wire sDAC_mem_35Z0Z_4;
    wire sDAC_mem_35Z0Z_5;
    wire sDAC_mem_35Z0Z_6;
    wire sDAC_mem_35_1_sqmuxa;
    wire sDAC_mem_21Z0Z_4;
    wire sDAC_mem_21Z0Z_5;
    wire sDAC_mem_21Z0Z_6;
    wire sDAC_mem_21Z0Z_7;
    wire sDAC_mem_21_1_sqmuxa;
    wire sDAC_mem_7Z0Z_3;
    wire sDAC_data_2_13_bm_1_6_cascade_;
    wire sDAC_mem_39Z0Z_3;
    wire sDAC_mem_6Z0Z_3;
    wire sDAC_mem_6Z0Z_4;
    wire sDAC_mem_6Z0Z_5;
    wire sDAC_mem_7Z0Z_5;
    wire sDAC_data_2_13_bm_1_8_cascade_;
    wire sDAC_mem_39Z0Z_5;
    wire sDAC_data_RNO_21Z0Z_8;
    wire sDAC_data_RNO_20Z0Z_8;
    wire sDAC_data_RNO_29Z0Z_8;
    wire sDAC_data_RNO_30Z0Z_8;
    wire sDAC_data_2_32_ns_1_8;
    wire sDAC_data_RNO_15Z0Z_8;
    wire sDAC_data_RNO_14Z0Z_8;
    wire sDAC_data_RNO_5Z0Z_8;
    wire sDAC_data_2_14_ns_1_8_cascade_;
    wire sDAC_data_RNO_4Z0Z_8;
    wire sDAC_data_RNO_10Z0Z_8;
    wire sDAC_data_RNO_11Z0Z_8;
    wire sDAC_data_2_41_ns_1_8_cascade_;
    wire sDAC_data_RNO_1Z0Z_8;
    wire sDAC_data_2_8_cascade_;
    wire sDAC_dataZ0Z_8;
    wire sDAC_mem_2Z0Z_1;
    wire sDAC_mem_34Z0Z_1;
    wire sDAC_mem_35Z0Z_1;
    wire sDAC_data_2_6_bm_1_4_cascade_;
    wire sDAC_mem_3Z0Z_1;
    wire sDAC_data_RNO_17Z0Z_6_cascade_;
    wire sDAC_mem_8Z0Z_3;
    wire sDAC_data_2_20_am_1_6_cascade_;
    wire sDAC_data_2_24_ns_1_6;
    wire sDAC_data_RNO_7Z0Z_6_cascade_;
    wire sDAC_data_RNO_8Z0Z_6;
    wire sDAC_data_RNO_10Z0Z_4_cascade_;
    wire sDAC_data_RNO_30Z0Z_4;
    wire sDAC_data_2_32_ns_1_4;
    wire sDAC_data_RNO_15Z0Z_4;
    wire sDAC_data_RNO_14Z0Z_4;
    wire sDAC_data_RNO_5Z0Z_4;
    wire sDAC_data_2_14_ns_1_4_cascade_;
    wire sDAC_data_RNO_4Z0Z_4;
    wire sDAC_data_RNO_1Z0Z_4_cascade_;
    wire sDAC_data_2_41_ns_1_4;
    wire sDAC_data_2_4_cascade_;
    wire sDAC_dataZ0Z_4;
    wire sDAC_data_RNO_21Z0Z_3;
    wire sDAC_data_RNO_10Z0Z_3_cascade_;
    wire sDAC_data_RNO_30Z0Z_3;
    wire sDAC_data_2_32_ns_1_3;
    wire sDAC_data_RNO_15Z0Z_3;
    wire sDAC_data_RNO_14Z0Z_3;
    wire sDAC_data_RNO_5Z0Z_3;
    wire sDAC_data_2_14_ns_1_3_cascade_;
    wire sDAC_data_RNO_4Z0Z_3;
    wire sDAC_data_RNO_1Z0Z_3_cascade_;
    wire sDAC_data_2_41_ns_1_3;
    wire sDAC_data_2_3_cascade_;
    wire sDAC_dataZ0Z_3;
    wire sDAC_mem_16Z0Z_7;
    wire sDAC_mem_17Z0Z_7;
    wire sDAC_data_RNO_29Z0Z_10;
    wire sDAC_mem_19Z0Z_3;
    wire sDAC_mem_18Z0Z_3;
    wire sDAC_mem_23Z0Z_1;
    wire sDAC_mem_22Z0Z_1;
    wire sDAC_data_RNO_21Z0Z_4;
    wire sDAC_mem_27Z0Z_2;
    wire sDAC_mem_27Z0Z_3;
    wire sDAC_mem_27Z0Z_4;
    wire sDAC_mem_27Z0Z_5;
    wire sDAC_mem_27Z0Z_6;
    wire sDAC_mem_27Z0Z_7;
    wire sEEADC_freqZ0Z_0;
    wire sEEADC_freqZ0Z_6;
    wire sEEADC_freqZ0Z_7;
    wire sDAC_mem_31Z0Z_0;
    wire sDAC_mem_30Z0Z_0;
    wire sDAC_mem_29Z0Z_0;
    wire sDAC_data_RNO_24Z0Z_3;
    wire sDAC_data_RNO_23Z0Z_3_cascade_;
    wire sDAC_data_2_39_ns_1_3;
    wire sDAC_data_RNO_11Z0Z_3;
    wire sDAC_mem_28Z0Z_0;
    wire sDAC_mem_24Z0Z_1;
    wire sDAC_data_RNO_31Z0Z_4_cascade_;
    wire sDAC_data_RNO_24Z0Z_4;
    wire sDAC_data_2_39_ns_1_4_cascade_;
    wire sDAC_data_RNO_23Z0Z_4;
    wire sDAC_data_RNO_11Z0Z_4;
    wire sDAC_mem_26Z0Z_1;
    wire sDAC_mem_27Z0Z_1;
    wire sDAC_data_RNO_32Z0Z_4;
    wire sDAC_mem_28Z0Z_1;
    wire sDAC_mem_28Z0Z_2;
    wire sDAC_mem_28Z0Z_4;
    wire sDAC_mem_28Z0Z_5;
    wire sDAC_mem_28Z0Z_7;
    wire sDAC_mem_28_1_sqmuxa;
    wire sDAC_mem_25Z0Z_1;
    wire sDAC_mem_25_1_sqmuxa;
    wire sDAC_mem_17Z0Z_1;
    wire sDAC_data_RNO_29Z0Z_4;
    wire sDAC_mem_38Z0Z_0;
    wire sDAC_mem_38Z0Z_2;
    wire sDAC_mem_38Z0Z_3;
    wire sDAC_mem_38Z0Z_4;
    wire sDAC_mem_38Z0Z_5;
    wire sDAC_mem_38Z0Z_7;
    wire sDAC_mem_38_1_sqmuxa;
    wire sDAC_mem_40Z0Z_2;
    wire sDAC_mem_40Z0Z_3;
    wire sDAC_mem_40Z0Z_4;
    wire sDAC_mem_40Z0Z_6;
    wire sDAC_mem_40Z0Z_7;
    wire sDAC_mem_40_1_sqmuxa;
    wire sDAC_mem_21Z0Z_0;
    wire sDAC_data_RNO_20Z0Z_3;
    wire sDAC_mem_20Z0Z_0;
    wire sDAC_mem_21Z0Z_1;
    wire sDAC_data_RNO_20Z0Z_4;
    wire sDAC_mem_20Z0Z_1;
    wire sDAC_mem_21Z0Z_2;
    wire sDAC_data_RNO_20Z0Z_5;
    wire sDAC_mem_20Z0Z_2;
    wire sDAC_mem_21Z0Z_3;
    wire sDAC_mem_20Z0Z_3;
    wire sDAC_mem_33Z0Z_3;
    wire sDAC_data_RNO_26Z0Z_6_cascade_;
    wire sDAC_mem_32Z0Z_3;
    wire sDAC_data_RNO_27Z0Z_6;
    wire sDAC_mem_1Z0Z_3;
    wire sDAC_mem_33Z0Z_4;
    wire sDAC_data_RNO_26Z0Z_7_cascade_;
    wire sDAC_data_RNO_14Z0Z_7;
    wire sDAC_mem_32Z0Z_4;
    wire sDAC_data_RNO_27Z0Z_7;
    wire sDAC_mem_1Z0Z_4;
    wire sDAC_mem_1_1_sqmuxa;
    wire sDAC_data_RNO_5Z0Z_6;
    wire sDAC_data_RNO_4Z0Z_6;
    wire sDAC_data_RNO_14Z0Z_6;
    wire sDAC_data_2_14_ns_1_6;
    wire sDAC_data_RNO_29Z0Z_6;
    wire sDAC_data_RNO_30Z0Z_6;
    wire sDAC_data_RNO_21Z0Z_6;
    wire sDAC_data_2_32_ns_1_6_cascade_;
    wire sDAC_data_RNO_20Z0Z_6;
    wire sDAC_mem_pointerZ0Z_3;
    wire sDAC_data_RNO_10Z0Z_6_cascade_;
    wire sDAC_data_RNO_11Z0Z_6;
    wire sDAC_mem_pointerZ0Z_4;
    wire sDAC_data_RNO_2Z0Z_6;
    wire sDAC_data_2_41_ns_1_6_cascade_;
    wire sDAC_data_RNO_1Z0Z_6;
    wire un5_sdacdyn_cry_23_c_RNIELGZ0Z28;
    wire sDAC_data_2_6_cascade_;
    wire sDAC_dataZ0Z_6;
    wire op_eq_scounterdac10_g;
    wire sDAC_mem_2Z0Z_3;
    wire sDAC_mem_34Z0Z_3;
    wire sDAC_mem_35Z0Z_3;
    wire sDAC_data_2_6_bm_1_6_cascade_;
    wire sDAC_mem_3Z0Z_3;
    wire sDAC_data_RNO_15Z0Z_6;
    wire sDAC_data_RNO_17Z0Z_8_cascade_;
    wire sDAC_mem_40Z0Z_5;
    wire sDAC_mem_8Z0Z_5;
    wire sDAC_data_2_20_am_1_8_cascade_;
    wire sDAC_data_RNO_7Z0Z_8_cascade_;
    wire sDAC_data_RNO_8Z0Z_8;
    wire sDAC_data_RNO_2Z0Z_8;
    wire sDAC_mem_38Z0Z_6;
    wire sDAC_mem_39Z0Z_6;
    wire sDAC_data_2_13_bm_1_9_cascade_;
    wire sDAC_mem_7Z0Z_6;
    wire sDAC_data_RNO_5Z0Z_9;
    wire sDAC_mem_6Z0Z_6;
    wire sDAC_mem_6_1_sqmuxa;
    wire sDAC_mem_40Z0Z_0;
    wire sDAC_mem_8Z0Z_0;
    wire sDAC_data_2_20_am_1_3_cascade_;
    wire sDAC_data_RNO_17Z0Z_3_cascade_;
    wire sDAC_data_RNO_8Z0Z_3_cascade_;
    wire sDAC_data_RNO_7Z0Z_3;
    wire sDAC_data_RNO_2Z0Z_3;
    wire sDAC_mem_3_1_sqmuxa;
    wire sDAC_mem_34Z0Z_7;
    wire sDAC_mem_2Z0Z_7;
    wire sDAC_mem_35Z0Z_7;
    wire sDAC_data_2_6_bm_1_10_cascade_;
    wire sDAC_mem_3Z0Z_7;
    wire sDAC_data_RNO_15Z0Z_10;
    wire sDAC_mem_40Z0Z_1;
    wire sDAC_mem_8Z0Z_1;
    wire sDAC_data_2_20_am_1_4_cascade_;
    wire sDAC_mem_pointerZ0Z_5;
    wire sDAC_data_RNO_17Z0Z_4_cascade_;
    wire sDAC_data_RNO_8Z0Z_4_cascade_;
    wire sDAC_data_RNO_7Z0Z_4;
    wire sDAC_data_RNO_2Z0Z_4;
    wire N_284_cascade_;
    wire N_284;
    wire N_280;
    wire sPointerZ0Z_1;
    wire un1_spointer11_0;
    wire sDAC_mem_14Z0Z_2;
    wire sDAC_mem_14Z0Z_3;
    wire sDAC_mem_14Z0Z_6;
    wire sDAC_mem_14_1_sqmuxa;
    wire sDAC_mem_14Z0Z_4;
    wire sDAC_data_RNO_18Z0Z_7_cascade_;
    wire sDAC_data_RNO_19Z0Z_7;
    wire sDAC_data_2_24_ns_1_7;
    wire sDAC_data_RNO_18Z0Z_8_cascade_;
    wire sDAC_data_2_24_ns_1_8;
    wire sDAC_mem_12Z0Z_4;
    wire sDAC_mem_14Z0Z_5;
    wire sDAC_data_RNO_19Z0Z_8;
    wire sDAC_mem_12Z0Z_5;
    wire sEEADC_freqZ0Z_1;
    wire sEEADC_freq_1_sqmuxa;
    wire sDAC_mem_17Z0Z_0;
    wire sDAC_mem_16Z0Z_0;
    wire sDAC_data_RNO_29Z0Z_3;
    wire sDAC_mem_16Z0Z_3;
    wire sDAC_mem_20Z0Z_7;
    wire sDAC_mem_20_1_sqmuxa;
    wire sDAC_mem_41Z0Z_0;
    wire sDAC_mem_41Z0Z_1;
    wire sDAC_mem_41Z0Z_2;
    wire sDAC_mem_41Z0Z_3;
    wire sDAC_mem_41Z0Z_4;
    wire sDAC_mem_41Z0Z_5;
    wire sDAC_mem_41Z0Z_6;
    wire sDAC_mem_41Z0Z_7;
    wire sDAC_mem_42Z0Z_0;
    wire sDAC_mem_42Z0Z_1;
    wire sDAC_mem_42Z0Z_2;
    wire sDAC_mem_42Z0Z_3;
    wire sDAC_mem_42Z0Z_4;
    wire sDAC_mem_42Z0Z_5;
    wire sDAC_mem_42Z0Z_6;
    wire sDAC_mem_42Z0Z_7;
    wire sDAC_mem_10Z0Z_0;
    wire sDAC_mem_10Z0Z_1;
    wire sDAC_mem_10Z0Z_2;
    wire sDAC_mem_10Z0Z_3;
    wire sDAC_mem_10Z0Z_4;
    wire sDAC_mem_10Z0Z_5;
    wire sDAC_mem_10Z0Z_6;
    wire sDAC_mem_10_1_sqmuxa;
    wire sDAC_mem_42_1_sqmuxa;
    wire sAddressZ0Z_2;
    wire sAddressZ0Z_1;
    wire sDAC_mem_30_1_sqmuxa_0_a2_1_0;
    wire N_275;
    wire sAddressZ0Z_4;
    wire N_286;
    wire N_278_cascade_;
    wire N_142;
    wire sDAC_mem_15Z0Z_2;
    wire sDAC_mem_15Z0Z_3;
    wire sDAC_mem_15Z0Z_4;
    wire sDAC_mem_15Z0Z_5;
    wire sDAC_mem_15Z0Z_6;
    wire sDAC_mem_15_1_sqmuxa;
    wire sDAC_mem_11Z0Z_0;
    wire sDAC_mem_11Z0Z_1;
    wire sDAC_mem_11Z0Z_2;
    wire sDAC_mem_11Z0Z_3;
    wire sDAC_mem_11Z0Z_4;
    wire sDAC_mem_11Z0Z_5;
    wire sDAC_mem_11Z0Z_6;
    wire sDAC_mem_11Z0Z_7;
    wire sDAC_mem_11_1_sqmuxa;
    wire sDAC_mem_15Z0Z_0;
    wire sDAC_mem_14Z0Z_0;
    wire sDAC_data_RNO_18Z0Z_3_cascade_;
    wire sDAC_data_RNO_19Z0Z_3;
    wire sDAC_data_2_24_ns_1_3;
    wire sDAC_mem_pointerZ0Z_2;
    wire sDAC_mem_pointerZ0Z_1;
    wire sDAC_data_RNO_18Z0Z_4_cascade_;
    wire sDAC_data_2_24_ns_1_4;
    wire sDAC_mem_12Z0Z_0;
    wire sDAC_mem_15Z0Z_1;
    wire sDAC_mem_14Z0Z_1;
    wire sDAC_data_RNO_19Z0Z_4;
    wire sDAC_mem_12Z0Z_1;
    wire sDAC_mem_27Z0Z_0;
    wire sDAC_mem_27_1_sqmuxa;
    wire sDAC_mem_13Z0Z_6;
    wire sDAC_mem_13Z0Z_5;
    wire sDAC_mem_16Z0Z_1;
    wire sDAC_mem_16_1_sqmuxa;
    wire sEEDACZ0Z_7;
    wire sAddressZ0Z_5;
    wire N_139;
    wire N_278;
    wire sDAC_mem_41_1_sqmuxa;
    wire N_285;
    wire N_1480;
    wire N_360;
    wire sEEDACZ0Z_0;
    wire sEEDACZ0Z_1;
    wire sEEDACZ0Z_2;
    wire sEEDACZ0Z_3;
    wire sEEDACZ0Z_4;
    wire sEEDACZ0Z_5;
    wire sEEDACZ0Z_6;
    wire sEEDAC_1_sqmuxa;
    wire sDAC_mem_9Z0Z_0;
    wire sDAC_mem_9Z0Z_1;
    wire sDAC_mem_9Z0Z_2;
    wire sDAC_mem_9Z0Z_3;
    wire sDAC_mem_9Z0Z_4;
    wire spi_data_mosi_5;
    wire sDAC_mem_9Z0Z_5;
    wire sDAC_mem_9Z0Z_6;
    wire sDAC_mem_9Z0Z_7;
    wire sDAC_mem_9_1_sqmuxa;
    wire N_14_3_cascade_;
    wire N_8_cascade_;
    wire sDAC_spi_startZ0;
    wire un1_scounterdac8_i_a2_1_2;
    wire un1_scounterdac8_i_a2_0;
    wire sDAC_data_RNO_18Z0Z_10;
    wire sDAC_mem_pointerZ0Z_0;
    wire sDAC_mem_15Z0Z_7;
    wire sDAC_mem_14Z0Z_7;
    wire sDAC_data_RNO_19Z0Z_10;
    wire spi_data_mosi_0;
    wire sDAC_mem_13Z0Z_0;
    wire spi_data_mosi_1;
    wire sDAC_mem_13Z0Z_1;
    wire spi_data_mosi_2;
    wire sDAC_mem_13Z0Z_2;
    wire spi_data_mosi_3;
    wire sDAC_mem_13Z0Z_3;
    wire spi_data_mosi_4;
    wire sDAC_mem_13Z0Z_4;
    wire sDAC_mem_13Z0Z_7;
    wire sDAC_mem_13_1_sqmuxa;
    wire spi_data_mosi_7;
    wire sDAC_mem_12Z0Z_7;
    wire spi_data_mosi_6;
    wire sDAC_mem_12Z0Z_6;
    wire pll_clk128_g;
    wire sDAC_mem_12_1_sqmuxa;
    wire N_14_3;
    wire bfn_22_10_0_;
    wire un2_scounterdac_cry_1;
    wire sCounterDACZ0Z_3;
    wire un2_scounterdac_cry_2;
    wire un2_scounterdac_cry_3;
    wire sCounterDACZ0Z_5;
    wire un2_scounterdac_cry_4;
    wire un2_scounterdac_cry_5_THRU_CO;
    wire un2_scounterdac_cry_5;
    wire un2_scounterdac_cry_6;
    wire sCounterDACZ0Z_8;
    wire un2_scounterdac_cry_7_THRU_CO;
    wire un2_scounterdac_cry_7;
    wire un2_scounterdac_cry_8;
    wire bfn_22_11_0_;
    wire pll_clk64_0_g;
    wire LED3_c_i_g;
    wire spi_mosi_rpi_c;
    wire spi_mosi_flash_c;
    wire sCounterDACZ0Z_4;
    wire sCounterDACZ0Z_1;
    wire sCounterDACZ0Z_7;
    wire sCounterDACZ0Z_2;
    wire sCounterDACZ0Z_9;
    wire sCounterDACZ0Z_6;
    wire spi_cs_rpi_c;
    wire spi_cs_flash_c;
    wire spi_sclk_rpi_c;
    wire cs_rpi2flash_c;
    wire spi_sclk_flash_c;
    wire op_eq_scounterdac10_0_a2_0;
    wire N_23;
    wire sCounterDACZ0Z_0;
    wire N_22;
    wire op_eq_scounterdac10;
    wire _gnd_net_;

    defparam \pll128M2_inst.pll128M2_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll128M2_inst.pll128M2_inst .TEST_MODE=1'b0;
    defparam \pll128M2_inst.pll128M2_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll128M2_inst.pll128M2_inst .PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam \pll128M2_inst.pll128M2_inst .PLLOUT_SELECT_PORTA="GENCLK";
    defparam \pll128M2_inst.pll128M2_inst .FILTER_RANGE=3'b001;
    defparam \pll128M2_inst.pll128M2_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll128M2_inst.pll128M2_inst .FDA_RELATIVE=4'b0000;
    defparam \pll128M2_inst.pll128M2_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll128M2_inst.pll128M2_inst .ENABLE_ICEGATE_PORTB=1'b0;
    defparam \pll128M2_inst.pll128M2_inst .ENABLE_ICEGATE_PORTA=1'b0;
    defparam \pll128M2_inst.pll128M2_inst .DIVR=4'b0000;
    defparam \pll128M2_inst.pll128M2_inst .DIVQ=3'b011;
    defparam \pll128M2_inst.pll128M2_inst .DIVF=7'b1010100;
    defparam \pll128M2_inst.pll128M2_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE \pll128M2_inst.pll128M2_inst  (
            .EXTFEEDBACK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(\pll128M2_inst.pll_clk64_0 ),
            .REFERENCECLK(N__20538),
            .RESETB(N__32326),
            .BYPASS(GNDG0),
            .PLLOUTCOREA(\pll128M2_inst.pll_clk128 ),
            .SDI(GNDG0),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(GNDG0),
            .PLLOUTGLOBALA(),
            .SCLK(GNDG0));
    IO_PAD RAM_ADD_obuf_5_iopad (
            .OE(N__54196),
            .DIN(N__54195),
            .DOUT(N__54194),
            .PACKAGEPIN(RAM_ADD[5]));
    defparam RAM_ADD_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_5_preio (
            .PADOEN(N__54196),
            .PADOUT(N__54195),
            .PADIN(N__54194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28581),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_mosi_rpi_ibuf_iopad (
            .OE(N__54187),
            .DIN(N__54186),
            .DOUT(N__54185),
            .PACKAGEPIN(spi_mosi_rpi));
    defparam spi_mosi_rpi_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_mosi_rpi_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_mosi_rpi_ibuf_preio (
            .PADOEN(N__54187),
            .PADOUT(N__54186),
            .PADIN(N__54185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_mosi_rpi_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_sclk_rpi_ibuf_iopad (
            .OE(N__54178),
            .DIN(N__54177),
            .DOUT(N__54176),
            .PACKAGEPIN(spi_sclk_rpi));
    defparam spi_sclk_rpi_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_sclk_rpi_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_sclk_rpi_ibuf_preio (
            .PADOEN(N__54178),
            .PADOUT(N__54177),
            .PADIN(N__54176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_sclk_rpi_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_miso_ft_obuf_iopad (
            .OE(N__54169),
            .DIN(N__54168),
            .DOUT(N__54167),
            .PACKAGEPIN(spi_miso_ft));
    defparam spi_miso_ft_obuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_miso_ft_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO spi_miso_ft_obuf_preio (
            .PADOEN(N__54169),
            .PADOUT(N__54168),
            .PADIN(N__54167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__38490),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC5_ibuf_iopad (
            .OE(N__54160),
            .DIN(N__54159),
            .DOUT(N__54158),
            .PACKAGEPIN(ADC5));
    defparam ADC5_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC5_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC5_ibuf_preio (
            .PADOEN(N__54160),
            .PADOUT(N__54159),
            .PADIN(N__54158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC5_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_ACQ_obuf_iopad (
            .OE(N__54151),
            .DIN(N__54150),
            .DOUT(N__54149),
            .PACKAGEPIN(LED_ACQ));
    defparam LED_ACQ_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED_ACQ_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_ACQ_obuf_preio (
            .PADOEN(N__54151),
            .PADOUT(N__54150),
            .PADIN(N__54149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22260),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD reset_rpi_ibuf_iopad (
            .OE(N__54142),
            .DIN(N__54141),
            .DOUT(N__54140),
            .PACKAGEPIN(reset_rpi));
    defparam reset_rpi_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam reset_rpi_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_rpi_ibuf_preio (
            .PADOEN(N__54142),
            .PADOUT(N__54141),
            .PADIN(N__54140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(LED3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_6_iopad (
            .OE(N__54133),
            .DIN(N__54132),
            .DOUT(N__54131),
            .PACKAGEPIN(RAM_DATA[6]));
    defparam RAM_DATA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_6_preio (
            .PADOEN(N__54133),
            .PADOUT(N__54132),
            .PADIN(N__54131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__30558),
            .DIN0(RAM_DATA_in_6),
            .DOUT0(N__31539),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_9_iopad (
            .OE(N__54124),
            .DIN(N__54123),
            .DOUT(N__54122),
            .PACKAGEPIN(RAM_ADD[9]));
    defparam RAM_ADD_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_9_preio (
            .PADOEN(N__54124),
            .PADOUT(N__54123),
            .PADIN(N__54122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28392),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_11_iopad (
            .OE(N__54115),
            .DIN(N__54114),
            .DOUT(N__54113),
            .PACKAGEPIN(RAM_DATA[11]));
    defparam RAM_DATA_iobuf_11_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_11_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_11_preio (
            .PADOEN(N__54115),
            .PADOUT(N__54114),
            .PADIN(N__54113),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__31773),
            .DIN0(RAM_DATA_in_11),
            .DOUT0(N__31455),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD trig_rpi_ibuf_iopad (
            .OE(N__54106),
            .DIN(N__54105),
            .DOUT(N__54104),
            .PACKAGEPIN(trig_rpi));
    defparam trig_rpi_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam trig_rpi_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO trig_rpi_ibuf_preio (
            .PADOEN(N__54106),
            .PADOUT(N__54105),
            .PADIN(N__54104),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(trig_rpi_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_0_iopad (
            .OE(N__54097),
            .DIN(N__54096),
            .DOUT(N__54095),
            .PACKAGEPIN(RAM_DATA[0]));
    defparam RAM_DATA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_0_preio (
            .PADOEN(N__54097),
            .PADOUT(N__54096),
            .PADIN(N__54095),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__26865),
            .DIN0(RAM_DATA_in_0),
            .DOUT0(N__30186),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC2_ibuf_iopad (
            .OE(N__54088),
            .DIN(N__54087),
            .DOUT(N__54086),
            .PACKAGEPIN(ADC2));
    defparam ADC2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC2_ibuf_preio (
            .PADOEN(N__54088),
            .PADOUT(N__54087),
            .PADIN(N__54086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_18_iopad (
            .OE(N__54079),
            .DIN(N__54078),
            .DOUT(N__54077),
            .PACKAGEPIN(RAM_ADD[18]));
    defparam RAM_ADD_obuf_18_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_18_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_18_preio (
            .PADOEN(N__54079),
            .PADOUT(N__54078),
            .PADIN(N__54077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28098),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_2_iopad (
            .OE(N__54070),
            .DIN(N__54069),
            .DOUT(N__54068),
            .PACKAGEPIN(RAM_ADD[2]));
    defparam RAM_ADD_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_2_preio (
            .PADOEN(N__54070),
            .PADOUT(N__54069),
            .PADIN(N__54068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28056),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DAC_mosi_obuf_iopad (
            .OE(N__54061),
            .DIN(N__54060),
            .DOUT(N__54059),
            .PACKAGEPIN(DAC_mosi));
    defparam DAC_mosi_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DAC_mosi_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DAC_mosi_obuf_preio (
            .PADOEN(N__54061),
            .PADOUT(N__54060),
            .PADIN(N__54059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21147),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_13_iopad (
            .OE(N__54052),
            .DIN(N__54051),
            .DOUT(N__54050),
            .PACKAGEPIN(RAM_ADD[13]));
    defparam RAM_ADD_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_13_preio (
            .PADOEN(N__54052),
            .PADOUT(N__54051),
            .PADIN(N__54050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__30291),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_nWE_obuf_iopad (
            .OE(N__54043),
            .DIN(N__54042),
            .DOUT(N__54041),
            .PACKAGEPIN(RAM_nWE));
    defparam RAM_nWE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAM_nWE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_nWE_obuf_preio (
            .PADOEN(N__54043),
            .PADOUT(N__54042),
            .PADIN(N__54041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27660),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_7_iopad (
            .OE(N__54034),
            .DIN(N__54033),
            .DOUT(N__54032),
            .PACKAGEPIN(RAM_DATA[7]));
    defparam RAM_DATA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_7_preio (
            .PADOEN(N__54034),
            .PADOUT(N__54033),
            .PADIN(N__54032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__30486),
            .DIN0(RAM_DATA_in_7),
            .DOUT0(N__30579),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC0_ibuf_iopad (
            .OE(N__54025),
            .DIN(N__54024),
            .DOUT(N__54023),
            .PACKAGEPIN(ADC0));
    defparam ADC0_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC0_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC0_ibuf_preio (
            .PADOEN(N__54025),
            .PADOUT(N__54024),
            .PADIN(N__54023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC0_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_nLB_obuf_iopad (
            .OE(N__54016),
            .DIN(N__54015),
            .DOUT(N__54014),
            .PACKAGEPIN(RAM_nLB));
    defparam RAM_nLB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAM_nLB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_nLB_obuf_preio (
            .PADOEN(N__54016),
            .PADOUT(N__54015),
            .PADIN(N__54014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_10_iopad (
            .OE(N__54007),
            .DIN(N__54006),
            .DOUT(N__54005),
            .PACKAGEPIN(RAM_DATA[10]));
    defparam RAM_DATA_iobuf_10_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_10_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_10_preio (
            .PADOEN(N__54007),
            .PADOUT(N__54006),
            .PADIN(N__54005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__31746),
            .DIN0(RAM_DATA_in_10),
            .DOUT0(N__31500),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_1_iopad (
            .OE(N__53998),
            .DIN(N__53997),
            .DOUT(N__53996),
            .PACKAGEPIN(RAM_DATA[1]));
    defparam RAM_DATA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_1_preio (
            .PADOEN(N__53998),
            .PADOUT(N__53997),
            .PADIN(N__53996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__28326),
            .DIN0(RAM_DATA_in_1),
            .DOUT0(N__30105),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_select_ibuf_iopad (
            .OE(N__53989),
            .DIN(N__53988),
            .DOUT(N__53987),
            .PACKAGEPIN(spi_select));
    defparam spi_select_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_select_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_select_ibuf_preio (
            .PADOEN(N__53989),
            .PADOUT(N__53988),
            .PADIN(N__53987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_select_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_nCE_obuf_iopad (
            .OE(N__53980),
            .DIN(N__53979),
            .DOUT(N__53978),
            .PACKAGEPIN(RAM_nCE));
    defparam RAM_nCE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAM_nCE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_nCE_obuf_preio (
            .PADOEN(N__53980),
            .PADOUT(N__53979),
            .PADIN(N__53978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_sclk_flash_obuf_iopad (
            .OE(N__53971),
            .DIN(N__53970),
            .DOUT(N__53969),
            .PACKAGEPIN(spi_sclk_flash));
    defparam spi_sclk_flash_obuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_sclk_flash_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO spi_sclk_flash_obuf_preio (
            .PADOEN(N__53971),
            .PADOUT(N__53970),
            .PADIN(N__53969),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__52272),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_3_iopad (
            .OE(N__53962),
            .DIN(N__53961),
            .DOUT(N__53960),
            .PACKAGEPIN(RAM_ADD[3]));
    defparam RAM_ADD_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_3_preio (
            .PADOEN(N__53962),
            .PADOUT(N__53961),
            .PADIN(N__53960),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28662),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_12_iopad (
            .OE(N__53953),
            .DIN(N__53952),
            .DOUT(N__53951),
            .PACKAGEPIN(RAM_ADD[12]));
    defparam RAM_ADD_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_12_preio (
            .PADOEN(N__53953),
            .PADOUT(N__53952),
            .PADIN(N__53951),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__30327),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC3_ibuf_iopad (
            .OE(N__53944),
            .DIN(N__53943),
            .DOUT(N__53942),
            .PACKAGEPIN(ADC3));
    defparam ADC3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC3_ibuf_preio (
            .PADOEN(N__53944),
            .PADOUT(N__53943),
            .PADIN(N__53942),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_15_iopad (
            .OE(N__53935),
            .DIN(N__53934),
            .DOUT(N__53933),
            .PACKAGEPIN(RAM_DATA[15]));
    defparam RAM_DATA_iobuf_15_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_15_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_15_preio (
            .PADOEN(N__53935),
            .PADOUT(N__53934),
            .PADIN(N__53933),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__32721),
            .DIN0(RAM_DATA_in_15),
            .DOUT0(N__30600),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pon_obuf_iopad (
            .OE(N__53926),
            .DIN(N__53925),
            .DOUT(N__53924),
            .PACKAGEPIN(pon));
    defparam pon_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pon_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pon_obuf_preio (
            .PADOEN(N__53926),
            .PADOUT(N__53925),
            .PADIN(N__53924),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21918),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DAC_sclk_obuf_iopad (
            .OE(N__53917),
            .DIN(N__53916),
            .DOUT(N__53915),
            .PACKAGEPIN(DAC_sclk));
    defparam DAC_sclk_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DAC_sclk_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DAC_sclk_obuf_preio (
            .PADOEN(N__53917),
            .PADOUT(N__53916),
            .PADIN(N__53915),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21069),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_4_iopad (
            .OE(N__53908),
            .DIN(N__53907),
            .DOUT(N__53906),
            .PACKAGEPIN(RAM_DATA[4]));
    defparam RAM_DATA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_4_preio (
            .PADOEN(N__53908),
            .PADOUT(N__53907),
            .PADIN(N__53906),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__27822),
            .DIN0(RAM_DATA_in_4),
            .DOUT0(N__31572),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC1_ibuf_iopad (
            .OE(N__53899),
            .DIN(N__53898),
            .DOUT(N__53897),
            .PACKAGEPIN(ADC1));
    defparam ADC1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC1_ibuf_preio (
            .PADOEN(N__53899),
            .PADOUT(N__53898),
            .PADIN(N__53897),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_cs_flash_obuf_iopad (
            .OE(N__53890),
            .DIN(N__53889),
            .DOUT(N__53888),
            .PACKAGEPIN(spi_cs_flash));
    defparam spi_cs_flash_obuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_cs_flash_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO spi_cs_flash_obuf_preio (
            .PADOEN(N__53890),
            .PADOUT(N__53889),
            .PADIN(N__53888),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__52362),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_miso_flash_ibuf_iopad (
            .OE(N__53881),
            .DIN(N__53880),
            .DOUT(N__53879),
            .PACKAGEPIN(spi_miso_flash));
    defparam spi_miso_flash_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_miso_flash_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_miso_flash_ibuf_preio (
            .PADOEN(N__53881),
            .PADOUT(N__53880),
            .PADIN(N__53879),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_miso_flash_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD trig_ext_ibuf_iopad (
            .OE(N__53872),
            .DIN(N__53871),
            .DOUT(N__53870),
            .PACKAGEPIN(trig_ext));
    defparam trig_ext_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam trig_ext_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO trig_ext_ibuf_preio (
            .PADOEN(N__53872),
            .PADOUT(N__53871),
            .PADIN(N__53870),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(trig_ext_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_6_iopad (
            .OE(N__53863),
            .DIN(N__53862),
            .DOUT(N__53861),
            .PACKAGEPIN(RAM_ADD[6]));
    defparam RAM_ADD_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_6_preio (
            .PADOEN(N__53863),
            .PADOUT(N__53862),
            .PADIN(N__53861),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28536),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD top_tour1_ibuf_iopad (
            .OE(N__53854),
            .DIN(N__53853),
            .DOUT(N__53852),
            .PACKAGEPIN(top_tour1));
    defparam top_tour1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam top_tour1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO top_tour1_ibuf_preio (
            .PADOEN(N__53854),
            .PADOUT(N__53853),
            .PADIN(N__53852),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(top_tour1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_17_iopad (
            .OE(N__53845),
            .DIN(N__53844),
            .DOUT(N__53843),
            .PACKAGEPIN(RAM_ADD[17]));
    defparam RAM_ADD_obuf_17_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_17_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_17_preio (
            .PADOEN(N__53845),
            .PADOUT(N__53844),
            .PADIN(N__53843),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28140),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_0_iopad (
            .OE(N__53836),
            .DIN(N__53835),
            .DOUT(N__53834),
            .PACKAGEPIN(RAM_ADD[0]));
    defparam RAM_ADD_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_0_preio (
            .PADOEN(N__53836),
            .PADOUT(N__53835),
            .PADIN(N__53834),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29739),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED_MODE_obuf_iopad (
            .OE(N__53827),
            .DIN(N__53826),
            .DOUT(N__53825),
            .PACKAGEPIN(LED_MODE));
    defparam LED_MODE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED_MODE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_MODE_obuf_preio (
            .PADOEN(N__53827),
            .PADOUT(N__53826),
            .PADIN(N__53825),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24321),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_nUB_obuf_iopad (
            .OE(N__53818),
            .DIN(N__53817),
            .DOUT(N__53816),
            .PACKAGEPIN(RAM_nUB));
    defparam RAM_nUB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAM_nUB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_nUB_obuf_preio (
            .PADOEN(N__53818),
            .PADOUT(N__53817),
            .PADIN(N__53816),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_11_iopad (
            .OE(N__53809),
            .DIN(N__53808),
            .DOUT(N__53807),
            .PACKAGEPIN(RAM_ADD[11]));
    defparam RAM_ADD_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_11_preio (
            .PADOEN(N__53809),
            .PADOUT(N__53808),
            .PADIN(N__53807),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__30381),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_14_iopad (
            .OE(N__53800),
            .DIN(N__53799),
            .DOUT(N__53798),
            .PACKAGEPIN(RAM_DATA[14]));
    defparam RAM_DATA_iobuf_14_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_14_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_14_preio (
            .PADOEN(N__53800),
            .PADOUT(N__53799),
            .PADIN(N__53798),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__32754),
            .DIN0(RAM_DATA_in_14),
            .DOUT0(N__31230),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DAC_cs_obuf_iopad (
            .OE(N__53791),
            .DIN(N__53790),
            .DOUT(N__53789),
            .PACKAGEPIN(DAC_cs));
    defparam DAC_cs_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DAC_cs_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DAC_cs_obuf_preio (
            .PADOEN(N__53791),
            .PADOUT(N__53790),
            .PADIN(N__53789),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20574),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC8_ibuf_iopad (
            .OE(N__53782),
            .DIN(N__53781),
            .DOUT(N__53780),
            .PACKAGEPIN(ADC8));
    defparam ADC8_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC8_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC8_ibuf_preio (
            .PADOEN(N__53782),
            .PADOUT(N__53781),
            .PADIN(N__53780),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC8_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_5_iopad (
            .OE(N__53773),
            .DIN(N__53772),
            .DOUT(N__53771),
            .PACKAGEPIN(RAM_DATA[5]));
    defparam RAM_DATA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_5_preio (
            .PADOEN(N__53773),
            .PADOUT(N__53772),
            .PADIN(N__53771),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__26931),
            .DIN0(RAM_DATA_in_5),
            .DOUT0(N__30147),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC_clk_obuf_iopad (
            .OE(N__53764),
            .DIN(N__53763),
            .DOUT(N__53762),
            .PACKAGEPIN(ADC_clk));
    defparam ADC_clk_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC_clk_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ADC_clk_obuf_preio (
            .PADOEN(N__53764),
            .PADOUT(N__53763),
            .PADIN(N__53762),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27615),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_7_iopad (
            .OE(N__53755),
            .DIN(N__53754),
            .DOUT(N__53753),
            .PACKAGEPIN(RAM_ADD[7]));
    defparam RAM_ADD_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_7_preio (
            .PADOEN(N__53755),
            .PADOUT(N__53754),
            .PADIN(N__53753),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28488),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD poff_obuf_iopad (
            .OE(N__53746),
            .DIN(N__53745),
            .DOUT(N__53744),
            .PACKAGEPIN(poff));
    defparam poff_obuf_preio.NEG_TRIGGER=1'b0;
    defparam poff_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO poff_obuf_preio (
            .PADOEN(N__53746),
            .PADOUT(N__53745),
            .PADIN(N__53744),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25335),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC4_ibuf_iopad (
            .OE(N__53737),
            .DIN(N__53736),
            .DOUT(N__53735),
            .PACKAGEPIN(ADC4));
    defparam ADC4_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC4_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC4_ibuf_preio (
            .PADOEN(N__53737),
            .PADOUT(N__53736),
            .PADIN(N__53735),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC4_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC6_ibuf_iopad (
            .OE(N__53728),
            .DIN(N__53727),
            .DOUT(N__53726),
            .PACKAGEPIN(ADC6));
    defparam ADC6_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC6_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC6_ibuf_preio (
            .PADOEN(N__53728),
            .PADOUT(N__53727),
            .PADIN(N__53726),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC6_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_16_iopad (
            .OE(N__53719),
            .DIN(N__53718),
            .DOUT(N__53717),
            .PACKAGEPIN(RAM_ADD[16]));
    defparam RAM_ADD_obuf_16_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_16_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_16_preio (
            .PADOEN(N__53719),
            .PADOUT(N__53718),
            .PADIN(N__53717),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28185),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_1_iopad (
            .OE(N__53710),
            .DIN(N__53709),
            .DOUT(N__53708),
            .PACKAGEPIN(RAM_ADD[1]));
    defparam RAM_ADD_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_1_preio (
            .PADOEN(N__53710),
            .PADOUT(N__53709),
            .PADIN(N__53708),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29664),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC7_ibuf_iopad (
            .OE(N__53701),
            .DIN(N__53700),
            .DOUT(N__53699),
            .PACKAGEPIN(ADC7));
    defparam ADC7_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC7_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC7_ibuf_preio (
            .PADOEN(N__53701),
            .PADOUT(N__53700),
            .PADIN(N__53699),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC7_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD button_mode_ibuf_iopad (
            .OE(N__53692),
            .DIN(N__53691),
            .DOUT(N__53690),
            .PACKAGEPIN(button_mode));
    defparam button_mode_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam button_mode_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO button_mode_ibuf_preio (
            .PADOEN(N__53692),
            .PADOUT(N__53691),
            .PADIN(N__53690),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(button_mode_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_sclk_ft_ibuf_iopad (
            .OE(N__53683),
            .DIN(N__53682),
            .DOUT(N__53681),
            .PACKAGEPIN(spi_sclk_ft));
    defparam spi_sclk_ft_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_sclk_ft_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_sclk_ft_ibuf_preio (
            .PADOEN(N__53683),
            .PADOUT(N__53682),
            .PADIN(N__53681),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_sclk_ft_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_8_iopad (
            .OE(N__53674),
            .DIN(N__53673),
            .DOUT(N__53672),
            .PACKAGEPIN(RAM_DATA[8]));
    defparam RAM_DATA_iobuf_8_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_8_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_8_preio (
            .PADOEN(N__53674),
            .PADOUT(N__53673),
            .PADIN(N__53672),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__26646),
            .DIN0(RAM_DATA_in_8),
            .DOUT0(N__30075),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_10_iopad (
            .OE(N__53665),
            .DIN(N__53664),
            .DOUT(N__53663),
            .PACKAGEPIN(RAM_ADD[10]));
    defparam RAM_ADD_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_10_preio (
            .PADOEN(N__53665),
            .PADOUT(N__53664),
            .PADIN(N__53663),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29616),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_13_iopad (
            .OE(N__53656),
            .DIN(N__53655),
            .DOUT(N__53654),
            .PACKAGEPIN(RAM_DATA[13]));
    defparam RAM_DATA_iobuf_13_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_13_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_13_preio (
            .PADOEN(N__53656),
            .PADOUT(N__53655),
            .PADIN(N__53654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__30522),
            .DIN0(RAM_DATA_in_13),
            .DOUT0(N__31317),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD trig_ft_ibuf_iopad (
            .OE(N__53647),
            .DIN(N__53646),
            .DOUT(N__53645),
            .PACKAGEPIN(trig_ft));
    defparam trig_ft_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam trig_ft_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO trig_ft_ibuf_preio (
            .PADOEN(N__53647),
            .PADOUT(N__53646),
            .PADIN(N__53645),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(trig_ft_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADC9_ibuf_iopad (
            .OE(N__53638),
            .DIN(N__53637),
            .DOUT(N__53636),
            .PACKAGEPIN(ADC9));
    defparam ADC9_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ADC9_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ADC9_ibuf_preio (
            .PADOEN(N__53638),
            .PADOUT(N__53637),
            .PADIN(N__53636),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ADC9_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_2_iopad (
            .OE(N__53629),
            .DIN(N__53628),
            .DOUT(N__53627),
            .PACKAGEPIN(RAM_DATA[2]));
    defparam RAM_DATA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_2_preio (
            .PADOEN(N__53629),
            .PADOUT(N__53628),
            .PADIN(N__53627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__30447),
            .DIN0(RAM_DATA_in_2),
            .DOUT0(N__31197),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD cs_rpi2flash_ibuf_iopad (
            .OE(N__53620),
            .DIN(N__53619),
            .DOUT(N__53618),
            .PACKAGEPIN(cs_rpi2flash));
    defparam cs_rpi2flash_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam cs_rpi2flash_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO cs_rpi2flash_ibuf_preio (
            .PADOEN(N__53620),
            .PADOUT(N__53619),
            .PADIN(N__53618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(cs_rpi2flash_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED3_obuf_iopad (
            .OE(N__53611),
            .DIN(N__53610),
            .DOUT(N__53609),
            .PACKAGEPIN(LED3));
    defparam LED3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED3_obuf_preio (
            .PADOEN(N__53611),
            .PADOUT(N__53610),
            .PADIN(N__53609),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32583),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_mosi_ft_ibuf_iopad (
            .OE(N__53602),
            .DIN(N__53601),
            .DOUT(N__53600),
            .PACKAGEPIN(spi_mosi_ft));
    defparam spi_mosi_ft_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_mosi_ft_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_mosi_ft_ibuf_preio (
            .PADOEN(N__53602),
            .PADOUT(N__53601),
            .PADIN(N__53600),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_mosi_ft_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_nOE_obuf_iopad (
            .OE(N__53593),
            .DIN(N__53592),
            .DOUT(N__53591),
            .PACKAGEPIN(RAM_nOE));
    defparam RAM_nOE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAM_nOE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_nOE_obuf_preio (
            .PADOEN(N__53593),
            .PADOUT(N__53592),
            .PADIN(N__53591),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_4_iopad (
            .OE(N__53584),
            .DIN(N__53583),
            .DOUT(N__53582),
            .PACKAGEPIN(RAM_ADD[4]));
    defparam RAM_ADD_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_4_preio (
            .PADOEN(N__53584),
            .PADOUT(N__53583),
            .PADIN(N__53582),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28626),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_ibuf_iopad (
            .OE(N__53575),
            .DIN(N__53574),
            .DOUT(N__53573),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_preio (
            .PADOEN(N__53575),
            .PADOUT(N__53574),
            .PADIN(N__53573),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD top_tour2_ibuf_iopad (
            .OE(N__53566),
            .DIN(N__53565),
            .DOUT(N__53564),
            .PACKAGEPIN(top_tour2));
    defparam top_tour2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam top_tour2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO top_tour2_ibuf_preio (
            .PADOEN(N__53566),
            .PADOUT(N__53565),
            .PADIN(N__53564),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(top_tour2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_cs_rpi_ibuf_iopad (
            .OE(N__53557),
            .DIN(N__53556),
            .DOUT(N__53555),
            .PACKAGEPIN(spi_cs_rpi));
    defparam spi_cs_rpi_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_cs_rpi_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_cs_rpi_ibuf_preio (
            .PADOEN(N__53557),
            .PADOUT(N__53556),
            .PADIN(N__53555),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_cs_rpi_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_15_iopad (
            .OE(N__53548),
            .DIN(N__53547),
            .DOUT(N__53546),
            .PACKAGEPIN(RAM_ADD[15]));
    defparam RAM_ADD_obuf_15_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_15_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_15_preio (
            .PADOEN(N__53548),
            .PADOUT(N__53547),
            .PADIN(N__53546),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28230),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_miso_rpi_obuf_iopad (
            .OE(N__53539),
            .DIN(N__53538),
            .DOUT(N__53537),
            .PACKAGEPIN(spi_miso_rpi));
    defparam spi_miso_rpi_obuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_miso_rpi_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO spi_miso_rpi_obuf_preio (
            .PADOEN(N__53539),
            .PADOUT(N__53538),
            .PADIN(N__53537),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33120),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_9_iopad (
            .OE(N__53530),
            .DIN(N__53529),
            .DOUT(N__53528),
            .PACKAGEPIN(RAM_DATA[9]));
    defparam RAM_DATA_iobuf_9_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_9_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_9_preio (
            .PADOEN(N__53530),
            .PADOUT(N__53529),
            .PADIN(N__53528),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__28362),
            .DIN0(RAM_DATA_in_9),
            .DOUT0(N__30624),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_8_iopad (
            .OE(N__53521),
            .DIN(N__53520),
            .DOUT(N__53519),
            .PACKAGEPIN(RAM_ADD[8]));
    defparam RAM_ADD_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_8_preio (
            .PADOEN(N__53521),
            .PADOUT(N__53520),
            .PADIN(N__53519),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28440),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_12_iopad (
            .OE(N__53512),
            .DIN(N__53511),
            .DOUT(N__53510),
            .PACKAGEPIN(RAM_DATA[12]));
    defparam RAM_DATA_iobuf_12_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_12_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_12_preio (
            .PADOEN(N__53512),
            .PADOUT(N__53511),
            .PADIN(N__53510),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__26898),
            .DIN0(RAM_DATA_in_12),
            .DOUT0(N__31413),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_DATA_iobuf_3_iopad (
            .OE(N__53503),
            .DIN(N__53502),
            .DOUT(N__53501),
            .PACKAGEPIN(RAM_DATA[3]));
    defparam RAM_DATA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam RAM_DATA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO RAM_DATA_iobuf_3_preio (
            .PADOEN(N__53503),
            .PADOUT(N__53502),
            .PADIN(N__53501),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__27792),
            .DIN0(RAM_DATA_in_3),
            .DOUT0(N__30222),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_cs_ft_ibuf_iopad (
            .OE(N__53494),
            .DIN(N__53493),
            .DOUT(N__53492),
            .PACKAGEPIN(spi_cs_ft));
    defparam spi_cs_ft_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_cs_ft_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO spi_cs_ft_ibuf_preio (
            .PADOEN(N__53494),
            .PADOUT(N__53493),
            .PADIN(N__53492),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(spi_cs_ft_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD spi_mosi_flash_obuf_iopad (
            .OE(N__53485),
            .DIN(N__53484),
            .DOUT(N__53483),
            .PACKAGEPIN(spi_mosi_flash));
    defparam spi_mosi_flash_obuf_preio.NEG_TRIGGER=1'b0;
    defparam spi_mosi_flash_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO spi_mosi_flash_obuf_preio (
            .PADOEN(N__53485),
            .PADOUT(N__53484),
            .PADIN(N__53483),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__52563),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAM_ADD_obuf_14_iopad (
            .OE(N__53476),
            .DIN(N__53475),
            .DOUT(N__53474),
            .PACKAGEPIN(RAM_ADD[14]));
    defparam RAM_ADD_obuf_14_preio.NEG_TRIGGER=1'b0;
    defparam RAM_ADD_obuf_14_preio.PIN_TYPE=6'b011001;
    PRE_IO RAM_ADD_obuf_14_preio (
            .PADOEN(N__53476),
            .PADOUT(N__53475),
            .PADIN(N__53474),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28275),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__12722 (
            .O(N__53457),
            .I(N__53454));
    LocalMux I__12721 (
            .O(N__53454),
            .I(op_eq_scounterdac10_0_a2_0));
    InMux I__12720 (
            .O(N__53451),
            .I(N__53446));
    InMux I__12719 (
            .O(N__53450),
            .I(N__53443));
    InMux I__12718 (
            .O(N__53449),
            .I(N__53440));
    LocalMux I__12717 (
            .O(N__53446),
            .I(N__53437));
    LocalMux I__12716 (
            .O(N__53443),
            .I(N__53433));
    LocalMux I__12715 (
            .O(N__53440),
            .I(N__53430));
    Span4Mux_v I__12714 (
            .O(N__53437),
            .I(N__53427));
    InMux I__12713 (
            .O(N__53436),
            .I(N__53424));
    Odrv4 I__12712 (
            .O(N__53433),
            .I(N_23));
    Odrv4 I__12711 (
            .O(N__53430),
            .I(N_23));
    Odrv4 I__12710 (
            .O(N__53427),
            .I(N_23));
    LocalMux I__12709 (
            .O(N__53424),
            .I(N_23));
    CascadeMux I__12708 (
            .O(N__53415),
            .I(N__53411));
    CascadeMux I__12707 (
            .O(N__53414),
            .I(N__53407));
    InMux I__12706 (
            .O(N__53411),
            .I(N__53402));
    InMux I__12705 (
            .O(N__53410),
            .I(N__53399));
    InMux I__12704 (
            .O(N__53407),
            .I(N__53396));
    InMux I__12703 (
            .O(N__53406),
            .I(N__53390));
    InMux I__12702 (
            .O(N__53405),
            .I(N__53390));
    LocalMux I__12701 (
            .O(N__53402),
            .I(N__53387));
    LocalMux I__12700 (
            .O(N__53399),
            .I(N__53382));
    LocalMux I__12699 (
            .O(N__53396),
            .I(N__53382));
    CascadeMux I__12698 (
            .O(N__53395),
            .I(N__53379));
    LocalMux I__12697 (
            .O(N__53390),
            .I(N__53372));
    Span4Mux_v I__12696 (
            .O(N__53387),
            .I(N__53372));
    Span4Mux_v I__12695 (
            .O(N__53382),
            .I(N__53372));
    InMux I__12694 (
            .O(N__53379),
            .I(N__53369));
    Odrv4 I__12693 (
            .O(N__53372),
            .I(sCounterDACZ0Z_0));
    LocalMux I__12692 (
            .O(N__53369),
            .I(sCounterDACZ0Z_0));
    InMux I__12691 (
            .O(N__53364),
            .I(N__53361));
    LocalMux I__12690 (
            .O(N__53361),
            .I(N__53358));
    Span4Mux_v I__12689 (
            .O(N__53358),
            .I(N__53354));
    InMux I__12688 (
            .O(N__53357),
            .I(N__53351));
    Odrv4 I__12687 (
            .O(N__53354),
            .I(N_22));
    LocalMux I__12686 (
            .O(N__53351),
            .I(N_22));
    IoInMux I__12685 (
            .O(N__53346),
            .I(N__53343));
    LocalMux I__12684 (
            .O(N__53343),
            .I(N__53340));
    Odrv12 I__12683 (
            .O(N__53340),
            .I(op_eq_scounterdac10));
    InMux I__12682 (
            .O(N__53337),
            .I(N__53332));
    InMux I__12681 (
            .O(N__53336),
            .I(N__53326));
    InMux I__12680 (
            .O(N__53335),
            .I(N__53326));
    LocalMux I__12679 (
            .O(N__53332),
            .I(N__53323));
    InMux I__12678 (
            .O(N__53331),
            .I(N__53319));
    LocalMux I__12677 (
            .O(N__53326),
            .I(N__53316));
    Span12Mux_h I__12676 (
            .O(N__53323),
            .I(N__53313));
    InMux I__12675 (
            .O(N__53322),
            .I(N__53310));
    LocalMux I__12674 (
            .O(N__53319),
            .I(N__53305));
    Span4Mux_h I__12673 (
            .O(N__53316),
            .I(N__53305));
    Odrv12 I__12672 (
            .O(N__53313),
            .I(sCounterDACZ0Z_8));
    LocalMux I__12671 (
            .O(N__53310),
            .I(sCounterDACZ0Z_8));
    Odrv4 I__12670 (
            .O(N__53305),
            .I(sCounterDACZ0Z_8));
    InMux I__12669 (
            .O(N__53298),
            .I(N__53295));
    LocalMux I__12668 (
            .O(N__53295),
            .I(N__53292));
    Odrv4 I__12667 (
            .O(N__53292),
            .I(un2_scounterdac_cry_7_THRU_CO));
    InMux I__12666 (
            .O(N__53289),
            .I(un2_scounterdac_cry_7));
    InMux I__12665 (
            .O(N__53286),
            .I(bfn_22_11_0_));
    ClkMux I__12664 (
            .O(N__53283),
            .I(N__53154));
    ClkMux I__12663 (
            .O(N__53282),
            .I(N__53154));
    ClkMux I__12662 (
            .O(N__53281),
            .I(N__53154));
    ClkMux I__12661 (
            .O(N__53280),
            .I(N__53154));
    ClkMux I__12660 (
            .O(N__53279),
            .I(N__53154));
    ClkMux I__12659 (
            .O(N__53278),
            .I(N__53154));
    ClkMux I__12658 (
            .O(N__53277),
            .I(N__53154));
    ClkMux I__12657 (
            .O(N__53276),
            .I(N__53154));
    ClkMux I__12656 (
            .O(N__53275),
            .I(N__53154));
    ClkMux I__12655 (
            .O(N__53274),
            .I(N__53154));
    ClkMux I__12654 (
            .O(N__53273),
            .I(N__53154));
    ClkMux I__12653 (
            .O(N__53272),
            .I(N__53154));
    ClkMux I__12652 (
            .O(N__53271),
            .I(N__53154));
    ClkMux I__12651 (
            .O(N__53270),
            .I(N__53154));
    ClkMux I__12650 (
            .O(N__53269),
            .I(N__53154));
    ClkMux I__12649 (
            .O(N__53268),
            .I(N__53154));
    ClkMux I__12648 (
            .O(N__53267),
            .I(N__53154));
    ClkMux I__12647 (
            .O(N__53266),
            .I(N__53154));
    ClkMux I__12646 (
            .O(N__53265),
            .I(N__53154));
    ClkMux I__12645 (
            .O(N__53264),
            .I(N__53154));
    ClkMux I__12644 (
            .O(N__53263),
            .I(N__53154));
    ClkMux I__12643 (
            .O(N__53262),
            .I(N__53154));
    ClkMux I__12642 (
            .O(N__53261),
            .I(N__53154));
    ClkMux I__12641 (
            .O(N__53260),
            .I(N__53154));
    ClkMux I__12640 (
            .O(N__53259),
            .I(N__53154));
    ClkMux I__12639 (
            .O(N__53258),
            .I(N__53154));
    ClkMux I__12638 (
            .O(N__53257),
            .I(N__53154));
    ClkMux I__12637 (
            .O(N__53256),
            .I(N__53154));
    ClkMux I__12636 (
            .O(N__53255),
            .I(N__53154));
    ClkMux I__12635 (
            .O(N__53254),
            .I(N__53154));
    ClkMux I__12634 (
            .O(N__53253),
            .I(N__53154));
    ClkMux I__12633 (
            .O(N__53252),
            .I(N__53154));
    ClkMux I__12632 (
            .O(N__53251),
            .I(N__53154));
    ClkMux I__12631 (
            .O(N__53250),
            .I(N__53154));
    ClkMux I__12630 (
            .O(N__53249),
            .I(N__53154));
    ClkMux I__12629 (
            .O(N__53248),
            .I(N__53154));
    ClkMux I__12628 (
            .O(N__53247),
            .I(N__53154));
    ClkMux I__12627 (
            .O(N__53246),
            .I(N__53154));
    ClkMux I__12626 (
            .O(N__53245),
            .I(N__53154));
    ClkMux I__12625 (
            .O(N__53244),
            .I(N__53154));
    ClkMux I__12624 (
            .O(N__53243),
            .I(N__53154));
    ClkMux I__12623 (
            .O(N__53242),
            .I(N__53154));
    ClkMux I__12622 (
            .O(N__53241),
            .I(N__53154));
    GlobalMux I__12621 (
            .O(N__53154),
            .I(N__53151));
    gio2CtrlBuf I__12620 (
            .O(N__53151),
            .I(pll_clk64_0_g));
    SRMux I__12619 (
            .O(N__53148),
            .I(N__52602));
    SRMux I__12618 (
            .O(N__53147),
            .I(N__52602));
    SRMux I__12617 (
            .O(N__53146),
            .I(N__52602));
    SRMux I__12616 (
            .O(N__53145),
            .I(N__52602));
    SRMux I__12615 (
            .O(N__53144),
            .I(N__52602));
    SRMux I__12614 (
            .O(N__53143),
            .I(N__52602));
    SRMux I__12613 (
            .O(N__53142),
            .I(N__52602));
    SRMux I__12612 (
            .O(N__53141),
            .I(N__52602));
    SRMux I__12611 (
            .O(N__53140),
            .I(N__52602));
    SRMux I__12610 (
            .O(N__53139),
            .I(N__52602));
    SRMux I__12609 (
            .O(N__53138),
            .I(N__52602));
    SRMux I__12608 (
            .O(N__53137),
            .I(N__52602));
    SRMux I__12607 (
            .O(N__53136),
            .I(N__52602));
    SRMux I__12606 (
            .O(N__53135),
            .I(N__52602));
    SRMux I__12605 (
            .O(N__53134),
            .I(N__52602));
    SRMux I__12604 (
            .O(N__53133),
            .I(N__52602));
    SRMux I__12603 (
            .O(N__53132),
            .I(N__52602));
    SRMux I__12602 (
            .O(N__53131),
            .I(N__52602));
    SRMux I__12601 (
            .O(N__53130),
            .I(N__52602));
    SRMux I__12600 (
            .O(N__53129),
            .I(N__52602));
    SRMux I__12599 (
            .O(N__53128),
            .I(N__52602));
    SRMux I__12598 (
            .O(N__53127),
            .I(N__52602));
    SRMux I__12597 (
            .O(N__53126),
            .I(N__52602));
    SRMux I__12596 (
            .O(N__53125),
            .I(N__52602));
    SRMux I__12595 (
            .O(N__53124),
            .I(N__52602));
    SRMux I__12594 (
            .O(N__53123),
            .I(N__52602));
    SRMux I__12593 (
            .O(N__53122),
            .I(N__52602));
    SRMux I__12592 (
            .O(N__53121),
            .I(N__52602));
    SRMux I__12591 (
            .O(N__53120),
            .I(N__52602));
    SRMux I__12590 (
            .O(N__53119),
            .I(N__52602));
    SRMux I__12589 (
            .O(N__53118),
            .I(N__52602));
    SRMux I__12588 (
            .O(N__53117),
            .I(N__52602));
    SRMux I__12587 (
            .O(N__53116),
            .I(N__52602));
    SRMux I__12586 (
            .O(N__53115),
            .I(N__52602));
    SRMux I__12585 (
            .O(N__53114),
            .I(N__52602));
    SRMux I__12584 (
            .O(N__53113),
            .I(N__52602));
    SRMux I__12583 (
            .O(N__53112),
            .I(N__52602));
    SRMux I__12582 (
            .O(N__53111),
            .I(N__52602));
    SRMux I__12581 (
            .O(N__53110),
            .I(N__52602));
    SRMux I__12580 (
            .O(N__53109),
            .I(N__52602));
    SRMux I__12579 (
            .O(N__53108),
            .I(N__52602));
    SRMux I__12578 (
            .O(N__53107),
            .I(N__52602));
    SRMux I__12577 (
            .O(N__53106),
            .I(N__52602));
    SRMux I__12576 (
            .O(N__53105),
            .I(N__52602));
    SRMux I__12575 (
            .O(N__53104),
            .I(N__52602));
    SRMux I__12574 (
            .O(N__53103),
            .I(N__52602));
    SRMux I__12573 (
            .O(N__53102),
            .I(N__52602));
    SRMux I__12572 (
            .O(N__53101),
            .I(N__52602));
    SRMux I__12571 (
            .O(N__53100),
            .I(N__52602));
    SRMux I__12570 (
            .O(N__53099),
            .I(N__52602));
    SRMux I__12569 (
            .O(N__53098),
            .I(N__52602));
    SRMux I__12568 (
            .O(N__53097),
            .I(N__52602));
    SRMux I__12567 (
            .O(N__53096),
            .I(N__52602));
    SRMux I__12566 (
            .O(N__53095),
            .I(N__52602));
    SRMux I__12565 (
            .O(N__53094),
            .I(N__52602));
    SRMux I__12564 (
            .O(N__53093),
            .I(N__52602));
    SRMux I__12563 (
            .O(N__53092),
            .I(N__52602));
    SRMux I__12562 (
            .O(N__53091),
            .I(N__52602));
    SRMux I__12561 (
            .O(N__53090),
            .I(N__52602));
    SRMux I__12560 (
            .O(N__53089),
            .I(N__52602));
    SRMux I__12559 (
            .O(N__53088),
            .I(N__52602));
    SRMux I__12558 (
            .O(N__53087),
            .I(N__52602));
    SRMux I__12557 (
            .O(N__53086),
            .I(N__52602));
    SRMux I__12556 (
            .O(N__53085),
            .I(N__52602));
    SRMux I__12555 (
            .O(N__53084),
            .I(N__52602));
    SRMux I__12554 (
            .O(N__53083),
            .I(N__52602));
    SRMux I__12553 (
            .O(N__53082),
            .I(N__52602));
    SRMux I__12552 (
            .O(N__53081),
            .I(N__52602));
    SRMux I__12551 (
            .O(N__53080),
            .I(N__52602));
    SRMux I__12550 (
            .O(N__53079),
            .I(N__52602));
    SRMux I__12549 (
            .O(N__53078),
            .I(N__52602));
    SRMux I__12548 (
            .O(N__53077),
            .I(N__52602));
    SRMux I__12547 (
            .O(N__53076),
            .I(N__52602));
    SRMux I__12546 (
            .O(N__53075),
            .I(N__52602));
    SRMux I__12545 (
            .O(N__53074),
            .I(N__52602));
    SRMux I__12544 (
            .O(N__53073),
            .I(N__52602));
    SRMux I__12543 (
            .O(N__53072),
            .I(N__52602));
    SRMux I__12542 (
            .O(N__53071),
            .I(N__52602));
    SRMux I__12541 (
            .O(N__53070),
            .I(N__52602));
    SRMux I__12540 (
            .O(N__53069),
            .I(N__52602));
    SRMux I__12539 (
            .O(N__53068),
            .I(N__52602));
    SRMux I__12538 (
            .O(N__53067),
            .I(N__52602));
    SRMux I__12537 (
            .O(N__53066),
            .I(N__52602));
    SRMux I__12536 (
            .O(N__53065),
            .I(N__52602));
    SRMux I__12535 (
            .O(N__53064),
            .I(N__52602));
    SRMux I__12534 (
            .O(N__53063),
            .I(N__52602));
    SRMux I__12533 (
            .O(N__53062),
            .I(N__52602));
    SRMux I__12532 (
            .O(N__53061),
            .I(N__52602));
    SRMux I__12531 (
            .O(N__53060),
            .I(N__52602));
    SRMux I__12530 (
            .O(N__53059),
            .I(N__52602));
    SRMux I__12529 (
            .O(N__53058),
            .I(N__52602));
    SRMux I__12528 (
            .O(N__53057),
            .I(N__52602));
    SRMux I__12527 (
            .O(N__53056),
            .I(N__52602));
    SRMux I__12526 (
            .O(N__53055),
            .I(N__52602));
    SRMux I__12525 (
            .O(N__53054),
            .I(N__52602));
    SRMux I__12524 (
            .O(N__53053),
            .I(N__52602));
    SRMux I__12523 (
            .O(N__53052),
            .I(N__52602));
    SRMux I__12522 (
            .O(N__53051),
            .I(N__52602));
    SRMux I__12521 (
            .O(N__53050),
            .I(N__52602));
    SRMux I__12520 (
            .O(N__53049),
            .I(N__52602));
    SRMux I__12519 (
            .O(N__53048),
            .I(N__52602));
    SRMux I__12518 (
            .O(N__53047),
            .I(N__52602));
    SRMux I__12517 (
            .O(N__53046),
            .I(N__52602));
    SRMux I__12516 (
            .O(N__53045),
            .I(N__52602));
    SRMux I__12515 (
            .O(N__53044),
            .I(N__52602));
    SRMux I__12514 (
            .O(N__53043),
            .I(N__52602));
    SRMux I__12513 (
            .O(N__53042),
            .I(N__52602));
    SRMux I__12512 (
            .O(N__53041),
            .I(N__52602));
    SRMux I__12511 (
            .O(N__53040),
            .I(N__52602));
    SRMux I__12510 (
            .O(N__53039),
            .I(N__52602));
    SRMux I__12509 (
            .O(N__53038),
            .I(N__52602));
    SRMux I__12508 (
            .O(N__53037),
            .I(N__52602));
    SRMux I__12507 (
            .O(N__53036),
            .I(N__52602));
    SRMux I__12506 (
            .O(N__53035),
            .I(N__52602));
    SRMux I__12505 (
            .O(N__53034),
            .I(N__52602));
    SRMux I__12504 (
            .O(N__53033),
            .I(N__52602));
    SRMux I__12503 (
            .O(N__53032),
            .I(N__52602));
    SRMux I__12502 (
            .O(N__53031),
            .I(N__52602));
    SRMux I__12501 (
            .O(N__53030),
            .I(N__52602));
    SRMux I__12500 (
            .O(N__53029),
            .I(N__52602));
    SRMux I__12499 (
            .O(N__53028),
            .I(N__52602));
    SRMux I__12498 (
            .O(N__53027),
            .I(N__52602));
    SRMux I__12497 (
            .O(N__53026),
            .I(N__52602));
    SRMux I__12496 (
            .O(N__53025),
            .I(N__52602));
    SRMux I__12495 (
            .O(N__53024),
            .I(N__52602));
    SRMux I__12494 (
            .O(N__53023),
            .I(N__52602));
    SRMux I__12493 (
            .O(N__53022),
            .I(N__52602));
    SRMux I__12492 (
            .O(N__53021),
            .I(N__52602));
    SRMux I__12491 (
            .O(N__53020),
            .I(N__52602));
    SRMux I__12490 (
            .O(N__53019),
            .I(N__52602));
    SRMux I__12489 (
            .O(N__53018),
            .I(N__52602));
    SRMux I__12488 (
            .O(N__53017),
            .I(N__52602));
    SRMux I__12487 (
            .O(N__53016),
            .I(N__52602));
    SRMux I__12486 (
            .O(N__53015),
            .I(N__52602));
    SRMux I__12485 (
            .O(N__53014),
            .I(N__52602));
    SRMux I__12484 (
            .O(N__53013),
            .I(N__52602));
    SRMux I__12483 (
            .O(N__53012),
            .I(N__52602));
    SRMux I__12482 (
            .O(N__53011),
            .I(N__52602));
    SRMux I__12481 (
            .O(N__53010),
            .I(N__52602));
    SRMux I__12480 (
            .O(N__53009),
            .I(N__52602));
    SRMux I__12479 (
            .O(N__53008),
            .I(N__52602));
    SRMux I__12478 (
            .O(N__53007),
            .I(N__52602));
    SRMux I__12477 (
            .O(N__53006),
            .I(N__52602));
    SRMux I__12476 (
            .O(N__53005),
            .I(N__52602));
    SRMux I__12475 (
            .O(N__53004),
            .I(N__52602));
    SRMux I__12474 (
            .O(N__53003),
            .I(N__52602));
    SRMux I__12473 (
            .O(N__53002),
            .I(N__52602));
    SRMux I__12472 (
            .O(N__53001),
            .I(N__52602));
    SRMux I__12471 (
            .O(N__53000),
            .I(N__52602));
    SRMux I__12470 (
            .O(N__52999),
            .I(N__52602));
    SRMux I__12469 (
            .O(N__52998),
            .I(N__52602));
    SRMux I__12468 (
            .O(N__52997),
            .I(N__52602));
    SRMux I__12467 (
            .O(N__52996),
            .I(N__52602));
    SRMux I__12466 (
            .O(N__52995),
            .I(N__52602));
    SRMux I__12465 (
            .O(N__52994),
            .I(N__52602));
    SRMux I__12464 (
            .O(N__52993),
            .I(N__52602));
    SRMux I__12463 (
            .O(N__52992),
            .I(N__52602));
    SRMux I__12462 (
            .O(N__52991),
            .I(N__52602));
    SRMux I__12461 (
            .O(N__52990),
            .I(N__52602));
    SRMux I__12460 (
            .O(N__52989),
            .I(N__52602));
    SRMux I__12459 (
            .O(N__52988),
            .I(N__52602));
    SRMux I__12458 (
            .O(N__52987),
            .I(N__52602));
    SRMux I__12457 (
            .O(N__52986),
            .I(N__52602));
    SRMux I__12456 (
            .O(N__52985),
            .I(N__52602));
    SRMux I__12455 (
            .O(N__52984),
            .I(N__52602));
    SRMux I__12454 (
            .O(N__52983),
            .I(N__52602));
    SRMux I__12453 (
            .O(N__52982),
            .I(N__52602));
    SRMux I__12452 (
            .O(N__52981),
            .I(N__52602));
    SRMux I__12451 (
            .O(N__52980),
            .I(N__52602));
    SRMux I__12450 (
            .O(N__52979),
            .I(N__52602));
    SRMux I__12449 (
            .O(N__52978),
            .I(N__52602));
    SRMux I__12448 (
            .O(N__52977),
            .I(N__52602));
    SRMux I__12447 (
            .O(N__52976),
            .I(N__52602));
    SRMux I__12446 (
            .O(N__52975),
            .I(N__52602));
    SRMux I__12445 (
            .O(N__52974),
            .I(N__52602));
    SRMux I__12444 (
            .O(N__52973),
            .I(N__52602));
    SRMux I__12443 (
            .O(N__52972),
            .I(N__52602));
    SRMux I__12442 (
            .O(N__52971),
            .I(N__52602));
    SRMux I__12441 (
            .O(N__52970),
            .I(N__52602));
    SRMux I__12440 (
            .O(N__52969),
            .I(N__52602));
    SRMux I__12439 (
            .O(N__52968),
            .I(N__52602));
    SRMux I__12438 (
            .O(N__52967),
            .I(N__52602));
    GlobalMux I__12437 (
            .O(N__52602),
            .I(N__52599));
    gio2CtrlBuf I__12436 (
            .O(N__52599),
            .I(LED3_c_i_g));
    InMux I__12435 (
            .O(N__52596),
            .I(N__52593));
    LocalMux I__12434 (
            .O(N__52593),
            .I(N__52589));
    InMux I__12433 (
            .O(N__52592),
            .I(N__52586));
    Span4Mux_v I__12432 (
            .O(N__52589),
            .I(N__52583));
    LocalMux I__12431 (
            .O(N__52586),
            .I(N__52580));
    Sp12to4 I__12430 (
            .O(N__52583),
            .I(N__52577));
    Span4Mux_v I__12429 (
            .O(N__52580),
            .I(N__52574));
    Span12Mux_h I__12428 (
            .O(N__52577),
            .I(N__52569));
    Sp12to4 I__12427 (
            .O(N__52574),
            .I(N__52569));
    Span12Mux_h I__12426 (
            .O(N__52569),
            .I(N__52566));
    Odrv12 I__12425 (
            .O(N__52566),
            .I(spi_mosi_rpi_c));
    IoInMux I__12424 (
            .O(N__52563),
            .I(N__52560));
    LocalMux I__12423 (
            .O(N__52560),
            .I(N__52557));
    Span4Mux_s2_v I__12422 (
            .O(N__52557),
            .I(N__52554));
    Span4Mux_v I__12421 (
            .O(N__52554),
            .I(N__52551));
    Odrv4 I__12420 (
            .O(N__52551),
            .I(spi_mosi_flash_c));
    InMux I__12419 (
            .O(N__52548),
            .I(N__52542));
    InMux I__12418 (
            .O(N__52547),
            .I(N__52542));
    LocalMux I__12417 (
            .O(N__52542),
            .I(N__52537));
    InMux I__12416 (
            .O(N__52541),
            .I(N__52534));
    InMux I__12415 (
            .O(N__52540),
            .I(N__52531));
    Odrv4 I__12414 (
            .O(N__52537),
            .I(sCounterDACZ0Z_4));
    LocalMux I__12413 (
            .O(N__52534),
            .I(sCounterDACZ0Z_4));
    LocalMux I__12412 (
            .O(N__52531),
            .I(sCounterDACZ0Z_4));
    InMux I__12411 (
            .O(N__52524),
            .I(N__52521));
    LocalMux I__12410 (
            .O(N__52521),
            .I(N__52516));
    InMux I__12409 (
            .O(N__52520),
            .I(N__52513));
    InMux I__12408 (
            .O(N__52519),
            .I(N__52508));
    Span4Mux_v I__12407 (
            .O(N__52516),
            .I(N__52503));
    LocalMux I__12406 (
            .O(N__52513),
            .I(N__52503));
    InMux I__12405 (
            .O(N__52512),
            .I(N__52500));
    InMux I__12404 (
            .O(N__52511),
            .I(N__52497));
    LocalMux I__12403 (
            .O(N__52508),
            .I(sCounterDACZ0Z_1));
    Odrv4 I__12402 (
            .O(N__52503),
            .I(sCounterDACZ0Z_1));
    LocalMux I__12401 (
            .O(N__52500),
            .I(sCounterDACZ0Z_1));
    LocalMux I__12400 (
            .O(N__52497),
            .I(sCounterDACZ0Z_1));
    InMux I__12399 (
            .O(N__52488),
            .I(N__52484));
    InMux I__12398 (
            .O(N__52487),
            .I(N__52481));
    LocalMux I__12397 (
            .O(N__52484),
            .I(sCounterDACZ0Z_7));
    LocalMux I__12396 (
            .O(N__52481),
            .I(sCounterDACZ0Z_7));
    InMux I__12395 (
            .O(N__52476),
            .I(N__52472));
    InMux I__12394 (
            .O(N__52475),
            .I(N__52469));
    LocalMux I__12393 (
            .O(N__52472),
            .I(sCounterDACZ0Z_2));
    LocalMux I__12392 (
            .O(N__52469),
            .I(sCounterDACZ0Z_2));
    CascadeMux I__12391 (
            .O(N__52464),
            .I(N__52460));
    InMux I__12390 (
            .O(N__52463),
            .I(N__52457));
    InMux I__12389 (
            .O(N__52460),
            .I(N__52454));
    LocalMux I__12388 (
            .O(N__52457),
            .I(sCounterDACZ0Z_9));
    LocalMux I__12387 (
            .O(N__52454),
            .I(sCounterDACZ0Z_9));
    CascadeMux I__12386 (
            .O(N__52449),
            .I(N__52446));
    InMux I__12385 (
            .O(N__52446),
            .I(N__52441));
    InMux I__12384 (
            .O(N__52445),
            .I(N__52438));
    InMux I__12383 (
            .O(N__52444),
            .I(N__52435));
    LocalMux I__12382 (
            .O(N__52441),
            .I(N__52430));
    LocalMux I__12381 (
            .O(N__52438),
            .I(N__52430));
    LocalMux I__12380 (
            .O(N__52435),
            .I(sCounterDACZ0Z_6));
    Odrv12 I__12379 (
            .O(N__52430),
            .I(sCounterDACZ0Z_6));
    InMux I__12378 (
            .O(N__52425),
            .I(N__52422));
    LocalMux I__12377 (
            .O(N__52422),
            .I(N__52416));
    InMux I__12376 (
            .O(N__52421),
            .I(N__52407));
    InMux I__12375 (
            .O(N__52420),
            .I(N__52407));
    InMux I__12374 (
            .O(N__52419),
            .I(N__52407));
    Span4Mux_h I__12373 (
            .O(N__52416),
            .I(N__52404));
    InMux I__12372 (
            .O(N__52415),
            .I(N__52401));
    InMux I__12371 (
            .O(N__52414),
            .I(N__52398));
    LocalMux I__12370 (
            .O(N__52407),
            .I(N__52395));
    Sp12to4 I__12369 (
            .O(N__52404),
            .I(N__52390));
    LocalMux I__12368 (
            .O(N__52401),
            .I(N__52390));
    LocalMux I__12367 (
            .O(N__52398),
            .I(N__52387));
    Span12Mux_v I__12366 (
            .O(N__52395),
            .I(N__52384));
    Span12Mux_v I__12365 (
            .O(N__52390),
            .I(N__52381));
    Span4Mux_v I__12364 (
            .O(N__52387),
            .I(N__52378));
    Span12Mux_h I__12363 (
            .O(N__52384),
            .I(N__52375));
    Span12Mux_h I__12362 (
            .O(N__52381),
            .I(N__52372));
    Span4Mux_v I__12361 (
            .O(N__52378),
            .I(N__52369));
    Odrv12 I__12360 (
            .O(N__52375),
            .I(spi_cs_rpi_c));
    Odrv12 I__12359 (
            .O(N__52372),
            .I(spi_cs_rpi_c));
    Odrv4 I__12358 (
            .O(N__52369),
            .I(spi_cs_rpi_c));
    IoInMux I__12357 (
            .O(N__52362),
            .I(N__52359));
    LocalMux I__12356 (
            .O(N__52359),
            .I(N__52356));
    Span4Mux_s2_v I__12355 (
            .O(N__52356),
            .I(N__52353));
    Span4Mux_v I__12354 (
            .O(N__52353),
            .I(N__52350));
    Odrv4 I__12353 (
            .O(N__52350),
            .I(spi_cs_flash_c));
    InMux I__12352 (
            .O(N__52347),
            .I(N__52344));
    LocalMux I__12351 (
            .O(N__52344),
            .I(N__52340));
    InMux I__12350 (
            .O(N__52343),
            .I(N__52337));
    Span4Mux_v I__12349 (
            .O(N__52340),
            .I(N__52334));
    LocalMux I__12348 (
            .O(N__52337),
            .I(N__52331));
    Sp12to4 I__12347 (
            .O(N__52334),
            .I(N__52328));
    Span4Mux_v I__12346 (
            .O(N__52331),
            .I(N__52325));
    Span12Mux_h I__12345 (
            .O(N__52328),
            .I(N__52320));
    Sp12to4 I__12344 (
            .O(N__52325),
            .I(N__52320));
    Span12Mux_h I__12343 (
            .O(N__52320),
            .I(N__52317));
    Odrv12 I__12342 (
            .O(N__52317),
            .I(spi_sclk_rpi_c));
    InMux I__12341 (
            .O(N__52314),
            .I(N__52311));
    LocalMux I__12340 (
            .O(N__52311),
            .I(N__52308));
    Span4Mux_h I__12339 (
            .O(N__52308),
            .I(N__52305));
    Span4Mux_h I__12338 (
            .O(N__52305),
            .I(N__52301));
    InMux I__12337 (
            .O(N__52304),
            .I(N__52298));
    Span4Mux_h I__12336 (
            .O(N__52301),
            .I(N__52291));
    LocalMux I__12335 (
            .O(N__52298),
            .I(N__52291));
    InMux I__12334 (
            .O(N__52297),
            .I(N__52288));
    InMux I__12333 (
            .O(N__52296),
            .I(N__52285));
    Sp12to4 I__12332 (
            .O(N__52291),
            .I(N__52278));
    LocalMux I__12331 (
            .O(N__52288),
            .I(N__52278));
    LocalMux I__12330 (
            .O(N__52285),
            .I(N__52278));
    Span12Mux_v I__12329 (
            .O(N__52278),
            .I(N__52275));
    Odrv12 I__12328 (
            .O(N__52275),
            .I(cs_rpi2flash_c));
    IoInMux I__12327 (
            .O(N__52272),
            .I(N__52269));
    LocalMux I__12326 (
            .O(N__52269),
            .I(N__52266));
    Span12Mux_s6_v I__12325 (
            .O(N__52266),
            .I(N__52263));
    Odrv12 I__12324 (
            .O(N__52263),
            .I(spi_sclk_flash_c));
    CascadeMux I__12323 (
            .O(N__52260),
            .I(N__52257));
    InMux I__12322 (
            .O(N__52257),
            .I(N__52254));
    LocalMux I__12321 (
            .O(N__52254),
            .I(N__52250));
    CascadeMux I__12320 (
            .O(N__52253),
            .I(N__52247));
    Span4Mux_v I__12319 (
            .O(N__52250),
            .I(N__52244));
    InMux I__12318 (
            .O(N__52247),
            .I(N__52241));
    Odrv4 I__12317 (
            .O(N__52244),
            .I(N_14_3));
    LocalMux I__12316 (
            .O(N__52241),
            .I(N_14_3));
    InMux I__12315 (
            .O(N__52236),
            .I(un2_scounterdac_cry_1));
    InMux I__12314 (
            .O(N__52233),
            .I(N__52229));
    InMux I__12313 (
            .O(N__52232),
            .I(N__52226));
    LocalMux I__12312 (
            .O(N__52229),
            .I(N__52222));
    LocalMux I__12311 (
            .O(N__52226),
            .I(N__52219));
    InMux I__12310 (
            .O(N__52225),
            .I(N__52216));
    Span4Mux_h I__12309 (
            .O(N__52222),
            .I(N__52213));
    Odrv4 I__12308 (
            .O(N__52219),
            .I(sCounterDACZ0Z_3));
    LocalMux I__12307 (
            .O(N__52216),
            .I(sCounterDACZ0Z_3));
    Odrv4 I__12306 (
            .O(N__52213),
            .I(sCounterDACZ0Z_3));
    InMux I__12305 (
            .O(N__52206),
            .I(un2_scounterdac_cry_2));
    InMux I__12304 (
            .O(N__52203),
            .I(un2_scounterdac_cry_3));
    InMux I__12303 (
            .O(N__52200),
            .I(N__52194));
    InMux I__12302 (
            .O(N__52199),
            .I(N__52194));
    LocalMux I__12301 (
            .O(N__52194),
            .I(N__52190));
    InMux I__12300 (
            .O(N__52193),
            .I(N__52187));
    Span4Mux_v I__12299 (
            .O(N__52190),
            .I(N__52184));
    LocalMux I__12298 (
            .O(N__52187),
            .I(sCounterDACZ0Z_5));
    Odrv4 I__12297 (
            .O(N__52184),
            .I(sCounterDACZ0Z_5));
    InMux I__12296 (
            .O(N__52179),
            .I(un2_scounterdac_cry_4));
    InMux I__12295 (
            .O(N__52176),
            .I(N__52173));
    LocalMux I__12294 (
            .O(N__52173),
            .I(N__52170));
    Odrv4 I__12293 (
            .O(N__52170),
            .I(un2_scounterdac_cry_5_THRU_CO));
    InMux I__12292 (
            .O(N__52167),
            .I(un2_scounterdac_cry_5));
    InMux I__12291 (
            .O(N__52164),
            .I(un2_scounterdac_cry_6));
    InMux I__12290 (
            .O(N__52161),
            .I(N__52132));
    InMux I__12289 (
            .O(N__52160),
            .I(N__52132));
    InMux I__12288 (
            .O(N__52159),
            .I(N__52123));
    InMux I__12287 (
            .O(N__52158),
            .I(N__52123));
    InMux I__12286 (
            .O(N__52157),
            .I(N__52123));
    InMux I__12285 (
            .O(N__52156),
            .I(N__52123));
    InMux I__12284 (
            .O(N__52155),
            .I(N__52099));
    InMux I__12283 (
            .O(N__52154),
            .I(N__52099));
    InMux I__12282 (
            .O(N__52153),
            .I(N__52096));
    InMux I__12281 (
            .O(N__52152),
            .I(N__52084));
    InMux I__12280 (
            .O(N__52151),
            .I(N__52084));
    InMux I__12279 (
            .O(N__52150),
            .I(N__52084));
    InMux I__12278 (
            .O(N__52149),
            .I(N__52068));
    InMux I__12277 (
            .O(N__52148),
            .I(N__52068));
    InMux I__12276 (
            .O(N__52147),
            .I(N__52059));
    InMux I__12275 (
            .O(N__52146),
            .I(N__52059));
    InMux I__12274 (
            .O(N__52145),
            .I(N__52054));
    InMux I__12273 (
            .O(N__52144),
            .I(N__52054));
    InMux I__12272 (
            .O(N__52143),
            .I(N__52047));
    InMux I__12271 (
            .O(N__52142),
            .I(N__52047));
    InMux I__12270 (
            .O(N__52141),
            .I(N__52047));
    InMux I__12269 (
            .O(N__52140),
            .I(N__52042));
    InMux I__12268 (
            .O(N__52139),
            .I(N__52042));
    InMux I__12267 (
            .O(N__52138),
            .I(N__52036));
    InMux I__12266 (
            .O(N__52137),
            .I(N__52036));
    LocalMux I__12265 (
            .O(N__52132),
            .I(N__52031));
    LocalMux I__12264 (
            .O(N__52123),
            .I(N__52031));
    InMux I__12263 (
            .O(N__52122),
            .I(N__52028));
    InMux I__12262 (
            .O(N__52121),
            .I(N__52023));
    InMux I__12261 (
            .O(N__52120),
            .I(N__52023));
    InMux I__12260 (
            .O(N__52119),
            .I(N__52020));
    CascadeMux I__12259 (
            .O(N__52118),
            .I(N__52009));
    InMux I__12258 (
            .O(N__52117),
            .I(N__51986));
    InMux I__12257 (
            .O(N__52116),
            .I(N__51986));
    InMux I__12256 (
            .O(N__52115),
            .I(N__51986));
    InMux I__12255 (
            .O(N__52114),
            .I(N__51980));
    InMux I__12254 (
            .O(N__52113),
            .I(N__51975));
    InMux I__12253 (
            .O(N__52112),
            .I(N__51975));
    InMux I__12252 (
            .O(N__52111),
            .I(N__51963));
    InMux I__12251 (
            .O(N__52110),
            .I(N__51963));
    InMux I__12250 (
            .O(N__52109),
            .I(N__51963));
    InMux I__12249 (
            .O(N__52108),
            .I(N__51958));
    InMux I__12248 (
            .O(N__52107),
            .I(N__51958));
    InMux I__12247 (
            .O(N__52106),
            .I(N__51951));
    InMux I__12246 (
            .O(N__52105),
            .I(N__51951));
    InMux I__12245 (
            .O(N__52104),
            .I(N__51951));
    LocalMux I__12244 (
            .O(N__52099),
            .I(N__51948));
    LocalMux I__12243 (
            .O(N__52096),
            .I(N__51945));
    InMux I__12242 (
            .O(N__52095),
            .I(N__51934));
    InMux I__12241 (
            .O(N__52094),
            .I(N__51934));
    InMux I__12240 (
            .O(N__52093),
            .I(N__51934));
    InMux I__12239 (
            .O(N__52092),
            .I(N__51934));
    InMux I__12238 (
            .O(N__52091),
            .I(N__51934));
    LocalMux I__12237 (
            .O(N__52084),
            .I(N__51931));
    InMux I__12236 (
            .O(N__52083),
            .I(N__51924));
    InMux I__12235 (
            .O(N__52082),
            .I(N__51924));
    InMux I__12234 (
            .O(N__52081),
            .I(N__51924));
    InMux I__12233 (
            .O(N__52080),
            .I(N__51917));
    InMux I__12232 (
            .O(N__52079),
            .I(N__51917));
    InMux I__12231 (
            .O(N__52078),
            .I(N__51917));
    InMux I__12230 (
            .O(N__52077),
            .I(N__51914));
    InMux I__12229 (
            .O(N__52076),
            .I(N__51911));
    InMux I__12228 (
            .O(N__52075),
            .I(N__51897));
    InMux I__12227 (
            .O(N__52074),
            .I(N__51897));
    InMux I__12226 (
            .O(N__52073),
            .I(N__51882));
    LocalMux I__12225 (
            .O(N__52068),
            .I(N__51875));
    InMux I__12224 (
            .O(N__52067),
            .I(N__51868));
    InMux I__12223 (
            .O(N__52066),
            .I(N__51868));
    InMux I__12222 (
            .O(N__52065),
            .I(N__51868));
    InMux I__12221 (
            .O(N__52064),
            .I(N__51861));
    LocalMux I__12220 (
            .O(N__52059),
            .I(N__51858));
    LocalMux I__12219 (
            .O(N__52054),
            .I(N__51851));
    LocalMux I__12218 (
            .O(N__52047),
            .I(N__51851));
    LocalMux I__12217 (
            .O(N__52042),
            .I(N__51851));
    InMux I__12216 (
            .O(N__52041),
            .I(N__51848));
    LocalMux I__12215 (
            .O(N__52036),
            .I(N__51843));
    Span4Mux_h I__12214 (
            .O(N__52031),
            .I(N__51843));
    LocalMux I__12213 (
            .O(N__52028),
            .I(N__51836));
    LocalMux I__12212 (
            .O(N__52023),
            .I(N__51836));
    LocalMux I__12211 (
            .O(N__52020),
            .I(N__51836));
    InMux I__12210 (
            .O(N__52019),
            .I(N__51831));
    InMux I__12209 (
            .O(N__52018),
            .I(N__51831));
    InMux I__12208 (
            .O(N__52017),
            .I(N__51826));
    InMux I__12207 (
            .O(N__52016),
            .I(N__51826));
    InMux I__12206 (
            .O(N__52015),
            .I(N__51819));
    InMux I__12205 (
            .O(N__52014),
            .I(N__51819));
    InMux I__12204 (
            .O(N__52013),
            .I(N__51819));
    CascadeMux I__12203 (
            .O(N__52012),
            .I(N__51805));
    InMux I__12202 (
            .O(N__52009),
            .I(N__51794));
    InMux I__12201 (
            .O(N__52008),
            .I(N__51794));
    InMux I__12200 (
            .O(N__52007),
            .I(N__51794));
    InMux I__12199 (
            .O(N__52006),
            .I(N__51785));
    InMux I__12198 (
            .O(N__52005),
            .I(N__51785));
    InMux I__12197 (
            .O(N__52004),
            .I(N__51785));
    InMux I__12196 (
            .O(N__52003),
            .I(N__51785));
    InMux I__12195 (
            .O(N__52002),
            .I(N__51778));
    InMux I__12194 (
            .O(N__52001),
            .I(N__51778));
    InMux I__12193 (
            .O(N__52000),
            .I(N__51778));
    InMux I__12192 (
            .O(N__51999),
            .I(N__51773));
    InMux I__12191 (
            .O(N__51998),
            .I(N__51773));
    InMux I__12190 (
            .O(N__51997),
            .I(N__51763));
    InMux I__12189 (
            .O(N__51996),
            .I(N__51763));
    InMux I__12188 (
            .O(N__51995),
            .I(N__51763));
    InMux I__12187 (
            .O(N__51994),
            .I(N__51758));
    InMux I__12186 (
            .O(N__51993),
            .I(N__51758));
    LocalMux I__12185 (
            .O(N__51986),
            .I(N__51755));
    InMux I__12184 (
            .O(N__51985),
            .I(N__51752));
    InMux I__12183 (
            .O(N__51984),
            .I(N__51747));
    InMux I__12182 (
            .O(N__51983),
            .I(N__51747));
    LocalMux I__12181 (
            .O(N__51980),
            .I(N__51742));
    LocalMux I__12180 (
            .O(N__51975),
            .I(N__51742));
    InMux I__12179 (
            .O(N__51974),
            .I(N__51737));
    InMux I__12178 (
            .O(N__51973),
            .I(N__51737));
    InMux I__12177 (
            .O(N__51972),
            .I(N__51730));
    InMux I__12176 (
            .O(N__51971),
            .I(N__51730));
    InMux I__12175 (
            .O(N__51970),
            .I(N__51730));
    LocalMux I__12174 (
            .O(N__51963),
            .I(N__51727));
    LocalMux I__12173 (
            .O(N__51958),
            .I(N__51722));
    LocalMux I__12172 (
            .O(N__51951),
            .I(N__51722));
    Span4Mux_h I__12171 (
            .O(N__51948),
            .I(N__51711));
    Span4Mux_v I__12170 (
            .O(N__51945),
            .I(N__51711));
    LocalMux I__12169 (
            .O(N__51934),
            .I(N__51711));
    Span4Mux_v I__12168 (
            .O(N__51931),
            .I(N__51711));
    LocalMux I__12167 (
            .O(N__51924),
            .I(N__51711));
    LocalMux I__12166 (
            .O(N__51917),
            .I(N__51704));
    LocalMux I__12165 (
            .O(N__51914),
            .I(N__51704));
    LocalMux I__12164 (
            .O(N__51911),
            .I(N__51704));
    InMux I__12163 (
            .O(N__51910),
            .I(N__51695));
    InMux I__12162 (
            .O(N__51909),
            .I(N__51695));
    InMux I__12161 (
            .O(N__51908),
            .I(N__51695));
    InMux I__12160 (
            .O(N__51907),
            .I(N__51695));
    InMux I__12159 (
            .O(N__51906),
            .I(N__51684));
    InMux I__12158 (
            .O(N__51905),
            .I(N__51684));
    InMux I__12157 (
            .O(N__51904),
            .I(N__51684));
    InMux I__12156 (
            .O(N__51903),
            .I(N__51684));
    InMux I__12155 (
            .O(N__51902),
            .I(N__51684));
    LocalMux I__12154 (
            .O(N__51897),
            .I(N__51681));
    InMux I__12153 (
            .O(N__51896),
            .I(N__51678));
    InMux I__12152 (
            .O(N__51895),
            .I(N__51671));
    InMux I__12151 (
            .O(N__51894),
            .I(N__51671));
    InMux I__12150 (
            .O(N__51893),
            .I(N__51671));
    InMux I__12149 (
            .O(N__51892),
            .I(N__51666));
    InMux I__12148 (
            .O(N__51891),
            .I(N__51666));
    InMux I__12147 (
            .O(N__51890),
            .I(N__51663));
    InMux I__12146 (
            .O(N__51889),
            .I(N__51656));
    InMux I__12145 (
            .O(N__51888),
            .I(N__51656));
    InMux I__12144 (
            .O(N__51887),
            .I(N__51656));
    InMux I__12143 (
            .O(N__51886),
            .I(N__51651));
    InMux I__12142 (
            .O(N__51885),
            .I(N__51651));
    LocalMux I__12141 (
            .O(N__51882),
            .I(N__51648));
    InMux I__12140 (
            .O(N__51881),
            .I(N__51645));
    InMux I__12139 (
            .O(N__51880),
            .I(N__51638));
    InMux I__12138 (
            .O(N__51879),
            .I(N__51638));
    InMux I__12137 (
            .O(N__51878),
            .I(N__51638));
    Span4Mux_v I__12136 (
            .O(N__51875),
            .I(N__51633));
    LocalMux I__12135 (
            .O(N__51868),
            .I(N__51633));
    InMux I__12134 (
            .O(N__51867),
            .I(N__51624));
    InMux I__12133 (
            .O(N__51866),
            .I(N__51624));
    InMux I__12132 (
            .O(N__51865),
            .I(N__51624));
    InMux I__12131 (
            .O(N__51864),
            .I(N__51624));
    LocalMux I__12130 (
            .O(N__51861),
            .I(N__51617));
    Span4Mux_v I__12129 (
            .O(N__51858),
            .I(N__51617));
    Span4Mux_v I__12128 (
            .O(N__51851),
            .I(N__51617));
    LocalMux I__12127 (
            .O(N__51848),
            .I(N__51610));
    Span4Mux_v I__12126 (
            .O(N__51843),
            .I(N__51610));
    Span4Mux_h I__12125 (
            .O(N__51836),
            .I(N__51610));
    LocalMux I__12124 (
            .O(N__51831),
            .I(N__51603));
    LocalMux I__12123 (
            .O(N__51826),
            .I(N__51603));
    LocalMux I__12122 (
            .O(N__51819),
            .I(N__51603));
    InMux I__12121 (
            .O(N__51818),
            .I(N__51589));
    InMux I__12120 (
            .O(N__51817),
            .I(N__51589));
    InMux I__12119 (
            .O(N__51816),
            .I(N__51582));
    InMux I__12118 (
            .O(N__51815),
            .I(N__51582));
    InMux I__12117 (
            .O(N__51814),
            .I(N__51582));
    InMux I__12116 (
            .O(N__51813),
            .I(N__51577));
    InMux I__12115 (
            .O(N__51812),
            .I(N__51577));
    InMux I__12114 (
            .O(N__51811),
            .I(N__51570));
    InMux I__12113 (
            .O(N__51810),
            .I(N__51570));
    InMux I__12112 (
            .O(N__51809),
            .I(N__51570));
    InMux I__12111 (
            .O(N__51808),
            .I(N__51565));
    InMux I__12110 (
            .O(N__51805),
            .I(N__51565));
    InMux I__12109 (
            .O(N__51804),
            .I(N__51556));
    InMux I__12108 (
            .O(N__51803),
            .I(N__51556));
    InMux I__12107 (
            .O(N__51802),
            .I(N__51556));
    InMux I__12106 (
            .O(N__51801),
            .I(N__51556));
    LocalMux I__12105 (
            .O(N__51794),
            .I(N__51542));
    LocalMux I__12104 (
            .O(N__51785),
            .I(N__51542));
    LocalMux I__12103 (
            .O(N__51778),
            .I(N__51542));
    LocalMux I__12102 (
            .O(N__51773),
            .I(N__51542));
    InMux I__12101 (
            .O(N__51772),
            .I(N__51530));
    InMux I__12100 (
            .O(N__51771),
            .I(N__51530));
    InMux I__12099 (
            .O(N__51770),
            .I(N__51530));
    LocalMux I__12098 (
            .O(N__51763),
            .I(N__51521));
    LocalMux I__12097 (
            .O(N__51758),
            .I(N__51521));
    Span4Mux_v I__12096 (
            .O(N__51755),
            .I(N__51521));
    LocalMux I__12095 (
            .O(N__51752),
            .I(N__51521));
    LocalMux I__12094 (
            .O(N__51747),
            .I(N__51514));
    Span4Mux_h I__12093 (
            .O(N__51742),
            .I(N__51514));
    LocalMux I__12092 (
            .O(N__51737),
            .I(N__51514));
    LocalMux I__12091 (
            .O(N__51730),
            .I(N__51503));
    Span4Mux_v I__12090 (
            .O(N__51727),
            .I(N__51503));
    Span4Mux_v I__12089 (
            .O(N__51722),
            .I(N__51503));
    Span4Mux_h I__12088 (
            .O(N__51711),
            .I(N__51503));
    Span4Mux_h I__12087 (
            .O(N__51704),
            .I(N__51503));
    LocalMux I__12086 (
            .O(N__51695),
            .I(N__51496));
    LocalMux I__12085 (
            .O(N__51684),
            .I(N__51496));
    Span4Mux_h I__12084 (
            .O(N__51681),
            .I(N__51490));
    LocalMux I__12083 (
            .O(N__51678),
            .I(N__51481));
    LocalMux I__12082 (
            .O(N__51671),
            .I(N__51481));
    LocalMux I__12081 (
            .O(N__51666),
            .I(N__51481));
    LocalMux I__12080 (
            .O(N__51663),
            .I(N__51481));
    LocalMux I__12079 (
            .O(N__51656),
            .I(N__51472));
    LocalMux I__12078 (
            .O(N__51651),
            .I(N__51472));
    Span4Mux_h I__12077 (
            .O(N__51648),
            .I(N__51461));
    LocalMux I__12076 (
            .O(N__51645),
            .I(N__51461));
    LocalMux I__12075 (
            .O(N__51638),
            .I(N__51461));
    Span4Mux_h I__12074 (
            .O(N__51633),
            .I(N__51461));
    LocalMux I__12073 (
            .O(N__51624),
            .I(N__51461));
    Span4Mux_h I__12072 (
            .O(N__51617),
            .I(N__51454));
    Span4Mux_v I__12071 (
            .O(N__51610),
            .I(N__51454));
    Span4Mux_v I__12070 (
            .O(N__51603),
            .I(N__51454));
    InMux I__12069 (
            .O(N__51602),
            .I(N__51443));
    InMux I__12068 (
            .O(N__51601),
            .I(N__51443));
    InMux I__12067 (
            .O(N__51600),
            .I(N__51443));
    InMux I__12066 (
            .O(N__51599),
            .I(N__51443));
    InMux I__12065 (
            .O(N__51598),
            .I(N__51443));
    InMux I__12064 (
            .O(N__51597),
            .I(N__51434));
    InMux I__12063 (
            .O(N__51596),
            .I(N__51434));
    InMux I__12062 (
            .O(N__51595),
            .I(N__51434));
    InMux I__12061 (
            .O(N__51594),
            .I(N__51434));
    LocalMux I__12060 (
            .O(N__51589),
            .I(N__51421));
    LocalMux I__12059 (
            .O(N__51582),
            .I(N__51421));
    LocalMux I__12058 (
            .O(N__51577),
            .I(N__51421));
    LocalMux I__12057 (
            .O(N__51570),
            .I(N__51421));
    LocalMux I__12056 (
            .O(N__51565),
            .I(N__51421));
    LocalMux I__12055 (
            .O(N__51556),
            .I(N__51421));
    InMux I__12054 (
            .O(N__51555),
            .I(N__51412));
    InMux I__12053 (
            .O(N__51554),
            .I(N__51412));
    InMux I__12052 (
            .O(N__51553),
            .I(N__51412));
    InMux I__12051 (
            .O(N__51552),
            .I(N__51412));
    InMux I__12050 (
            .O(N__51551),
            .I(N__51409));
    Span12Mux_h I__12049 (
            .O(N__51542),
            .I(N__51406));
    InMux I__12048 (
            .O(N__51541),
            .I(N__51395));
    InMux I__12047 (
            .O(N__51540),
            .I(N__51395));
    InMux I__12046 (
            .O(N__51539),
            .I(N__51395));
    InMux I__12045 (
            .O(N__51538),
            .I(N__51395));
    InMux I__12044 (
            .O(N__51537),
            .I(N__51395));
    LocalMux I__12043 (
            .O(N__51530),
            .I(N__51386));
    Span4Mux_v I__12042 (
            .O(N__51521),
            .I(N__51386));
    Span4Mux_h I__12041 (
            .O(N__51514),
            .I(N__51386));
    Span4Mux_v I__12040 (
            .O(N__51503),
            .I(N__51386));
    InMux I__12039 (
            .O(N__51502),
            .I(N__51383));
    InMux I__12038 (
            .O(N__51501),
            .I(N__51380));
    Span12Mux_v I__12037 (
            .O(N__51496),
            .I(N__51377));
    InMux I__12036 (
            .O(N__51495),
            .I(N__51370));
    InMux I__12035 (
            .O(N__51494),
            .I(N__51370));
    InMux I__12034 (
            .O(N__51493),
            .I(N__51370));
    Span4Mux_h I__12033 (
            .O(N__51490),
            .I(N__51365));
    Span4Mux_h I__12032 (
            .O(N__51481),
            .I(N__51365));
    InMux I__12031 (
            .O(N__51480),
            .I(N__51362));
    InMux I__12030 (
            .O(N__51479),
            .I(N__51355));
    InMux I__12029 (
            .O(N__51478),
            .I(N__51355));
    InMux I__12028 (
            .O(N__51477),
            .I(N__51355));
    Span4Mux_h I__12027 (
            .O(N__51472),
            .I(N__51348));
    Span4Mux_v I__12026 (
            .O(N__51461),
            .I(N__51348));
    Span4Mux_v I__12025 (
            .O(N__51454),
            .I(N__51348));
    LocalMux I__12024 (
            .O(N__51443),
            .I(N__51339));
    LocalMux I__12023 (
            .O(N__51434),
            .I(N__51339));
    Span12Mux_h I__12022 (
            .O(N__51421),
            .I(N__51339));
    LocalMux I__12021 (
            .O(N__51412),
            .I(N__51339));
    LocalMux I__12020 (
            .O(N__51409),
            .I(N__51334));
    Span12Mux_v I__12019 (
            .O(N__51406),
            .I(N__51334));
    LocalMux I__12018 (
            .O(N__51395),
            .I(N__51329));
    Span4Mux_v I__12017 (
            .O(N__51386),
            .I(N__51329));
    LocalMux I__12016 (
            .O(N__51383),
            .I(sDAC_mem_pointerZ0Z_0));
    LocalMux I__12015 (
            .O(N__51380),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv12 I__12014 (
            .O(N__51377),
            .I(sDAC_mem_pointerZ0Z_0));
    LocalMux I__12013 (
            .O(N__51370),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv4 I__12012 (
            .O(N__51365),
            .I(sDAC_mem_pointerZ0Z_0));
    LocalMux I__12011 (
            .O(N__51362),
            .I(sDAC_mem_pointerZ0Z_0));
    LocalMux I__12010 (
            .O(N__51355),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv4 I__12009 (
            .O(N__51348),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv12 I__12008 (
            .O(N__51339),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv12 I__12007 (
            .O(N__51334),
            .I(sDAC_mem_pointerZ0Z_0));
    Odrv4 I__12006 (
            .O(N__51329),
            .I(sDAC_mem_pointerZ0Z_0));
    InMux I__12005 (
            .O(N__51306),
            .I(N__51303));
    LocalMux I__12004 (
            .O(N__51303),
            .I(sDAC_mem_15Z0Z_7));
    InMux I__12003 (
            .O(N__51300),
            .I(N__51297));
    LocalMux I__12002 (
            .O(N__51297),
            .I(N__51294));
    Span4Mux_h I__12001 (
            .O(N__51294),
            .I(N__51291));
    Odrv4 I__12000 (
            .O(N__51291),
            .I(sDAC_mem_14Z0Z_7));
    InMux I__11999 (
            .O(N__51288),
            .I(N__51285));
    LocalMux I__11998 (
            .O(N__51285),
            .I(N__51282));
    Span4Mux_h I__11997 (
            .O(N__51282),
            .I(N__51279));
    Odrv4 I__11996 (
            .O(N__51279),
            .I(sDAC_data_RNO_19Z0Z_10));
    InMux I__11995 (
            .O(N__51276),
            .I(N__51273));
    LocalMux I__11994 (
            .O(N__51273),
            .I(N__51263));
    InMux I__11993 (
            .O(N__51272),
            .I(N__51254));
    InMux I__11992 (
            .O(N__51271),
            .I(N__51249));
    InMux I__11991 (
            .O(N__51270),
            .I(N__51243));
    InMux I__11990 (
            .O(N__51269),
            .I(N__51236));
    InMux I__11989 (
            .O(N__51268),
            .I(N__51233));
    InMux I__11988 (
            .O(N__51267),
            .I(N__51229));
    InMux I__11987 (
            .O(N__51266),
            .I(N__51226));
    Span4Mux_v I__11986 (
            .O(N__51263),
            .I(N__51223));
    InMux I__11985 (
            .O(N__51262),
            .I(N__51220));
    InMux I__11984 (
            .O(N__51261),
            .I(N__51217));
    InMux I__11983 (
            .O(N__51260),
            .I(N__51213));
    InMux I__11982 (
            .O(N__51259),
            .I(N__51210));
    InMux I__11981 (
            .O(N__51258),
            .I(N__51207));
    InMux I__11980 (
            .O(N__51257),
            .I(N__51204));
    LocalMux I__11979 (
            .O(N__51254),
            .I(N__51200));
    InMux I__11978 (
            .O(N__51253),
            .I(N__51197));
    InMux I__11977 (
            .O(N__51252),
            .I(N__51194));
    LocalMux I__11976 (
            .O(N__51249),
            .I(N__51191));
    InMux I__11975 (
            .O(N__51248),
            .I(N__51188));
    InMux I__11974 (
            .O(N__51247),
            .I(N__51185));
    InMux I__11973 (
            .O(N__51246),
            .I(N__51182));
    LocalMux I__11972 (
            .O(N__51243),
            .I(N__51178));
    InMux I__11971 (
            .O(N__51242),
            .I(N__51175));
    InMux I__11970 (
            .O(N__51241),
            .I(N__51172));
    InMux I__11969 (
            .O(N__51240),
            .I(N__51169));
    InMux I__11968 (
            .O(N__51239),
            .I(N__51165));
    LocalMux I__11967 (
            .O(N__51236),
            .I(N__51159));
    LocalMux I__11966 (
            .O(N__51233),
            .I(N__51159));
    InMux I__11965 (
            .O(N__51232),
            .I(N__51152));
    LocalMux I__11964 (
            .O(N__51229),
            .I(N__51147));
    LocalMux I__11963 (
            .O(N__51226),
            .I(N__51147));
    Span4Mux_v I__11962 (
            .O(N__51223),
            .I(N__51140));
    LocalMux I__11961 (
            .O(N__51220),
            .I(N__51140));
    LocalMux I__11960 (
            .O(N__51217),
            .I(N__51140));
    InMux I__11959 (
            .O(N__51216),
            .I(N__51135));
    LocalMux I__11958 (
            .O(N__51213),
            .I(N__51127));
    LocalMux I__11957 (
            .O(N__51210),
            .I(N__51127));
    LocalMux I__11956 (
            .O(N__51207),
            .I(N__51122));
    LocalMux I__11955 (
            .O(N__51204),
            .I(N__51122));
    InMux I__11954 (
            .O(N__51203),
            .I(N__51119));
    Span4Mux_h I__11953 (
            .O(N__51200),
            .I(N__51112));
    LocalMux I__11952 (
            .O(N__51197),
            .I(N__51112));
    LocalMux I__11951 (
            .O(N__51194),
            .I(N__51112));
    Span4Mux_v I__11950 (
            .O(N__51191),
            .I(N__51105));
    LocalMux I__11949 (
            .O(N__51188),
            .I(N__51105));
    LocalMux I__11948 (
            .O(N__51185),
            .I(N__51105));
    LocalMux I__11947 (
            .O(N__51182),
            .I(N__51102));
    InMux I__11946 (
            .O(N__51181),
            .I(N__51096));
    Span4Mux_v I__11945 (
            .O(N__51178),
            .I(N__51087));
    LocalMux I__11944 (
            .O(N__51175),
            .I(N__51087));
    LocalMux I__11943 (
            .O(N__51172),
            .I(N__51087));
    LocalMux I__11942 (
            .O(N__51169),
            .I(N__51087));
    InMux I__11941 (
            .O(N__51168),
            .I(N__51084));
    LocalMux I__11940 (
            .O(N__51165),
            .I(N__51075));
    InMux I__11939 (
            .O(N__51164),
            .I(N__51072));
    Span4Mux_v I__11938 (
            .O(N__51159),
            .I(N__51069));
    InMux I__11937 (
            .O(N__51158),
            .I(N__51066));
    InMux I__11936 (
            .O(N__51157),
            .I(N__51063));
    InMux I__11935 (
            .O(N__51156),
            .I(N__51060));
    InMux I__11934 (
            .O(N__51155),
            .I(N__51057));
    LocalMux I__11933 (
            .O(N__51152),
            .I(N__51054));
    Span4Mux_v I__11932 (
            .O(N__51147),
            .I(N__51051));
    Span4Mux_v I__11931 (
            .O(N__51140),
            .I(N__51048));
    InMux I__11930 (
            .O(N__51139),
            .I(N__51045));
    InMux I__11929 (
            .O(N__51138),
            .I(N__51042));
    LocalMux I__11928 (
            .O(N__51135),
            .I(N__51037));
    InMux I__11927 (
            .O(N__51134),
            .I(N__51034));
    InMux I__11926 (
            .O(N__51133),
            .I(N__51031));
    InMux I__11925 (
            .O(N__51132),
            .I(N__51028));
    Span4Mux_v I__11924 (
            .O(N__51127),
            .I(N__51017));
    Span4Mux_h I__11923 (
            .O(N__51122),
            .I(N__51017));
    LocalMux I__11922 (
            .O(N__51119),
            .I(N__51017));
    Span4Mux_v I__11921 (
            .O(N__51112),
            .I(N__51010));
    Span4Mux_v I__11920 (
            .O(N__51105),
            .I(N__51010));
    Span4Mux_h I__11919 (
            .O(N__51102),
            .I(N__51010));
    InMux I__11918 (
            .O(N__51101),
            .I(N__51007));
    InMux I__11917 (
            .O(N__51100),
            .I(N__51004));
    InMux I__11916 (
            .O(N__51099),
            .I(N__51001));
    LocalMux I__11915 (
            .O(N__51096),
            .I(N__50994));
    Span4Mux_v I__11914 (
            .O(N__51087),
            .I(N__50994));
    LocalMux I__11913 (
            .O(N__51084),
            .I(N__50994));
    InMux I__11912 (
            .O(N__51083),
            .I(N__50991));
    InMux I__11911 (
            .O(N__51082),
            .I(N__50988));
    InMux I__11910 (
            .O(N__51081),
            .I(N__50983));
    InMux I__11909 (
            .O(N__51080),
            .I(N__50978));
    InMux I__11908 (
            .O(N__51079),
            .I(N__50975));
    InMux I__11907 (
            .O(N__51078),
            .I(N__50972));
    Span4Mux_h I__11906 (
            .O(N__51075),
            .I(N__50967));
    LocalMux I__11905 (
            .O(N__51072),
            .I(N__50967));
    Span4Mux_v I__11904 (
            .O(N__51069),
            .I(N__50956));
    LocalMux I__11903 (
            .O(N__51066),
            .I(N__50956));
    LocalMux I__11902 (
            .O(N__51063),
            .I(N__50956));
    LocalMux I__11901 (
            .O(N__51060),
            .I(N__50956));
    LocalMux I__11900 (
            .O(N__51057),
            .I(N__50956));
    Span4Mux_v I__11899 (
            .O(N__51054),
            .I(N__50953));
    Span4Mux_v I__11898 (
            .O(N__51051),
            .I(N__50944));
    Span4Mux_h I__11897 (
            .O(N__51048),
            .I(N__50944));
    LocalMux I__11896 (
            .O(N__51045),
            .I(N__50944));
    LocalMux I__11895 (
            .O(N__51042),
            .I(N__50944));
    InMux I__11894 (
            .O(N__51041),
            .I(N__50941));
    InMux I__11893 (
            .O(N__51040),
            .I(N__50938));
    Span4Mux_v I__11892 (
            .O(N__51037),
            .I(N__50929));
    LocalMux I__11891 (
            .O(N__51034),
            .I(N__50929));
    LocalMux I__11890 (
            .O(N__51031),
            .I(N__50929));
    LocalMux I__11889 (
            .O(N__51028),
            .I(N__50929));
    InMux I__11888 (
            .O(N__51027),
            .I(N__50926));
    InMux I__11887 (
            .O(N__51026),
            .I(N__50923));
    InMux I__11886 (
            .O(N__51025),
            .I(N__50920));
    InMux I__11885 (
            .O(N__51024),
            .I(N__50917));
    Span4Mux_v I__11884 (
            .O(N__51017),
            .I(N__50914));
    Span4Mux_v I__11883 (
            .O(N__51010),
            .I(N__50905));
    LocalMux I__11882 (
            .O(N__51007),
            .I(N__50905));
    LocalMux I__11881 (
            .O(N__51004),
            .I(N__50905));
    LocalMux I__11880 (
            .O(N__51001),
            .I(N__50905));
    Span4Mux_v I__11879 (
            .O(N__50994),
            .I(N__50898));
    LocalMux I__11878 (
            .O(N__50991),
            .I(N__50898));
    LocalMux I__11877 (
            .O(N__50988),
            .I(N__50898));
    InMux I__11876 (
            .O(N__50987),
            .I(N__50895));
    InMux I__11875 (
            .O(N__50986),
            .I(N__50892));
    LocalMux I__11874 (
            .O(N__50983),
            .I(N__50889));
    InMux I__11873 (
            .O(N__50982),
            .I(N__50886));
    InMux I__11872 (
            .O(N__50981),
            .I(N__50883));
    LocalMux I__11871 (
            .O(N__50978),
            .I(N__50874));
    LocalMux I__11870 (
            .O(N__50975),
            .I(N__50874));
    LocalMux I__11869 (
            .O(N__50972),
            .I(N__50874));
    Span4Mux_v I__11868 (
            .O(N__50967),
            .I(N__50867));
    Span4Mux_v I__11867 (
            .O(N__50956),
            .I(N__50867));
    Span4Mux_h I__11866 (
            .O(N__50953),
            .I(N__50860));
    Span4Mux_v I__11865 (
            .O(N__50944),
            .I(N__50860));
    LocalMux I__11864 (
            .O(N__50941),
            .I(N__50860));
    LocalMux I__11863 (
            .O(N__50938),
            .I(N__50857));
    Span4Mux_v I__11862 (
            .O(N__50929),
            .I(N__50846));
    LocalMux I__11861 (
            .O(N__50926),
            .I(N__50846));
    LocalMux I__11860 (
            .O(N__50923),
            .I(N__50846));
    LocalMux I__11859 (
            .O(N__50920),
            .I(N__50846));
    LocalMux I__11858 (
            .O(N__50917),
            .I(N__50846));
    Span4Mux_h I__11857 (
            .O(N__50914),
            .I(N__50835));
    Span4Mux_v I__11856 (
            .O(N__50905),
            .I(N__50835));
    Span4Mux_h I__11855 (
            .O(N__50898),
            .I(N__50835));
    LocalMux I__11854 (
            .O(N__50895),
            .I(N__50835));
    LocalMux I__11853 (
            .O(N__50892),
            .I(N__50835));
    Sp12to4 I__11852 (
            .O(N__50889),
            .I(N__50828));
    LocalMux I__11851 (
            .O(N__50886),
            .I(N__50828));
    LocalMux I__11850 (
            .O(N__50883),
            .I(N__50828));
    InMux I__11849 (
            .O(N__50882),
            .I(N__50825));
    InMux I__11848 (
            .O(N__50881),
            .I(N__50822));
    Span4Mux_v I__11847 (
            .O(N__50874),
            .I(N__50819));
    InMux I__11846 (
            .O(N__50873),
            .I(N__50814));
    InMux I__11845 (
            .O(N__50872),
            .I(N__50814));
    Span4Mux_h I__11844 (
            .O(N__50867),
            .I(N__50807));
    Span4Mux_v I__11843 (
            .O(N__50860),
            .I(N__50807));
    Span4Mux_v I__11842 (
            .O(N__50857),
            .I(N__50807));
    Span4Mux_v I__11841 (
            .O(N__50846),
            .I(N__50804));
    Span4Mux_h I__11840 (
            .O(N__50835),
            .I(N__50801));
    Span12Mux_v I__11839 (
            .O(N__50828),
            .I(N__50796));
    LocalMux I__11838 (
            .O(N__50825),
            .I(N__50796));
    LocalMux I__11837 (
            .O(N__50822),
            .I(N__50789));
    Sp12to4 I__11836 (
            .O(N__50819),
            .I(N__50789));
    LocalMux I__11835 (
            .O(N__50814),
            .I(N__50789));
    Odrv4 I__11834 (
            .O(N__50807),
            .I(spi_data_mosi_0));
    Odrv4 I__11833 (
            .O(N__50804),
            .I(spi_data_mosi_0));
    Odrv4 I__11832 (
            .O(N__50801),
            .I(spi_data_mosi_0));
    Odrv12 I__11831 (
            .O(N__50796),
            .I(spi_data_mosi_0));
    Odrv12 I__11830 (
            .O(N__50789),
            .I(spi_data_mosi_0));
    InMux I__11829 (
            .O(N__50778),
            .I(N__50775));
    LocalMux I__11828 (
            .O(N__50775),
            .I(sDAC_mem_13Z0Z_0));
    InMux I__11827 (
            .O(N__50772),
            .I(N__50766));
    InMux I__11826 (
            .O(N__50771),
            .I(N__50763));
    InMux I__11825 (
            .O(N__50770),
            .I(N__50758));
    InMux I__11824 (
            .O(N__50769),
            .I(N__50755));
    LocalMux I__11823 (
            .O(N__50766),
            .I(N__50750));
    LocalMux I__11822 (
            .O(N__50763),
            .I(N__50747));
    InMux I__11821 (
            .O(N__50762),
            .I(N__50744));
    InMux I__11820 (
            .O(N__50761),
            .I(N__50741));
    LocalMux I__11819 (
            .O(N__50758),
            .I(N__50735));
    LocalMux I__11818 (
            .O(N__50755),
            .I(N__50735));
    InMux I__11817 (
            .O(N__50754),
            .I(N__50729));
    InMux I__11816 (
            .O(N__50753),
            .I(N__50726));
    Span4Mux_v I__11815 (
            .O(N__50750),
            .I(N__50714));
    Span4Mux_v I__11814 (
            .O(N__50747),
            .I(N__50714));
    LocalMux I__11813 (
            .O(N__50744),
            .I(N__50714));
    LocalMux I__11812 (
            .O(N__50741),
            .I(N__50714));
    InMux I__11811 (
            .O(N__50740),
            .I(N__50711));
    Span4Mux_v I__11810 (
            .O(N__50735),
            .I(N__50704));
    InMux I__11809 (
            .O(N__50734),
            .I(N__50701));
    InMux I__11808 (
            .O(N__50733),
            .I(N__50698));
    InMux I__11807 (
            .O(N__50732),
            .I(N__50695));
    LocalMux I__11806 (
            .O(N__50729),
            .I(N__50688));
    LocalMux I__11805 (
            .O(N__50726),
            .I(N__50682));
    InMux I__11804 (
            .O(N__50725),
            .I(N__50679));
    InMux I__11803 (
            .O(N__50724),
            .I(N__50669));
    InMux I__11802 (
            .O(N__50723),
            .I(N__50666));
    Span4Mux_v I__11801 (
            .O(N__50714),
            .I(N__50659));
    LocalMux I__11800 (
            .O(N__50711),
            .I(N__50659));
    InMux I__11799 (
            .O(N__50710),
            .I(N__50656));
    InMux I__11798 (
            .O(N__50709),
            .I(N__50653));
    InMux I__11797 (
            .O(N__50708),
            .I(N__50650));
    InMux I__11796 (
            .O(N__50707),
            .I(N__50647));
    Span4Mux_h I__11795 (
            .O(N__50704),
            .I(N__50638));
    LocalMux I__11794 (
            .O(N__50701),
            .I(N__50638));
    LocalMux I__11793 (
            .O(N__50698),
            .I(N__50638));
    LocalMux I__11792 (
            .O(N__50695),
            .I(N__50638));
    InMux I__11791 (
            .O(N__50694),
            .I(N__50635));
    InMux I__11790 (
            .O(N__50693),
            .I(N__50632));
    InMux I__11789 (
            .O(N__50692),
            .I(N__50629));
    InMux I__11788 (
            .O(N__50691),
            .I(N__50626));
    Span4Mux_v I__11787 (
            .O(N__50688),
            .I(N__50622));
    InMux I__11786 (
            .O(N__50687),
            .I(N__50619));
    InMux I__11785 (
            .O(N__50686),
            .I(N__50616));
    InMux I__11784 (
            .O(N__50685),
            .I(N__50613));
    Span4Mux_v I__11783 (
            .O(N__50682),
            .I(N__50608));
    LocalMux I__11782 (
            .O(N__50679),
            .I(N__50608));
    InMux I__11781 (
            .O(N__50678),
            .I(N__50605));
    InMux I__11780 (
            .O(N__50677),
            .I(N__50602));
    InMux I__11779 (
            .O(N__50676),
            .I(N__50596));
    InMux I__11778 (
            .O(N__50675),
            .I(N__50593));
    InMux I__11777 (
            .O(N__50674),
            .I(N__50589));
    InMux I__11776 (
            .O(N__50673),
            .I(N__50586));
    InMux I__11775 (
            .O(N__50672),
            .I(N__50577));
    LocalMux I__11774 (
            .O(N__50669),
            .I(N__50567));
    LocalMux I__11773 (
            .O(N__50666),
            .I(N__50567));
    InMux I__11772 (
            .O(N__50665),
            .I(N__50564));
    InMux I__11771 (
            .O(N__50664),
            .I(N__50561));
    Span4Mux_v I__11770 (
            .O(N__50659),
            .I(N__50549));
    LocalMux I__11769 (
            .O(N__50656),
            .I(N__50549));
    LocalMux I__11768 (
            .O(N__50653),
            .I(N__50549));
    LocalMux I__11767 (
            .O(N__50650),
            .I(N__50549));
    LocalMux I__11766 (
            .O(N__50647),
            .I(N__50549));
    Span4Mux_v I__11765 (
            .O(N__50638),
            .I(N__50542));
    LocalMux I__11764 (
            .O(N__50635),
            .I(N__50542));
    LocalMux I__11763 (
            .O(N__50632),
            .I(N__50542));
    LocalMux I__11762 (
            .O(N__50629),
            .I(N__50537));
    LocalMux I__11761 (
            .O(N__50626),
            .I(N__50537));
    InMux I__11760 (
            .O(N__50625),
            .I(N__50534));
    Span4Mux_v I__11759 (
            .O(N__50622),
            .I(N__50525));
    LocalMux I__11758 (
            .O(N__50619),
            .I(N__50525));
    LocalMux I__11757 (
            .O(N__50616),
            .I(N__50525));
    LocalMux I__11756 (
            .O(N__50613),
            .I(N__50525));
    Span4Mux_v I__11755 (
            .O(N__50608),
            .I(N__50518));
    LocalMux I__11754 (
            .O(N__50605),
            .I(N__50518));
    LocalMux I__11753 (
            .O(N__50602),
            .I(N__50518));
    InMux I__11752 (
            .O(N__50601),
            .I(N__50515));
    InMux I__11751 (
            .O(N__50600),
            .I(N__50512));
    InMux I__11750 (
            .O(N__50599),
            .I(N__50509));
    LocalMux I__11749 (
            .O(N__50596),
            .I(N__50504));
    LocalMux I__11748 (
            .O(N__50593),
            .I(N__50504));
    InMux I__11747 (
            .O(N__50592),
            .I(N__50501));
    LocalMux I__11746 (
            .O(N__50589),
            .I(N__50497));
    LocalMux I__11745 (
            .O(N__50586),
            .I(N__50494));
    InMux I__11744 (
            .O(N__50585),
            .I(N__50491));
    InMux I__11743 (
            .O(N__50584),
            .I(N__50488));
    InMux I__11742 (
            .O(N__50583),
            .I(N__50485));
    InMux I__11741 (
            .O(N__50582),
            .I(N__50482));
    InMux I__11740 (
            .O(N__50581),
            .I(N__50479));
    InMux I__11739 (
            .O(N__50580),
            .I(N__50476));
    LocalMux I__11738 (
            .O(N__50577),
            .I(N__50473));
    InMux I__11737 (
            .O(N__50576),
            .I(N__50470));
    InMux I__11736 (
            .O(N__50575),
            .I(N__50467));
    InMux I__11735 (
            .O(N__50574),
            .I(N__50464));
    InMux I__11734 (
            .O(N__50573),
            .I(N__50461));
    InMux I__11733 (
            .O(N__50572),
            .I(N__50458));
    Span4Mux_v I__11732 (
            .O(N__50567),
            .I(N__50451));
    LocalMux I__11731 (
            .O(N__50564),
            .I(N__50448));
    LocalMux I__11730 (
            .O(N__50561),
            .I(N__50445));
    InMux I__11729 (
            .O(N__50560),
            .I(N__50442));
    Span4Mux_v I__11728 (
            .O(N__50549),
            .I(N__50439));
    Span4Mux_v I__11727 (
            .O(N__50542),
            .I(N__50432));
    Span4Mux_h I__11726 (
            .O(N__50537),
            .I(N__50432));
    LocalMux I__11725 (
            .O(N__50534),
            .I(N__50432));
    Span4Mux_v I__11724 (
            .O(N__50525),
            .I(N__50423));
    Span4Mux_h I__11723 (
            .O(N__50518),
            .I(N__50423));
    LocalMux I__11722 (
            .O(N__50515),
            .I(N__50423));
    LocalMux I__11721 (
            .O(N__50512),
            .I(N__50423));
    LocalMux I__11720 (
            .O(N__50509),
            .I(N__50415));
    Sp12to4 I__11719 (
            .O(N__50504),
            .I(N__50415));
    LocalMux I__11718 (
            .O(N__50501),
            .I(N__50415));
    InMux I__11717 (
            .O(N__50500),
            .I(N__50412));
    Span12Mux_s11_v I__11716 (
            .O(N__50497),
            .I(N__50393));
    Sp12to4 I__11715 (
            .O(N__50494),
            .I(N__50393));
    LocalMux I__11714 (
            .O(N__50491),
            .I(N__50393));
    LocalMux I__11713 (
            .O(N__50488),
            .I(N__50393));
    LocalMux I__11712 (
            .O(N__50485),
            .I(N__50393));
    LocalMux I__11711 (
            .O(N__50482),
            .I(N__50393));
    LocalMux I__11710 (
            .O(N__50479),
            .I(N__50393));
    LocalMux I__11709 (
            .O(N__50476),
            .I(N__50393));
    Sp12to4 I__11708 (
            .O(N__50473),
            .I(N__50393));
    LocalMux I__11707 (
            .O(N__50470),
            .I(N__50386));
    LocalMux I__11706 (
            .O(N__50467),
            .I(N__50386));
    LocalMux I__11705 (
            .O(N__50464),
            .I(N__50386));
    LocalMux I__11704 (
            .O(N__50461),
            .I(N__50381));
    LocalMux I__11703 (
            .O(N__50458),
            .I(N__50381));
    InMux I__11702 (
            .O(N__50457),
            .I(N__50378));
    InMux I__11701 (
            .O(N__50456),
            .I(N__50375));
    InMux I__11700 (
            .O(N__50455),
            .I(N__50372));
    InMux I__11699 (
            .O(N__50454),
            .I(N__50369));
    Span4Mux_h I__11698 (
            .O(N__50451),
            .I(N__50360));
    Span4Mux_h I__11697 (
            .O(N__50448),
            .I(N__50360));
    Span4Mux_v I__11696 (
            .O(N__50445),
            .I(N__50360));
    LocalMux I__11695 (
            .O(N__50442),
            .I(N__50360));
    Span4Mux_h I__11694 (
            .O(N__50439),
            .I(N__50355));
    Span4Mux_v I__11693 (
            .O(N__50432),
            .I(N__50355));
    Span4Mux_h I__11692 (
            .O(N__50423),
            .I(N__50352));
    InMux I__11691 (
            .O(N__50422),
            .I(N__50349));
    Span12Mux_v I__11690 (
            .O(N__50415),
            .I(N__50342));
    LocalMux I__11689 (
            .O(N__50412),
            .I(N__50342));
    Span12Mux_v I__11688 (
            .O(N__50393),
            .I(N__50342));
    Span12Mux_h I__11687 (
            .O(N__50386),
            .I(N__50327));
    Span12Mux_v I__11686 (
            .O(N__50381),
            .I(N__50327));
    LocalMux I__11685 (
            .O(N__50378),
            .I(N__50327));
    LocalMux I__11684 (
            .O(N__50375),
            .I(N__50327));
    LocalMux I__11683 (
            .O(N__50372),
            .I(N__50327));
    LocalMux I__11682 (
            .O(N__50369),
            .I(N__50327));
    Sp12to4 I__11681 (
            .O(N__50360),
            .I(N__50327));
    Odrv4 I__11680 (
            .O(N__50355),
            .I(spi_data_mosi_1));
    Odrv4 I__11679 (
            .O(N__50352),
            .I(spi_data_mosi_1));
    LocalMux I__11678 (
            .O(N__50349),
            .I(spi_data_mosi_1));
    Odrv12 I__11677 (
            .O(N__50342),
            .I(spi_data_mosi_1));
    Odrv12 I__11676 (
            .O(N__50327),
            .I(spi_data_mosi_1));
    InMux I__11675 (
            .O(N__50316),
            .I(N__50313));
    LocalMux I__11674 (
            .O(N__50313),
            .I(sDAC_mem_13Z0Z_1));
    InMux I__11673 (
            .O(N__50310),
            .I(N__50302));
    InMux I__11672 (
            .O(N__50309),
            .I(N__50296));
    InMux I__11671 (
            .O(N__50308),
            .I(N__50293));
    InMux I__11670 (
            .O(N__50307),
            .I(N__50288));
    InMux I__11669 (
            .O(N__50306),
            .I(N__50278));
    InMux I__11668 (
            .O(N__50305),
            .I(N__50275));
    LocalMux I__11667 (
            .O(N__50302),
            .I(N__50271));
    InMux I__11666 (
            .O(N__50301),
            .I(N__50268));
    InMux I__11665 (
            .O(N__50300),
            .I(N__50265));
    InMux I__11664 (
            .O(N__50299),
            .I(N__50258));
    LocalMux I__11663 (
            .O(N__50296),
            .I(N__50250));
    LocalMux I__11662 (
            .O(N__50293),
            .I(N__50250));
    InMux I__11661 (
            .O(N__50292),
            .I(N__50247));
    InMux I__11660 (
            .O(N__50291),
            .I(N__50244));
    LocalMux I__11659 (
            .O(N__50288),
            .I(N__50237));
    InMux I__11658 (
            .O(N__50287),
            .I(N__50234));
    InMux I__11657 (
            .O(N__50286),
            .I(N__50231));
    InMux I__11656 (
            .O(N__50285),
            .I(N__50227));
    InMux I__11655 (
            .O(N__50284),
            .I(N__50224));
    InMux I__11654 (
            .O(N__50283),
            .I(N__50221));
    InMux I__11653 (
            .O(N__50282),
            .I(N__50218));
    InMux I__11652 (
            .O(N__50281),
            .I(N__50215));
    LocalMux I__11651 (
            .O(N__50278),
            .I(N__50210));
    LocalMux I__11650 (
            .O(N__50275),
            .I(N__50210));
    InMux I__11649 (
            .O(N__50274),
            .I(N__50207));
    Span4Mux_v I__11648 (
            .O(N__50271),
            .I(N__50200));
    LocalMux I__11647 (
            .O(N__50268),
            .I(N__50200));
    LocalMux I__11646 (
            .O(N__50265),
            .I(N__50200));
    InMux I__11645 (
            .O(N__50264),
            .I(N__50197));
    InMux I__11644 (
            .O(N__50263),
            .I(N__50194));
    InMux I__11643 (
            .O(N__50262),
            .I(N__50191));
    InMux I__11642 (
            .O(N__50261),
            .I(N__50188));
    LocalMux I__11641 (
            .O(N__50258),
            .I(N__50184));
    InMux I__11640 (
            .O(N__50257),
            .I(N__50181));
    InMux I__11639 (
            .O(N__50256),
            .I(N__50175));
    InMux I__11638 (
            .O(N__50255),
            .I(N__50171));
    Span4Mux_v I__11637 (
            .O(N__50250),
            .I(N__50164));
    LocalMux I__11636 (
            .O(N__50247),
            .I(N__50164));
    LocalMux I__11635 (
            .O(N__50244),
            .I(N__50164));
    InMux I__11634 (
            .O(N__50243),
            .I(N__50161));
    InMux I__11633 (
            .O(N__50242),
            .I(N__50158));
    InMux I__11632 (
            .O(N__50241),
            .I(N__50155));
    InMux I__11631 (
            .O(N__50240),
            .I(N__50152));
    Span4Mux_v I__11630 (
            .O(N__50237),
            .I(N__50144));
    LocalMux I__11629 (
            .O(N__50234),
            .I(N__50144));
    LocalMux I__11628 (
            .O(N__50231),
            .I(N__50144));
    InMux I__11627 (
            .O(N__50230),
            .I(N__50141));
    LocalMux I__11626 (
            .O(N__50227),
            .I(N__50132));
    LocalMux I__11625 (
            .O(N__50224),
            .I(N__50132));
    LocalMux I__11624 (
            .O(N__50221),
            .I(N__50132));
    LocalMux I__11623 (
            .O(N__50218),
            .I(N__50132));
    LocalMux I__11622 (
            .O(N__50215),
            .I(N__50129));
    Span4Mux_v I__11621 (
            .O(N__50210),
            .I(N__50124));
    LocalMux I__11620 (
            .O(N__50207),
            .I(N__50124));
    Span4Mux_v I__11619 (
            .O(N__50200),
            .I(N__50112));
    LocalMux I__11618 (
            .O(N__50197),
            .I(N__50112));
    LocalMux I__11617 (
            .O(N__50194),
            .I(N__50112));
    LocalMux I__11616 (
            .O(N__50191),
            .I(N__50112));
    LocalMux I__11615 (
            .O(N__50188),
            .I(N__50112));
    InMux I__11614 (
            .O(N__50187),
            .I(N__50109));
    Span4Mux_h I__11613 (
            .O(N__50184),
            .I(N__50100));
    LocalMux I__11612 (
            .O(N__50181),
            .I(N__50100));
    InMux I__11611 (
            .O(N__50180),
            .I(N__50097));
    InMux I__11610 (
            .O(N__50179),
            .I(N__50094));
    InMux I__11609 (
            .O(N__50178),
            .I(N__50087));
    LocalMux I__11608 (
            .O(N__50175),
            .I(N__50084));
    InMux I__11607 (
            .O(N__50174),
            .I(N__50081));
    LocalMux I__11606 (
            .O(N__50171),
            .I(N__50074));
    Span4Mux_h I__11605 (
            .O(N__50164),
            .I(N__50063));
    LocalMux I__11604 (
            .O(N__50161),
            .I(N__50063));
    LocalMux I__11603 (
            .O(N__50158),
            .I(N__50063));
    LocalMux I__11602 (
            .O(N__50155),
            .I(N__50063));
    LocalMux I__11601 (
            .O(N__50152),
            .I(N__50063));
    InMux I__11600 (
            .O(N__50151),
            .I(N__50060));
    Span4Mux_v I__11599 (
            .O(N__50144),
            .I(N__50055));
    LocalMux I__11598 (
            .O(N__50141),
            .I(N__50055));
    Span4Mux_v I__11597 (
            .O(N__50132),
            .I(N__50052));
    Span4Mux_h I__11596 (
            .O(N__50129),
            .I(N__50047));
    Span4Mux_v I__11595 (
            .O(N__50124),
            .I(N__50047));
    InMux I__11594 (
            .O(N__50123),
            .I(N__50044));
    Span4Mux_v I__11593 (
            .O(N__50112),
            .I(N__50039));
    LocalMux I__11592 (
            .O(N__50109),
            .I(N__50039));
    InMux I__11591 (
            .O(N__50108),
            .I(N__50036));
    InMux I__11590 (
            .O(N__50107),
            .I(N__50033));
    InMux I__11589 (
            .O(N__50106),
            .I(N__50030));
    InMux I__11588 (
            .O(N__50105),
            .I(N__50027));
    Span4Mux_v I__11587 (
            .O(N__50100),
            .I(N__50016));
    LocalMux I__11586 (
            .O(N__50097),
            .I(N__50016));
    LocalMux I__11585 (
            .O(N__50094),
            .I(N__50016));
    InMux I__11584 (
            .O(N__50093),
            .I(N__50013));
    InMux I__11583 (
            .O(N__50092),
            .I(N__50010));
    InMux I__11582 (
            .O(N__50091),
            .I(N__50007));
    InMux I__11581 (
            .O(N__50090),
            .I(N__50001));
    LocalMux I__11580 (
            .O(N__50087),
            .I(N__49998));
    Span4Mux_v I__11579 (
            .O(N__50084),
            .I(N__49993));
    LocalMux I__11578 (
            .O(N__50081),
            .I(N__49993));
    InMux I__11577 (
            .O(N__50080),
            .I(N__49990));
    InMux I__11576 (
            .O(N__50079),
            .I(N__49987));
    InMux I__11575 (
            .O(N__50078),
            .I(N__49984));
    InMux I__11574 (
            .O(N__50077),
            .I(N__49981));
    Span4Mux_h I__11573 (
            .O(N__50074),
            .I(N__49974));
    Span4Mux_v I__11572 (
            .O(N__50063),
            .I(N__49974));
    LocalMux I__11571 (
            .O(N__50060),
            .I(N__49974));
    Span4Mux_v I__11570 (
            .O(N__50055),
            .I(N__49971));
    Span4Mux_h I__11569 (
            .O(N__50052),
            .I(N__49964));
    Span4Mux_v I__11568 (
            .O(N__50047),
            .I(N__49964));
    LocalMux I__11567 (
            .O(N__50044),
            .I(N__49964));
    Span4Mux_v I__11566 (
            .O(N__50039),
            .I(N__49955));
    LocalMux I__11565 (
            .O(N__50036),
            .I(N__49955));
    LocalMux I__11564 (
            .O(N__50033),
            .I(N__49955));
    LocalMux I__11563 (
            .O(N__50030),
            .I(N__49955));
    LocalMux I__11562 (
            .O(N__50027),
            .I(N__49952));
    InMux I__11561 (
            .O(N__50026),
            .I(N__49949));
    InMux I__11560 (
            .O(N__50025),
            .I(N__49946));
    InMux I__11559 (
            .O(N__50024),
            .I(N__49943));
    InMux I__11558 (
            .O(N__50023),
            .I(N__49940));
    Span4Mux_v I__11557 (
            .O(N__50016),
            .I(N__49931));
    LocalMux I__11556 (
            .O(N__50013),
            .I(N__49931));
    LocalMux I__11555 (
            .O(N__50010),
            .I(N__49931));
    LocalMux I__11554 (
            .O(N__50007),
            .I(N__49931));
    InMux I__11553 (
            .O(N__50006),
            .I(N__49928));
    InMux I__11552 (
            .O(N__50005),
            .I(N__49925));
    InMux I__11551 (
            .O(N__50004),
            .I(N__49922));
    LocalMux I__11550 (
            .O(N__50001),
            .I(N__49907));
    Span12Mux_h I__11549 (
            .O(N__49998),
            .I(N__49907));
    Sp12to4 I__11548 (
            .O(N__49993),
            .I(N__49907));
    LocalMux I__11547 (
            .O(N__49990),
            .I(N__49907));
    LocalMux I__11546 (
            .O(N__49987),
            .I(N__49907));
    LocalMux I__11545 (
            .O(N__49984),
            .I(N__49907));
    LocalMux I__11544 (
            .O(N__49981),
            .I(N__49907));
    Span4Mux_h I__11543 (
            .O(N__49974),
            .I(N__49903));
    Span4Mux_h I__11542 (
            .O(N__49971),
            .I(N__49896));
    Span4Mux_v I__11541 (
            .O(N__49964),
            .I(N__49896));
    Span4Mux_v I__11540 (
            .O(N__49955),
            .I(N__49896));
    Span12Mux_h I__11539 (
            .O(N__49952),
            .I(N__49885));
    LocalMux I__11538 (
            .O(N__49949),
            .I(N__49885));
    LocalMux I__11537 (
            .O(N__49946),
            .I(N__49885));
    LocalMux I__11536 (
            .O(N__49943),
            .I(N__49885));
    LocalMux I__11535 (
            .O(N__49940),
            .I(N__49885));
    Span4Mux_v I__11534 (
            .O(N__49931),
            .I(N__49878));
    LocalMux I__11533 (
            .O(N__49928),
            .I(N__49878));
    LocalMux I__11532 (
            .O(N__49925),
            .I(N__49878));
    LocalMux I__11531 (
            .O(N__49922),
            .I(N__49873));
    Span12Mux_v I__11530 (
            .O(N__49907),
            .I(N__49873));
    InMux I__11529 (
            .O(N__49906),
            .I(N__49870));
    Odrv4 I__11528 (
            .O(N__49903),
            .I(spi_data_mosi_2));
    Odrv4 I__11527 (
            .O(N__49896),
            .I(spi_data_mosi_2));
    Odrv12 I__11526 (
            .O(N__49885),
            .I(spi_data_mosi_2));
    Odrv4 I__11525 (
            .O(N__49878),
            .I(spi_data_mosi_2));
    Odrv12 I__11524 (
            .O(N__49873),
            .I(spi_data_mosi_2));
    LocalMux I__11523 (
            .O(N__49870),
            .I(spi_data_mosi_2));
    InMux I__11522 (
            .O(N__49857),
            .I(N__49854));
    LocalMux I__11521 (
            .O(N__49854),
            .I(N__49851));
    Span12Mux_v I__11520 (
            .O(N__49851),
            .I(N__49848));
    Odrv12 I__11519 (
            .O(N__49848),
            .I(sDAC_mem_13Z0Z_2));
    InMux I__11518 (
            .O(N__49845),
            .I(N__49838));
    InMux I__11517 (
            .O(N__49844),
            .I(N__49830));
    InMux I__11516 (
            .O(N__49843),
            .I(N__49827));
    InMux I__11515 (
            .O(N__49842),
            .I(N__49815));
    InMux I__11514 (
            .O(N__49841),
            .I(N__49812));
    LocalMux I__11513 (
            .O(N__49838),
            .I(N__49808));
    InMux I__11512 (
            .O(N__49837),
            .I(N__49805));
    InMux I__11511 (
            .O(N__49836),
            .I(N__49802));
    InMux I__11510 (
            .O(N__49835),
            .I(N__49799));
    InMux I__11509 (
            .O(N__49834),
            .I(N__49791));
    InMux I__11508 (
            .O(N__49833),
            .I(N__49787));
    LocalMux I__11507 (
            .O(N__49830),
            .I(N__49779));
    LocalMux I__11506 (
            .O(N__49827),
            .I(N__49779));
    InMux I__11505 (
            .O(N__49826),
            .I(N__49776));
    InMux I__11504 (
            .O(N__49825),
            .I(N__49773));
    InMux I__11503 (
            .O(N__49824),
            .I(N__49770));
    InMux I__11502 (
            .O(N__49823),
            .I(N__49762));
    InMux I__11501 (
            .O(N__49822),
            .I(N__49759));
    InMux I__11500 (
            .O(N__49821),
            .I(N__49756));
    InMux I__11499 (
            .O(N__49820),
            .I(N__49753));
    InMux I__11498 (
            .O(N__49819),
            .I(N__49750));
    InMux I__11497 (
            .O(N__49818),
            .I(N__49747));
    LocalMux I__11496 (
            .O(N__49815),
            .I(N__49744));
    LocalMux I__11495 (
            .O(N__49812),
            .I(N__49741));
    InMux I__11494 (
            .O(N__49811),
            .I(N__49738));
    Span4Mux_h I__11493 (
            .O(N__49808),
            .I(N__49729));
    LocalMux I__11492 (
            .O(N__49805),
            .I(N__49729));
    LocalMux I__11491 (
            .O(N__49802),
            .I(N__49726));
    LocalMux I__11490 (
            .O(N__49799),
            .I(N__49723));
    InMux I__11489 (
            .O(N__49798),
            .I(N__49720));
    InMux I__11488 (
            .O(N__49797),
            .I(N__49717));
    InMux I__11487 (
            .O(N__49796),
            .I(N__49714));
    InMux I__11486 (
            .O(N__49795),
            .I(N__49711));
    InMux I__11485 (
            .O(N__49794),
            .I(N__49708));
    LocalMux I__11484 (
            .O(N__49791),
            .I(N__49705));
    InMux I__11483 (
            .O(N__49790),
            .I(N__49699));
    LocalMux I__11482 (
            .O(N__49787),
            .I(N__49696));
    InMux I__11481 (
            .O(N__49786),
            .I(N__49693));
    InMux I__11480 (
            .O(N__49785),
            .I(N__49690));
    InMux I__11479 (
            .O(N__49784),
            .I(N__49686));
    Span4Mux_v I__11478 (
            .O(N__49779),
            .I(N__49677));
    LocalMux I__11477 (
            .O(N__49776),
            .I(N__49677));
    LocalMux I__11476 (
            .O(N__49773),
            .I(N__49677));
    LocalMux I__11475 (
            .O(N__49770),
            .I(N__49677));
    InMux I__11474 (
            .O(N__49769),
            .I(N__49674));
    InMux I__11473 (
            .O(N__49768),
            .I(N__49671));
    InMux I__11472 (
            .O(N__49767),
            .I(N__49668));
    InMux I__11471 (
            .O(N__49766),
            .I(N__49665));
    InMux I__11470 (
            .O(N__49765),
            .I(N__49662));
    LocalMux I__11469 (
            .O(N__49762),
            .I(N__49652));
    LocalMux I__11468 (
            .O(N__49759),
            .I(N__49652));
    LocalMux I__11467 (
            .O(N__49756),
            .I(N__49652));
    LocalMux I__11466 (
            .O(N__49753),
            .I(N__49652));
    LocalMux I__11465 (
            .O(N__49750),
            .I(N__49646));
    LocalMux I__11464 (
            .O(N__49747),
            .I(N__49646));
    Span4Mux_v I__11463 (
            .O(N__49744),
            .I(N__49639));
    Span4Mux_v I__11462 (
            .O(N__49741),
            .I(N__49639));
    LocalMux I__11461 (
            .O(N__49738),
            .I(N__49639));
    InMux I__11460 (
            .O(N__49737),
            .I(N__49636));
    InMux I__11459 (
            .O(N__49736),
            .I(N__49633));
    InMux I__11458 (
            .O(N__49735),
            .I(N__49630));
    InMux I__11457 (
            .O(N__49734),
            .I(N__49627));
    Span4Mux_v I__11456 (
            .O(N__49729),
            .I(N__49611));
    Span4Mux_h I__11455 (
            .O(N__49726),
            .I(N__49611));
    Span4Mux_v I__11454 (
            .O(N__49723),
            .I(N__49611));
    LocalMux I__11453 (
            .O(N__49720),
            .I(N__49611));
    LocalMux I__11452 (
            .O(N__49717),
            .I(N__49611));
    LocalMux I__11451 (
            .O(N__49714),
            .I(N__49611));
    LocalMux I__11450 (
            .O(N__49711),
            .I(N__49611));
    LocalMux I__11449 (
            .O(N__49708),
            .I(N__49605));
    Span4Mux_h I__11448 (
            .O(N__49705),
            .I(N__49602));
    InMux I__11447 (
            .O(N__49704),
            .I(N__49599));
    InMux I__11446 (
            .O(N__49703),
            .I(N__49596));
    InMux I__11445 (
            .O(N__49702),
            .I(N__49593));
    LocalMux I__11444 (
            .O(N__49699),
            .I(N__49587));
    Span4Mux_v I__11443 (
            .O(N__49696),
            .I(N__49582));
    LocalMux I__11442 (
            .O(N__49693),
            .I(N__49582));
    LocalMux I__11441 (
            .O(N__49690),
            .I(N__49579));
    InMux I__11440 (
            .O(N__49689),
            .I(N__49576));
    LocalMux I__11439 (
            .O(N__49686),
            .I(N__49568));
    Span4Mux_h I__11438 (
            .O(N__49677),
            .I(N__49555));
    LocalMux I__11437 (
            .O(N__49674),
            .I(N__49555));
    LocalMux I__11436 (
            .O(N__49671),
            .I(N__49555));
    LocalMux I__11435 (
            .O(N__49668),
            .I(N__49555));
    LocalMux I__11434 (
            .O(N__49665),
            .I(N__49555));
    LocalMux I__11433 (
            .O(N__49662),
            .I(N__49555));
    InMux I__11432 (
            .O(N__49661),
            .I(N__49552));
    Span4Mux_v I__11431 (
            .O(N__49652),
            .I(N__49549));
    InMux I__11430 (
            .O(N__49651),
            .I(N__49546));
    Span4Mux_v I__11429 (
            .O(N__49646),
            .I(N__49533));
    Span4Mux_v I__11428 (
            .O(N__49639),
            .I(N__49533));
    LocalMux I__11427 (
            .O(N__49636),
            .I(N__49533));
    LocalMux I__11426 (
            .O(N__49633),
            .I(N__49533));
    LocalMux I__11425 (
            .O(N__49630),
            .I(N__49533));
    LocalMux I__11424 (
            .O(N__49627),
            .I(N__49533));
    InMux I__11423 (
            .O(N__49626),
            .I(N__49530));
    Span4Mux_v I__11422 (
            .O(N__49611),
            .I(N__49527));
    InMux I__11421 (
            .O(N__49610),
            .I(N__49524));
    InMux I__11420 (
            .O(N__49609),
            .I(N__49521));
    InMux I__11419 (
            .O(N__49608),
            .I(N__49518));
    Span4Mux_v I__11418 (
            .O(N__49605),
            .I(N__49515));
    Span4Mux_v I__11417 (
            .O(N__49602),
            .I(N__49506));
    LocalMux I__11416 (
            .O(N__49599),
            .I(N__49506));
    LocalMux I__11415 (
            .O(N__49596),
            .I(N__49506));
    LocalMux I__11414 (
            .O(N__49593),
            .I(N__49506));
    InMux I__11413 (
            .O(N__49592),
            .I(N__49503));
    InMux I__11412 (
            .O(N__49591),
            .I(N__49500));
    InMux I__11411 (
            .O(N__49590),
            .I(N__49497));
    Span4Mux_h I__11410 (
            .O(N__49587),
            .I(N__49493));
    Span4Mux_h I__11409 (
            .O(N__49582),
            .I(N__49486));
    Span4Mux_h I__11408 (
            .O(N__49579),
            .I(N__49486));
    LocalMux I__11407 (
            .O(N__49576),
            .I(N__49486));
    InMux I__11406 (
            .O(N__49575),
            .I(N__49483));
    InMux I__11405 (
            .O(N__49574),
            .I(N__49480));
    InMux I__11404 (
            .O(N__49573),
            .I(N__49477));
    InMux I__11403 (
            .O(N__49572),
            .I(N__49474));
    InMux I__11402 (
            .O(N__49571),
            .I(N__49471));
    Span4Mux_h I__11401 (
            .O(N__49568),
            .I(N__49464));
    Span4Mux_v I__11400 (
            .O(N__49555),
            .I(N__49464));
    LocalMux I__11399 (
            .O(N__49552),
            .I(N__49464));
    Span4Mux_h I__11398 (
            .O(N__49549),
            .I(N__49459));
    LocalMux I__11397 (
            .O(N__49546),
            .I(N__49459));
    Span4Mux_v I__11396 (
            .O(N__49533),
            .I(N__49454));
    LocalMux I__11395 (
            .O(N__49530),
            .I(N__49454));
    Span4Mux_v I__11394 (
            .O(N__49527),
            .I(N__49445));
    LocalMux I__11393 (
            .O(N__49524),
            .I(N__49445));
    LocalMux I__11392 (
            .O(N__49521),
            .I(N__49445));
    LocalMux I__11391 (
            .O(N__49518),
            .I(N__49445));
    Span4Mux_h I__11390 (
            .O(N__49515),
            .I(N__49434));
    Span4Mux_v I__11389 (
            .O(N__49506),
            .I(N__49434));
    LocalMux I__11388 (
            .O(N__49503),
            .I(N__49434));
    LocalMux I__11387 (
            .O(N__49500),
            .I(N__49434));
    LocalMux I__11386 (
            .O(N__49497),
            .I(N__49434));
    InMux I__11385 (
            .O(N__49496),
            .I(N__49431));
    Sp12to4 I__11384 (
            .O(N__49493),
            .I(N__49416));
    Sp12to4 I__11383 (
            .O(N__49486),
            .I(N__49416));
    LocalMux I__11382 (
            .O(N__49483),
            .I(N__49416));
    LocalMux I__11381 (
            .O(N__49480),
            .I(N__49416));
    LocalMux I__11380 (
            .O(N__49477),
            .I(N__49416));
    LocalMux I__11379 (
            .O(N__49474),
            .I(N__49416));
    LocalMux I__11378 (
            .O(N__49471),
            .I(N__49416));
    Span4Mux_h I__11377 (
            .O(N__49464),
            .I(N__49412));
    Span4Mux_v I__11376 (
            .O(N__49459),
            .I(N__49405));
    Span4Mux_h I__11375 (
            .O(N__49454),
            .I(N__49405));
    Span4Mux_v I__11374 (
            .O(N__49445),
            .I(N__49405));
    Span4Mux_v I__11373 (
            .O(N__49434),
            .I(N__49400));
    LocalMux I__11372 (
            .O(N__49431),
            .I(N__49400));
    Span12Mux_v I__11371 (
            .O(N__49416),
            .I(N__49397));
    InMux I__11370 (
            .O(N__49415),
            .I(N__49394));
    Odrv4 I__11369 (
            .O(N__49412),
            .I(spi_data_mosi_3));
    Odrv4 I__11368 (
            .O(N__49405),
            .I(spi_data_mosi_3));
    Odrv4 I__11367 (
            .O(N__49400),
            .I(spi_data_mosi_3));
    Odrv12 I__11366 (
            .O(N__49397),
            .I(spi_data_mosi_3));
    LocalMux I__11365 (
            .O(N__49394),
            .I(spi_data_mosi_3));
    InMux I__11364 (
            .O(N__49383),
            .I(N__49380));
    LocalMux I__11363 (
            .O(N__49380),
            .I(N__49377));
    Span4Mux_h I__11362 (
            .O(N__49377),
            .I(N__49374));
    Span4Mux_h I__11361 (
            .O(N__49374),
            .I(N__49371));
    Odrv4 I__11360 (
            .O(N__49371),
            .I(sDAC_mem_13Z0Z_3));
    InMux I__11359 (
            .O(N__49368),
            .I(N__49364));
    InMux I__11358 (
            .O(N__49367),
            .I(N__49351));
    LocalMux I__11357 (
            .O(N__49364),
            .I(N__49348));
    InMux I__11356 (
            .O(N__49363),
            .I(N__49340));
    InMux I__11355 (
            .O(N__49362),
            .I(N__49337));
    InMux I__11354 (
            .O(N__49361),
            .I(N__49331));
    InMux I__11353 (
            .O(N__49360),
            .I(N__49328));
    InMux I__11352 (
            .O(N__49359),
            .I(N__49323));
    InMux I__11351 (
            .O(N__49358),
            .I(N__49319));
    InMux I__11350 (
            .O(N__49357),
            .I(N__49316));
    InMux I__11349 (
            .O(N__49356),
            .I(N__49313));
    InMux I__11348 (
            .O(N__49355),
            .I(N__49309));
    InMux I__11347 (
            .O(N__49354),
            .I(N__49302));
    LocalMux I__11346 (
            .O(N__49351),
            .I(N__49297));
    Span4Mux_v I__11345 (
            .O(N__49348),
            .I(N__49297));
    InMux I__11344 (
            .O(N__49347),
            .I(N__49294));
    InMux I__11343 (
            .O(N__49346),
            .I(N__49291));
    InMux I__11342 (
            .O(N__49345),
            .I(N__49288));
    InMux I__11341 (
            .O(N__49344),
            .I(N__49285));
    InMux I__11340 (
            .O(N__49343),
            .I(N__49282));
    LocalMux I__11339 (
            .O(N__49340),
            .I(N__49276));
    LocalMux I__11338 (
            .O(N__49337),
            .I(N__49276));
    InMux I__11337 (
            .O(N__49336),
            .I(N__49273));
    InMux I__11336 (
            .O(N__49335),
            .I(N__49270));
    InMux I__11335 (
            .O(N__49334),
            .I(N__49267));
    LocalMux I__11334 (
            .O(N__49331),
            .I(N__49264));
    LocalMux I__11333 (
            .O(N__49328),
            .I(N__49261));
    InMux I__11332 (
            .O(N__49327),
            .I(N__49257));
    InMux I__11331 (
            .O(N__49326),
            .I(N__49254));
    LocalMux I__11330 (
            .O(N__49323),
            .I(N__49251));
    InMux I__11329 (
            .O(N__49322),
            .I(N__49248));
    LocalMux I__11328 (
            .O(N__49319),
            .I(N__49241));
    LocalMux I__11327 (
            .O(N__49316),
            .I(N__49241));
    LocalMux I__11326 (
            .O(N__49313),
            .I(N__49241));
    InMux I__11325 (
            .O(N__49312),
            .I(N__49238));
    LocalMux I__11324 (
            .O(N__49309),
            .I(N__49235));
    InMux I__11323 (
            .O(N__49308),
            .I(N__49232));
    InMux I__11322 (
            .O(N__49307),
            .I(N__49227));
    InMux I__11321 (
            .O(N__49306),
            .I(N__49223));
    InMux I__11320 (
            .O(N__49305),
            .I(N__49219));
    LocalMux I__11319 (
            .O(N__49302),
            .I(N__49208));
    Span4Mux_h I__11318 (
            .O(N__49297),
            .I(N__49208));
    LocalMux I__11317 (
            .O(N__49294),
            .I(N__49208));
    LocalMux I__11316 (
            .O(N__49291),
            .I(N__49208));
    LocalMux I__11315 (
            .O(N__49288),
            .I(N__49208));
    LocalMux I__11314 (
            .O(N__49285),
            .I(N__49202));
    LocalMux I__11313 (
            .O(N__49282),
            .I(N__49202));
    InMux I__11312 (
            .O(N__49281),
            .I(N__49199));
    Span4Mux_v I__11311 (
            .O(N__49276),
            .I(N__49190));
    LocalMux I__11310 (
            .O(N__49273),
            .I(N__49190));
    LocalMux I__11309 (
            .O(N__49270),
            .I(N__49190));
    LocalMux I__11308 (
            .O(N__49267),
            .I(N__49190));
    Span4Mux_h I__11307 (
            .O(N__49264),
            .I(N__49181));
    Span4Mux_v I__11306 (
            .O(N__49261),
            .I(N__49181));
    InMux I__11305 (
            .O(N__49260),
            .I(N__49178));
    LocalMux I__11304 (
            .O(N__49257),
            .I(N__49172));
    LocalMux I__11303 (
            .O(N__49254),
            .I(N__49172));
    Span4Mux_h I__11302 (
            .O(N__49251),
            .I(N__49167));
    LocalMux I__11301 (
            .O(N__49248),
            .I(N__49167));
    Span4Mux_v I__11300 (
            .O(N__49241),
            .I(N__49160));
    LocalMux I__11299 (
            .O(N__49238),
            .I(N__49160));
    Span4Mux_v I__11298 (
            .O(N__49235),
            .I(N__49155));
    LocalMux I__11297 (
            .O(N__49232),
            .I(N__49155));
    InMux I__11296 (
            .O(N__49231),
            .I(N__49152));
    InMux I__11295 (
            .O(N__49230),
            .I(N__49149));
    LocalMux I__11294 (
            .O(N__49227),
            .I(N__49146));
    InMux I__11293 (
            .O(N__49226),
            .I(N__49141));
    LocalMux I__11292 (
            .O(N__49223),
            .I(N__49138));
    InMux I__11291 (
            .O(N__49222),
            .I(N__49135));
    LocalMux I__11290 (
            .O(N__49219),
            .I(N__49132));
    Span4Mux_v I__11289 (
            .O(N__49208),
            .I(N__49126));
    InMux I__11288 (
            .O(N__49207),
            .I(N__49123));
    Span4Mux_v I__11287 (
            .O(N__49202),
            .I(N__49120));
    LocalMux I__11286 (
            .O(N__49199),
            .I(N__49115));
    Span4Mux_v I__11285 (
            .O(N__49190),
            .I(N__49115));
    InMux I__11284 (
            .O(N__49189),
            .I(N__49112));
    InMux I__11283 (
            .O(N__49188),
            .I(N__49106));
    InMux I__11282 (
            .O(N__49187),
            .I(N__49103));
    InMux I__11281 (
            .O(N__49186),
            .I(N__49100));
    Span4Mux_h I__11280 (
            .O(N__49181),
            .I(N__49095));
    LocalMux I__11279 (
            .O(N__49178),
            .I(N__49095));
    InMux I__11278 (
            .O(N__49177),
            .I(N__49092));
    Span4Mux_v I__11277 (
            .O(N__49172),
            .I(N__49088));
    Span4Mux_v I__11276 (
            .O(N__49167),
            .I(N__49085));
    InMux I__11275 (
            .O(N__49166),
            .I(N__49082));
    InMux I__11274 (
            .O(N__49165),
            .I(N__49079));
    Span4Mux_v I__11273 (
            .O(N__49160),
            .I(N__49068));
    Span4Mux_h I__11272 (
            .O(N__49155),
            .I(N__49068));
    LocalMux I__11271 (
            .O(N__49152),
            .I(N__49068));
    LocalMux I__11270 (
            .O(N__49149),
            .I(N__49063));
    Span4Mux_v I__11269 (
            .O(N__49146),
            .I(N__49063));
    InMux I__11268 (
            .O(N__49145),
            .I(N__49060));
    InMux I__11267 (
            .O(N__49144),
            .I(N__49057));
    LocalMux I__11266 (
            .O(N__49141),
            .I(N__49052));
    Span4Mux_h I__11265 (
            .O(N__49138),
            .I(N__49052));
    LocalMux I__11264 (
            .O(N__49135),
            .I(N__49047));
    Span4Mux_v I__11263 (
            .O(N__49132),
            .I(N__49047));
    InMux I__11262 (
            .O(N__49131),
            .I(N__49044));
    InMux I__11261 (
            .O(N__49130),
            .I(N__49041));
    InMux I__11260 (
            .O(N__49129),
            .I(N__49038));
    Sp12to4 I__11259 (
            .O(N__49126),
            .I(N__49035));
    LocalMux I__11258 (
            .O(N__49123),
            .I(N__49028));
    Sp12to4 I__11257 (
            .O(N__49120),
            .I(N__49028));
    Sp12to4 I__11256 (
            .O(N__49115),
            .I(N__49028));
    LocalMux I__11255 (
            .O(N__49112),
            .I(N__49025));
    InMux I__11254 (
            .O(N__49111),
            .I(N__49022));
    InMux I__11253 (
            .O(N__49110),
            .I(N__49019));
    InMux I__11252 (
            .O(N__49109),
            .I(N__49016));
    LocalMux I__11251 (
            .O(N__49106),
            .I(N__49009));
    LocalMux I__11250 (
            .O(N__49103),
            .I(N__49009));
    LocalMux I__11249 (
            .O(N__49100),
            .I(N__49009));
    Span4Mux_v I__11248 (
            .O(N__49095),
            .I(N__49004));
    LocalMux I__11247 (
            .O(N__49092),
            .I(N__49004));
    InMux I__11246 (
            .O(N__49091),
            .I(N__49001));
    Sp12to4 I__11245 (
            .O(N__49088),
            .I(N__48998));
    Sp12to4 I__11244 (
            .O(N__49085),
            .I(N__48993));
    LocalMux I__11243 (
            .O(N__49082),
            .I(N__48993));
    LocalMux I__11242 (
            .O(N__49079),
            .I(N__48990));
    InMux I__11241 (
            .O(N__49078),
            .I(N__48985));
    InMux I__11240 (
            .O(N__49077),
            .I(N__48982));
    InMux I__11239 (
            .O(N__49076),
            .I(N__48979));
    InMux I__11238 (
            .O(N__49075),
            .I(N__48976));
    Span4Mux_v I__11237 (
            .O(N__49068),
            .I(N__48973));
    Span4Mux_h I__11236 (
            .O(N__49063),
            .I(N__48962));
    LocalMux I__11235 (
            .O(N__49060),
            .I(N__48962));
    LocalMux I__11234 (
            .O(N__49057),
            .I(N__48962));
    Span4Mux_v I__11233 (
            .O(N__49052),
            .I(N__48962));
    Span4Mux_h I__11232 (
            .O(N__49047),
            .I(N__48962));
    LocalMux I__11231 (
            .O(N__49044),
            .I(N__48949));
    LocalMux I__11230 (
            .O(N__49041),
            .I(N__48949));
    LocalMux I__11229 (
            .O(N__49038),
            .I(N__48949));
    Span12Mux_h I__11228 (
            .O(N__49035),
            .I(N__48949));
    Span12Mux_h I__11227 (
            .O(N__49028),
            .I(N__48949));
    Span12Mux_h I__11226 (
            .O(N__49025),
            .I(N__48949));
    LocalMux I__11225 (
            .O(N__49022),
            .I(N__48930));
    LocalMux I__11224 (
            .O(N__49019),
            .I(N__48930));
    LocalMux I__11223 (
            .O(N__49016),
            .I(N__48930));
    Sp12to4 I__11222 (
            .O(N__49009),
            .I(N__48930));
    Sp12to4 I__11221 (
            .O(N__49004),
            .I(N__48930));
    LocalMux I__11220 (
            .O(N__49001),
            .I(N__48930));
    Span12Mux_s11_v I__11219 (
            .O(N__48998),
            .I(N__48930));
    Span12Mux_h I__11218 (
            .O(N__48993),
            .I(N__48930));
    Span12Mux_h I__11217 (
            .O(N__48990),
            .I(N__48930));
    InMux I__11216 (
            .O(N__48989),
            .I(N__48927));
    InMux I__11215 (
            .O(N__48988),
            .I(N__48924));
    LocalMux I__11214 (
            .O(N__48985),
            .I(N__48911));
    LocalMux I__11213 (
            .O(N__48982),
            .I(N__48911));
    LocalMux I__11212 (
            .O(N__48979),
            .I(N__48911));
    LocalMux I__11211 (
            .O(N__48976),
            .I(N__48911));
    Span4Mux_h I__11210 (
            .O(N__48973),
            .I(N__48911));
    Span4Mux_v I__11209 (
            .O(N__48962),
            .I(N__48911));
    Span12Mux_v I__11208 (
            .O(N__48949),
            .I(N__48907));
    Span12Mux_v I__11207 (
            .O(N__48930),
            .I(N__48904));
    LocalMux I__11206 (
            .O(N__48927),
            .I(N__48897));
    LocalMux I__11205 (
            .O(N__48924),
            .I(N__48897));
    Span4Mux_v I__11204 (
            .O(N__48911),
            .I(N__48897));
    InMux I__11203 (
            .O(N__48910),
            .I(N__48894));
    Odrv12 I__11202 (
            .O(N__48907),
            .I(spi_data_mosi_4));
    Odrv12 I__11201 (
            .O(N__48904),
            .I(spi_data_mosi_4));
    Odrv4 I__11200 (
            .O(N__48897),
            .I(spi_data_mosi_4));
    LocalMux I__11199 (
            .O(N__48894),
            .I(spi_data_mosi_4));
    InMux I__11198 (
            .O(N__48885),
            .I(N__48882));
    LocalMux I__11197 (
            .O(N__48882),
            .I(N__48879));
    Span4Mux_h I__11196 (
            .O(N__48879),
            .I(N__48876));
    Odrv4 I__11195 (
            .O(N__48876),
            .I(sDAC_mem_13Z0Z_4));
    InMux I__11194 (
            .O(N__48873),
            .I(N__48870));
    LocalMux I__11193 (
            .O(N__48870),
            .I(sDAC_mem_13Z0Z_7));
    CEMux I__11192 (
            .O(N__48867),
            .I(N__48863));
    CEMux I__11191 (
            .O(N__48866),
            .I(N__48860));
    LocalMux I__11190 (
            .O(N__48863),
            .I(N__48857));
    LocalMux I__11189 (
            .O(N__48860),
            .I(N__48854));
    Span4Mux_v I__11188 (
            .O(N__48857),
            .I(N__48851));
    Span4Mux_v I__11187 (
            .O(N__48854),
            .I(N__48848));
    Odrv4 I__11186 (
            .O(N__48851),
            .I(sDAC_mem_13_1_sqmuxa));
    Odrv4 I__11185 (
            .O(N__48848),
            .I(sDAC_mem_13_1_sqmuxa));
    InMux I__11184 (
            .O(N__48843),
            .I(N__48838));
    InMux I__11183 (
            .O(N__48842),
            .I(N__48835));
    InMux I__11182 (
            .O(N__48841),
            .I(N__48827));
    LocalMux I__11181 (
            .O(N__48838),
            .I(N__48822));
    LocalMux I__11180 (
            .O(N__48835),
            .I(N__48822));
    InMux I__11179 (
            .O(N__48834),
            .I(N__48819));
    InMux I__11178 (
            .O(N__48833),
            .I(N__48813));
    InMux I__11177 (
            .O(N__48832),
            .I(N__48809));
    InMux I__11176 (
            .O(N__48831),
            .I(N__48805));
    InMux I__11175 (
            .O(N__48830),
            .I(N__48802));
    LocalMux I__11174 (
            .O(N__48827),
            .I(N__48790));
    Span4Mux_h I__11173 (
            .O(N__48822),
            .I(N__48790));
    LocalMux I__11172 (
            .O(N__48819),
            .I(N__48790));
    InMux I__11171 (
            .O(N__48818),
            .I(N__48787));
    InMux I__11170 (
            .O(N__48817),
            .I(N__48783));
    InMux I__11169 (
            .O(N__48816),
            .I(N__48780));
    LocalMux I__11168 (
            .O(N__48813),
            .I(N__48773));
    InMux I__11167 (
            .O(N__48812),
            .I(N__48770));
    LocalMux I__11166 (
            .O(N__48809),
            .I(N__48765));
    InMux I__11165 (
            .O(N__48808),
            .I(N__48762));
    LocalMux I__11164 (
            .O(N__48805),
            .I(N__48757));
    LocalMux I__11163 (
            .O(N__48802),
            .I(N__48757));
    InMux I__11162 (
            .O(N__48801),
            .I(N__48754));
    InMux I__11161 (
            .O(N__48800),
            .I(N__48751));
    InMux I__11160 (
            .O(N__48799),
            .I(N__48748));
    InMux I__11159 (
            .O(N__48798),
            .I(N__48733));
    InMux I__11158 (
            .O(N__48797),
            .I(N__48730));
    Span4Mux_v I__11157 (
            .O(N__48790),
            .I(N__48723));
    LocalMux I__11156 (
            .O(N__48787),
            .I(N__48723));
    InMux I__11155 (
            .O(N__48786),
            .I(N__48720));
    LocalMux I__11154 (
            .O(N__48783),
            .I(N__48713));
    LocalMux I__11153 (
            .O(N__48780),
            .I(N__48713));
    InMux I__11152 (
            .O(N__48779),
            .I(N__48710));
    InMux I__11151 (
            .O(N__48778),
            .I(N__48707));
    InMux I__11150 (
            .O(N__48777),
            .I(N__48702));
    InMux I__11149 (
            .O(N__48776),
            .I(N__48699));
    Span4Mux_v I__11148 (
            .O(N__48773),
            .I(N__48694));
    LocalMux I__11147 (
            .O(N__48770),
            .I(N__48694));
    InMux I__11146 (
            .O(N__48769),
            .I(N__48691));
    InMux I__11145 (
            .O(N__48768),
            .I(N__48688));
    Span4Mux_h I__11144 (
            .O(N__48765),
            .I(N__48683));
    LocalMux I__11143 (
            .O(N__48762),
            .I(N__48683));
    Span4Mux_v I__11142 (
            .O(N__48757),
            .I(N__48678));
    LocalMux I__11141 (
            .O(N__48754),
            .I(N__48678));
    LocalMux I__11140 (
            .O(N__48751),
            .I(N__48673));
    LocalMux I__11139 (
            .O(N__48748),
            .I(N__48673));
    InMux I__11138 (
            .O(N__48747),
            .I(N__48664));
    InMux I__11137 (
            .O(N__48746),
            .I(N__48661));
    InMux I__11136 (
            .O(N__48745),
            .I(N__48658));
    InMux I__11135 (
            .O(N__48744),
            .I(N__48655));
    InMux I__11134 (
            .O(N__48743),
            .I(N__48652));
    InMux I__11133 (
            .O(N__48742),
            .I(N__48649));
    InMux I__11132 (
            .O(N__48741),
            .I(N__48646));
    InMux I__11131 (
            .O(N__48740),
            .I(N__48643));
    InMux I__11130 (
            .O(N__48739),
            .I(N__48640));
    InMux I__11129 (
            .O(N__48738),
            .I(N__48637));
    InMux I__11128 (
            .O(N__48737),
            .I(N__48634));
    InMux I__11127 (
            .O(N__48736),
            .I(N__48630));
    LocalMux I__11126 (
            .O(N__48733),
            .I(N__48627));
    LocalMux I__11125 (
            .O(N__48730),
            .I(N__48624));
    InMux I__11124 (
            .O(N__48729),
            .I(N__48621));
    InMux I__11123 (
            .O(N__48728),
            .I(N__48618));
    Span4Mux_v I__11122 (
            .O(N__48723),
            .I(N__48613));
    LocalMux I__11121 (
            .O(N__48720),
            .I(N__48613));
    InMux I__11120 (
            .O(N__48719),
            .I(N__48610));
    InMux I__11119 (
            .O(N__48718),
            .I(N__48607));
    Span4Mux_h I__11118 (
            .O(N__48713),
            .I(N__48600));
    LocalMux I__11117 (
            .O(N__48710),
            .I(N__48600));
    LocalMux I__11116 (
            .O(N__48707),
            .I(N__48600));
    InMux I__11115 (
            .O(N__48706),
            .I(N__48594));
    InMux I__11114 (
            .O(N__48705),
            .I(N__48589));
    LocalMux I__11113 (
            .O(N__48702),
            .I(N__48586));
    LocalMux I__11112 (
            .O(N__48699),
            .I(N__48583));
    Span4Mux_h I__11111 (
            .O(N__48694),
            .I(N__48580));
    LocalMux I__11110 (
            .O(N__48691),
            .I(N__48577));
    LocalMux I__11109 (
            .O(N__48688),
            .I(N__48572));
    Span4Mux_v I__11108 (
            .O(N__48683),
            .I(N__48569));
    Span4Mux_v I__11107 (
            .O(N__48678),
            .I(N__48564));
    Span4Mux_h I__11106 (
            .O(N__48673),
            .I(N__48564));
    CascadeMux I__11105 (
            .O(N__48672),
            .I(N__48561));
    InMux I__11104 (
            .O(N__48671),
            .I(N__48558));
    InMux I__11103 (
            .O(N__48670),
            .I(N__48555));
    InMux I__11102 (
            .O(N__48669),
            .I(N__48552));
    InMux I__11101 (
            .O(N__48668),
            .I(N__48549));
    InMux I__11100 (
            .O(N__48667),
            .I(N__48546));
    LocalMux I__11099 (
            .O(N__48664),
            .I(N__48540));
    LocalMux I__11098 (
            .O(N__48661),
            .I(N__48540));
    LocalMux I__11097 (
            .O(N__48658),
            .I(N__48531));
    LocalMux I__11096 (
            .O(N__48655),
            .I(N__48531));
    LocalMux I__11095 (
            .O(N__48652),
            .I(N__48531));
    LocalMux I__11094 (
            .O(N__48649),
            .I(N__48531));
    LocalMux I__11093 (
            .O(N__48646),
            .I(N__48520));
    LocalMux I__11092 (
            .O(N__48643),
            .I(N__48520));
    LocalMux I__11091 (
            .O(N__48640),
            .I(N__48520));
    LocalMux I__11090 (
            .O(N__48637),
            .I(N__48520));
    LocalMux I__11089 (
            .O(N__48634),
            .I(N__48520));
    InMux I__11088 (
            .O(N__48633),
            .I(N__48517));
    LocalMux I__11087 (
            .O(N__48630),
            .I(N__48512));
    Span4Mux_h I__11086 (
            .O(N__48627),
            .I(N__48512));
    Span4Mux_h I__11085 (
            .O(N__48624),
            .I(N__48507));
    LocalMux I__11084 (
            .O(N__48621),
            .I(N__48507));
    LocalMux I__11083 (
            .O(N__48618),
            .I(N__48502));
    Span4Mux_h I__11082 (
            .O(N__48613),
            .I(N__48502));
    LocalMux I__11081 (
            .O(N__48610),
            .I(N__48495));
    LocalMux I__11080 (
            .O(N__48607),
            .I(N__48495));
    Span4Mux_h I__11079 (
            .O(N__48600),
            .I(N__48495));
    InMux I__11078 (
            .O(N__48599),
            .I(N__48492));
    InMux I__11077 (
            .O(N__48598),
            .I(N__48489));
    InMux I__11076 (
            .O(N__48597),
            .I(N__48486));
    LocalMux I__11075 (
            .O(N__48594),
            .I(N__48483));
    InMux I__11074 (
            .O(N__48593),
            .I(N__48480));
    InMux I__11073 (
            .O(N__48592),
            .I(N__48477));
    LocalMux I__11072 (
            .O(N__48589),
            .I(N__48474));
    Span4Mux_h I__11071 (
            .O(N__48586),
            .I(N__48465));
    Span4Mux_v I__11070 (
            .O(N__48583),
            .I(N__48465));
    Span4Mux_h I__11069 (
            .O(N__48580),
            .I(N__48465));
    Span4Mux_h I__11068 (
            .O(N__48577),
            .I(N__48465));
    InMux I__11067 (
            .O(N__48576),
            .I(N__48462));
    InMux I__11066 (
            .O(N__48575),
            .I(N__48459));
    Span4Mux_h I__11065 (
            .O(N__48572),
            .I(N__48456));
    Sp12to4 I__11064 (
            .O(N__48569),
            .I(N__48453));
    Span4Mux_h I__11063 (
            .O(N__48564),
            .I(N__48450));
    InMux I__11062 (
            .O(N__48561),
            .I(N__48447));
    LocalMux I__11061 (
            .O(N__48558),
            .I(N__48436));
    LocalMux I__11060 (
            .O(N__48555),
            .I(N__48436));
    LocalMux I__11059 (
            .O(N__48552),
            .I(N__48436));
    LocalMux I__11058 (
            .O(N__48549),
            .I(N__48436));
    LocalMux I__11057 (
            .O(N__48546),
            .I(N__48436));
    InMux I__11056 (
            .O(N__48545),
            .I(N__48433));
    Span4Mux_v I__11055 (
            .O(N__48540),
            .I(N__48428));
    Span4Mux_v I__11054 (
            .O(N__48531),
            .I(N__48428));
    Span4Mux_v I__11053 (
            .O(N__48520),
            .I(N__48425));
    LocalMux I__11052 (
            .O(N__48517),
            .I(N__48420));
    Sp12to4 I__11051 (
            .O(N__48512),
            .I(N__48420));
    Sp12to4 I__11050 (
            .O(N__48507),
            .I(N__48413));
    Sp12to4 I__11049 (
            .O(N__48502),
            .I(N__48413));
    Sp12to4 I__11048 (
            .O(N__48495),
            .I(N__48413));
    LocalMux I__11047 (
            .O(N__48492),
            .I(N__48404));
    LocalMux I__11046 (
            .O(N__48489),
            .I(N__48404));
    LocalMux I__11045 (
            .O(N__48486),
            .I(N__48404));
    Span4Mux_h I__11044 (
            .O(N__48483),
            .I(N__48404));
    LocalMux I__11043 (
            .O(N__48480),
            .I(N__48401));
    LocalMux I__11042 (
            .O(N__48477),
            .I(N__48394));
    Span4Mux_v I__11041 (
            .O(N__48474),
            .I(N__48394));
    Span4Mux_h I__11040 (
            .O(N__48465),
            .I(N__48394));
    LocalMux I__11039 (
            .O(N__48462),
            .I(N__48381));
    LocalMux I__11038 (
            .O(N__48459),
            .I(N__48381));
    Sp12to4 I__11037 (
            .O(N__48456),
            .I(N__48381));
    Span12Mux_h I__11036 (
            .O(N__48453),
            .I(N__48381));
    Sp12to4 I__11035 (
            .O(N__48450),
            .I(N__48381));
    LocalMux I__11034 (
            .O(N__48447),
            .I(N__48381));
    Span12Mux_v I__11033 (
            .O(N__48436),
            .I(N__48378));
    LocalMux I__11032 (
            .O(N__48433),
            .I(N__48367));
    Sp12to4 I__11031 (
            .O(N__48428),
            .I(N__48367));
    Sp12to4 I__11030 (
            .O(N__48425),
            .I(N__48367));
    Span12Mux_v I__11029 (
            .O(N__48420),
            .I(N__48367));
    Span12Mux_v I__11028 (
            .O(N__48413),
            .I(N__48367));
    Sp12to4 I__11027 (
            .O(N__48404),
            .I(N__48358));
    Span12Mux_h I__11026 (
            .O(N__48401),
            .I(N__48358));
    Sp12to4 I__11025 (
            .O(N__48394),
            .I(N__48358));
    Span12Mux_v I__11024 (
            .O(N__48381),
            .I(N__48358));
    Odrv12 I__11023 (
            .O(N__48378),
            .I(spi_data_mosi_7));
    Odrv12 I__11022 (
            .O(N__48367),
            .I(spi_data_mosi_7));
    Odrv12 I__11021 (
            .O(N__48358),
            .I(spi_data_mosi_7));
    InMux I__11020 (
            .O(N__48351),
            .I(N__48348));
    LocalMux I__11019 (
            .O(N__48348),
            .I(N__48345));
    Odrv4 I__11018 (
            .O(N__48345),
            .I(sDAC_mem_12Z0Z_7));
    InMux I__11017 (
            .O(N__48342),
            .I(N__48333));
    InMux I__11016 (
            .O(N__48341),
            .I(N__48326));
    InMux I__11015 (
            .O(N__48340),
            .I(N__48321));
    InMux I__11014 (
            .O(N__48339),
            .I(N__48318));
    InMux I__11013 (
            .O(N__48338),
            .I(N__48315));
    InMux I__11012 (
            .O(N__48337),
            .I(N__48312));
    InMux I__11011 (
            .O(N__48336),
            .I(N__48307));
    LocalMux I__11010 (
            .O(N__48333),
            .I(N__48300));
    InMux I__11009 (
            .O(N__48332),
            .I(N__48297));
    InMux I__11008 (
            .O(N__48331),
            .I(N__48294));
    InMux I__11007 (
            .O(N__48330),
            .I(N__48291));
    InMux I__11006 (
            .O(N__48329),
            .I(N__48288));
    LocalMux I__11005 (
            .O(N__48326),
            .I(N__48285));
    InMux I__11004 (
            .O(N__48325),
            .I(N__48282));
    InMux I__11003 (
            .O(N__48324),
            .I(N__48275));
    LocalMux I__11002 (
            .O(N__48321),
            .I(N__48269));
    LocalMux I__11001 (
            .O(N__48318),
            .I(N__48262));
    LocalMux I__11000 (
            .O(N__48315),
            .I(N__48262));
    LocalMux I__10999 (
            .O(N__48312),
            .I(N__48262));
    InMux I__10998 (
            .O(N__48311),
            .I(N__48259));
    InMux I__10997 (
            .O(N__48310),
            .I(N__48256));
    LocalMux I__10996 (
            .O(N__48307),
            .I(N__48251));
    InMux I__10995 (
            .O(N__48306),
            .I(N__48248));
    InMux I__10994 (
            .O(N__48305),
            .I(N__48245));
    InMux I__10993 (
            .O(N__48304),
            .I(N__48241));
    InMux I__10992 (
            .O(N__48303),
            .I(N__48238));
    Span4Mux_v I__10991 (
            .O(N__48300),
            .I(N__48220));
    LocalMux I__10990 (
            .O(N__48297),
            .I(N__48220));
    LocalMux I__10989 (
            .O(N__48294),
            .I(N__48220));
    LocalMux I__10988 (
            .O(N__48291),
            .I(N__48215));
    LocalMux I__10987 (
            .O(N__48288),
            .I(N__48215));
    Span4Mux_v I__10986 (
            .O(N__48285),
            .I(N__48205));
    LocalMux I__10985 (
            .O(N__48282),
            .I(N__48205));
    InMux I__10984 (
            .O(N__48281),
            .I(N__48202));
    InMux I__10983 (
            .O(N__48280),
            .I(N__48199));
    InMux I__10982 (
            .O(N__48279),
            .I(N__48196));
    InMux I__10981 (
            .O(N__48278),
            .I(N__48193));
    LocalMux I__10980 (
            .O(N__48275),
            .I(N__48186));
    InMux I__10979 (
            .O(N__48274),
            .I(N__48183));
    InMux I__10978 (
            .O(N__48273),
            .I(N__48180));
    InMux I__10977 (
            .O(N__48272),
            .I(N__48177));
    Span4Mux_h I__10976 (
            .O(N__48269),
            .I(N__48168));
    Span4Mux_v I__10975 (
            .O(N__48262),
            .I(N__48168));
    LocalMux I__10974 (
            .O(N__48259),
            .I(N__48168));
    LocalMux I__10973 (
            .O(N__48256),
            .I(N__48168));
    InMux I__10972 (
            .O(N__48255),
            .I(N__48165));
    InMux I__10971 (
            .O(N__48254),
            .I(N__48162));
    Span4Mux_v I__10970 (
            .O(N__48251),
            .I(N__48154));
    LocalMux I__10969 (
            .O(N__48248),
            .I(N__48154));
    LocalMux I__10968 (
            .O(N__48245),
            .I(N__48150));
    InMux I__10967 (
            .O(N__48244),
            .I(N__48147));
    LocalMux I__10966 (
            .O(N__48241),
            .I(N__48143));
    LocalMux I__10965 (
            .O(N__48238),
            .I(N__48140));
    InMux I__10964 (
            .O(N__48237),
            .I(N__48137));
    InMux I__10963 (
            .O(N__48236),
            .I(N__48134));
    InMux I__10962 (
            .O(N__48235),
            .I(N__48131));
    InMux I__10961 (
            .O(N__48234),
            .I(N__48128));
    InMux I__10960 (
            .O(N__48233),
            .I(N__48125));
    InMux I__10959 (
            .O(N__48232),
            .I(N__48121));
    InMux I__10958 (
            .O(N__48231),
            .I(N__48118));
    InMux I__10957 (
            .O(N__48230),
            .I(N__48115));
    InMux I__10956 (
            .O(N__48229),
            .I(N__48112));
    InMux I__10955 (
            .O(N__48228),
            .I(N__48109));
    InMux I__10954 (
            .O(N__48227),
            .I(N__48106));
    Span4Mux_v I__10953 (
            .O(N__48220),
            .I(N__48101));
    Span4Mux_h I__10952 (
            .O(N__48215),
            .I(N__48101));
    InMux I__10951 (
            .O(N__48214),
            .I(N__48098));
    InMux I__10950 (
            .O(N__48213),
            .I(N__48095));
    InMux I__10949 (
            .O(N__48212),
            .I(N__48092));
    InMux I__10948 (
            .O(N__48211),
            .I(N__48089));
    InMux I__10947 (
            .O(N__48210),
            .I(N__48086));
    Span4Mux_v I__10946 (
            .O(N__48205),
            .I(N__48075));
    LocalMux I__10945 (
            .O(N__48202),
            .I(N__48075));
    LocalMux I__10944 (
            .O(N__48199),
            .I(N__48075));
    LocalMux I__10943 (
            .O(N__48196),
            .I(N__48075));
    LocalMux I__10942 (
            .O(N__48193),
            .I(N__48075));
    InMux I__10941 (
            .O(N__48192),
            .I(N__48072));
    InMux I__10940 (
            .O(N__48191),
            .I(N__48069));
    InMux I__10939 (
            .O(N__48190),
            .I(N__48066));
    InMux I__10938 (
            .O(N__48189),
            .I(N__48063));
    Span4Mux_h I__10937 (
            .O(N__48186),
            .I(N__48053));
    LocalMux I__10936 (
            .O(N__48183),
            .I(N__48053));
    LocalMux I__10935 (
            .O(N__48180),
            .I(N__48053));
    LocalMux I__10934 (
            .O(N__48177),
            .I(N__48053));
    Span4Mux_v I__10933 (
            .O(N__48168),
            .I(N__48046));
    LocalMux I__10932 (
            .O(N__48165),
            .I(N__48046));
    LocalMux I__10931 (
            .O(N__48162),
            .I(N__48046));
    InMux I__10930 (
            .O(N__48161),
            .I(N__48043));
    InMux I__10929 (
            .O(N__48160),
            .I(N__48040));
    InMux I__10928 (
            .O(N__48159),
            .I(N__48037));
    Span4Mux_v I__10927 (
            .O(N__48154),
            .I(N__48034));
    InMux I__10926 (
            .O(N__48153),
            .I(N__48031));
    Span4Mux_h I__10925 (
            .O(N__48150),
            .I(N__48026));
    LocalMux I__10924 (
            .O(N__48147),
            .I(N__48026));
    InMux I__10923 (
            .O(N__48146),
            .I(N__48023));
    Span4Mux_v I__10922 (
            .O(N__48143),
            .I(N__48014));
    Span4Mux_v I__10921 (
            .O(N__48140),
            .I(N__48014));
    LocalMux I__10920 (
            .O(N__48137),
            .I(N__48014));
    LocalMux I__10919 (
            .O(N__48134),
            .I(N__48014));
    LocalMux I__10918 (
            .O(N__48131),
            .I(N__48007));
    LocalMux I__10917 (
            .O(N__48128),
            .I(N__48007));
    LocalMux I__10916 (
            .O(N__48125),
            .I(N__48007));
    InMux I__10915 (
            .O(N__48124),
            .I(N__48004));
    LocalMux I__10914 (
            .O(N__48121),
            .I(N__48001));
    LocalMux I__10913 (
            .O(N__48118),
            .I(N__47996));
    LocalMux I__10912 (
            .O(N__48115),
            .I(N__47996));
    LocalMux I__10911 (
            .O(N__48112),
            .I(N__47989));
    LocalMux I__10910 (
            .O(N__48109),
            .I(N__47989));
    LocalMux I__10909 (
            .O(N__48106),
            .I(N__47989));
    Span4Mux_v I__10908 (
            .O(N__48101),
            .I(N__47976));
    LocalMux I__10907 (
            .O(N__48098),
            .I(N__47976));
    LocalMux I__10906 (
            .O(N__48095),
            .I(N__47976));
    LocalMux I__10905 (
            .O(N__48092),
            .I(N__47976));
    LocalMux I__10904 (
            .O(N__48089),
            .I(N__47976));
    LocalMux I__10903 (
            .O(N__48086),
            .I(N__47976));
    Span4Mux_v I__10902 (
            .O(N__48075),
            .I(N__47972));
    LocalMux I__10901 (
            .O(N__48072),
            .I(N__47963));
    LocalMux I__10900 (
            .O(N__48069),
            .I(N__47963));
    LocalMux I__10899 (
            .O(N__48066),
            .I(N__47963));
    LocalMux I__10898 (
            .O(N__48063),
            .I(N__47963));
    InMux I__10897 (
            .O(N__48062),
            .I(N__47960));
    Span4Mux_v I__10896 (
            .O(N__48053),
            .I(N__47949));
    Span4Mux_h I__10895 (
            .O(N__48046),
            .I(N__47949));
    LocalMux I__10894 (
            .O(N__48043),
            .I(N__47949));
    LocalMux I__10893 (
            .O(N__48040),
            .I(N__47949));
    LocalMux I__10892 (
            .O(N__48037),
            .I(N__47949));
    Sp12to4 I__10891 (
            .O(N__48034),
            .I(N__47943));
    LocalMux I__10890 (
            .O(N__48031),
            .I(N__47943));
    Span4Mux_v I__10889 (
            .O(N__48026),
            .I(N__47938));
    LocalMux I__10888 (
            .O(N__48023),
            .I(N__47938));
    Span4Mux_v I__10887 (
            .O(N__48014),
            .I(N__47931));
    Span4Mux_h I__10886 (
            .O(N__48007),
            .I(N__47931));
    LocalMux I__10885 (
            .O(N__48004),
            .I(N__47931));
    Span12Mux_h I__10884 (
            .O(N__48001),
            .I(N__47926));
    Span12Mux_s11_v I__10883 (
            .O(N__47996),
            .I(N__47926));
    Span4Mux_v I__10882 (
            .O(N__47989),
            .I(N__47923));
    Span4Mux_v I__10881 (
            .O(N__47976),
            .I(N__47920));
    InMux I__10880 (
            .O(N__47975),
            .I(N__47917));
    Span4Mux_h I__10879 (
            .O(N__47972),
            .I(N__47908));
    Span4Mux_v I__10878 (
            .O(N__47963),
            .I(N__47908));
    LocalMux I__10877 (
            .O(N__47960),
            .I(N__47908));
    Span4Mux_v I__10876 (
            .O(N__47949),
            .I(N__47908));
    CascadeMux I__10875 (
            .O(N__47948),
            .I(N__47905));
    Span12Mux_h I__10874 (
            .O(N__47943),
            .I(N__47902));
    Span4Mux_v I__10873 (
            .O(N__47938),
            .I(N__47899));
    Span4Mux_v I__10872 (
            .O(N__47931),
            .I(N__47896));
    Span12Mux_v I__10871 (
            .O(N__47926),
            .I(N__47887));
    Sp12to4 I__10870 (
            .O(N__47923),
            .I(N__47887));
    Sp12to4 I__10869 (
            .O(N__47920),
            .I(N__47887));
    LocalMux I__10868 (
            .O(N__47917),
            .I(N__47887));
    Span4Mux_h I__10867 (
            .O(N__47908),
            .I(N__47884));
    InMux I__10866 (
            .O(N__47905),
            .I(N__47881));
    Odrv12 I__10865 (
            .O(N__47902),
            .I(spi_data_mosi_6));
    Odrv4 I__10864 (
            .O(N__47899),
            .I(spi_data_mosi_6));
    Odrv4 I__10863 (
            .O(N__47896),
            .I(spi_data_mosi_6));
    Odrv12 I__10862 (
            .O(N__47887),
            .I(spi_data_mosi_6));
    Odrv4 I__10861 (
            .O(N__47884),
            .I(spi_data_mosi_6));
    LocalMux I__10860 (
            .O(N__47881),
            .I(spi_data_mosi_6));
    InMux I__10859 (
            .O(N__47868),
            .I(N__47865));
    LocalMux I__10858 (
            .O(N__47865),
            .I(N__47862));
    Span4Mux_h I__10857 (
            .O(N__47862),
            .I(N__47859));
    Span4Mux_h I__10856 (
            .O(N__47859),
            .I(N__47856));
    Odrv4 I__10855 (
            .O(N__47856),
            .I(sDAC_mem_12Z0Z_6));
    ClkMux I__10854 (
            .O(N__47853),
            .I(N__47397));
    ClkMux I__10853 (
            .O(N__47852),
            .I(N__47397));
    ClkMux I__10852 (
            .O(N__47851),
            .I(N__47397));
    ClkMux I__10851 (
            .O(N__47850),
            .I(N__47397));
    ClkMux I__10850 (
            .O(N__47849),
            .I(N__47397));
    ClkMux I__10849 (
            .O(N__47848),
            .I(N__47397));
    ClkMux I__10848 (
            .O(N__47847),
            .I(N__47397));
    ClkMux I__10847 (
            .O(N__47846),
            .I(N__47397));
    ClkMux I__10846 (
            .O(N__47845),
            .I(N__47397));
    ClkMux I__10845 (
            .O(N__47844),
            .I(N__47397));
    ClkMux I__10844 (
            .O(N__47843),
            .I(N__47397));
    ClkMux I__10843 (
            .O(N__47842),
            .I(N__47397));
    ClkMux I__10842 (
            .O(N__47841),
            .I(N__47397));
    ClkMux I__10841 (
            .O(N__47840),
            .I(N__47397));
    ClkMux I__10840 (
            .O(N__47839),
            .I(N__47397));
    ClkMux I__10839 (
            .O(N__47838),
            .I(N__47397));
    ClkMux I__10838 (
            .O(N__47837),
            .I(N__47397));
    ClkMux I__10837 (
            .O(N__47836),
            .I(N__47397));
    ClkMux I__10836 (
            .O(N__47835),
            .I(N__47397));
    ClkMux I__10835 (
            .O(N__47834),
            .I(N__47397));
    ClkMux I__10834 (
            .O(N__47833),
            .I(N__47397));
    ClkMux I__10833 (
            .O(N__47832),
            .I(N__47397));
    ClkMux I__10832 (
            .O(N__47831),
            .I(N__47397));
    ClkMux I__10831 (
            .O(N__47830),
            .I(N__47397));
    ClkMux I__10830 (
            .O(N__47829),
            .I(N__47397));
    ClkMux I__10829 (
            .O(N__47828),
            .I(N__47397));
    ClkMux I__10828 (
            .O(N__47827),
            .I(N__47397));
    ClkMux I__10827 (
            .O(N__47826),
            .I(N__47397));
    ClkMux I__10826 (
            .O(N__47825),
            .I(N__47397));
    ClkMux I__10825 (
            .O(N__47824),
            .I(N__47397));
    ClkMux I__10824 (
            .O(N__47823),
            .I(N__47397));
    ClkMux I__10823 (
            .O(N__47822),
            .I(N__47397));
    ClkMux I__10822 (
            .O(N__47821),
            .I(N__47397));
    ClkMux I__10821 (
            .O(N__47820),
            .I(N__47397));
    ClkMux I__10820 (
            .O(N__47819),
            .I(N__47397));
    ClkMux I__10819 (
            .O(N__47818),
            .I(N__47397));
    ClkMux I__10818 (
            .O(N__47817),
            .I(N__47397));
    ClkMux I__10817 (
            .O(N__47816),
            .I(N__47397));
    ClkMux I__10816 (
            .O(N__47815),
            .I(N__47397));
    ClkMux I__10815 (
            .O(N__47814),
            .I(N__47397));
    ClkMux I__10814 (
            .O(N__47813),
            .I(N__47397));
    ClkMux I__10813 (
            .O(N__47812),
            .I(N__47397));
    ClkMux I__10812 (
            .O(N__47811),
            .I(N__47397));
    ClkMux I__10811 (
            .O(N__47810),
            .I(N__47397));
    ClkMux I__10810 (
            .O(N__47809),
            .I(N__47397));
    ClkMux I__10809 (
            .O(N__47808),
            .I(N__47397));
    ClkMux I__10808 (
            .O(N__47807),
            .I(N__47397));
    ClkMux I__10807 (
            .O(N__47806),
            .I(N__47397));
    ClkMux I__10806 (
            .O(N__47805),
            .I(N__47397));
    ClkMux I__10805 (
            .O(N__47804),
            .I(N__47397));
    ClkMux I__10804 (
            .O(N__47803),
            .I(N__47397));
    ClkMux I__10803 (
            .O(N__47802),
            .I(N__47397));
    ClkMux I__10802 (
            .O(N__47801),
            .I(N__47397));
    ClkMux I__10801 (
            .O(N__47800),
            .I(N__47397));
    ClkMux I__10800 (
            .O(N__47799),
            .I(N__47397));
    ClkMux I__10799 (
            .O(N__47798),
            .I(N__47397));
    ClkMux I__10798 (
            .O(N__47797),
            .I(N__47397));
    ClkMux I__10797 (
            .O(N__47796),
            .I(N__47397));
    ClkMux I__10796 (
            .O(N__47795),
            .I(N__47397));
    ClkMux I__10795 (
            .O(N__47794),
            .I(N__47397));
    ClkMux I__10794 (
            .O(N__47793),
            .I(N__47397));
    ClkMux I__10793 (
            .O(N__47792),
            .I(N__47397));
    ClkMux I__10792 (
            .O(N__47791),
            .I(N__47397));
    ClkMux I__10791 (
            .O(N__47790),
            .I(N__47397));
    ClkMux I__10790 (
            .O(N__47789),
            .I(N__47397));
    ClkMux I__10789 (
            .O(N__47788),
            .I(N__47397));
    ClkMux I__10788 (
            .O(N__47787),
            .I(N__47397));
    ClkMux I__10787 (
            .O(N__47786),
            .I(N__47397));
    ClkMux I__10786 (
            .O(N__47785),
            .I(N__47397));
    ClkMux I__10785 (
            .O(N__47784),
            .I(N__47397));
    ClkMux I__10784 (
            .O(N__47783),
            .I(N__47397));
    ClkMux I__10783 (
            .O(N__47782),
            .I(N__47397));
    ClkMux I__10782 (
            .O(N__47781),
            .I(N__47397));
    ClkMux I__10781 (
            .O(N__47780),
            .I(N__47397));
    ClkMux I__10780 (
            .O(N__47779),
            .I(N__47397));
    ClkMux I__10779 (
            .O(N__47778),
            .I(N__47397));
    ClkMux I__10778 (
            .O(N__47777),
            .I(N__47397));
    ClkMux I__10777 (
            .O(N__47776),
            .I(N__47397));
    ClkMux I__10776 (
            .O(N__47775),
            .I(N__47397));
    ClkMux I__10775 (
            .O(N__47774),
            .I(N__47397));
    ClkMux I__10774 (
            .O(N__47773),
            .I(N__47397));
    ClkMux I__10773 (
            .O(N__47772),
            .I(N__47397));
    ClkMux I__10772 (
            .O(N__47771),
            .I(N__47397));
    ClkMux I__10771 (
            .O(N__47770),
            .I(N__47397));
    ClkMux I__10770 (
            .O(N__47769),
            .I(N__47397));
    ClkMux I__10769 (
            .O(N__47768),
            .I(N__47397));
    ClkMux I__10768 (
            .O(N__47767),
            .I(N__47397));
    ClkMux I__10767 (
            .O(N__47766),
            .I(N__47397));
    ClkMux I__10766 (
            .O(N__47765),
            .I(N__47397));
    ClkMux I__10765 (
            .O(N__47764),
            .I(N__47397));
    ClkMux I__10764 (
            .O(N__47763),
            .I(N__47397));
    ClkMux I__10763 (
            .O(N__47762),
            .I(N__47397));
    ClkMux I__10762 (
            .O(N__47761),
            .I(N__47397));
    ClkMux I__10761 (
            .O(N__47760),
            .I(N__47397));
    ClkMux I__10760 (
            .O(N__47759),
            .I(N__47397));
    ClkMux I__10759 (
            .O(N__47758),
            .I(N__47397));
    ClkMux I__10758 (
            .O(N__47757),
            .I(N__47397));
    ClkMux I__10757 (
            .O(N__47756),
            .I(N__47397));
    ClkMux I__10756 (
            .O(N__47755),
            .I(N__47397));
    ClkMux I__10755 (
            .O(N__47754),
            .I(N__47397));
    ClkMux I__10754 (
            .O(N__47753),
            .I(N__47397));
    ClkMux I__10753 (
            .O(N__47752),
            .I(N__47397));
    ClkMux I__10752 (
            .O(N__47751),
            .I(N__47397));
    ClkMux I__10751 (
            .O(N__47750),
            .I(N__47397));
    ClkMux I__10750 (
            .O(N__47749),
            .I(N__47397));
    ClkMux I__10749 (
            .O(N__47748),
            .I(N__47397));
    ClkMux I__10748 (
            .O(N__47747),
            .I(N__47397));
    ClkMux I__10747 (
            .O(N__47746),
            .I(N__47397));
    ClkMux I__10746 (
            .O(N__47745),
            .I(N__47397));
    ClkMux I__10745 (
            .O(N__47744),
            .I(N__47397));
    ClkMux I__10744 (
            .O(N__47743),
            .I(N__47397));
    ClkMux I__10743 (
            .O(N__47742),
            .I(N__47397));
    ClkMux I__10742 (
            .O(N__47741),
            .I(N__47397));
    ClkMux I__10741 (
            .O(N__47740),
            .I(N__47397));
    ClkMux I__10740 (
            .O(N__47739),
            .I(N__47397));
    ClkMux I__10739 (
            .O(N__47738),
            .I(N__47397));
    ClkMux I__10738 (
            .O(N__47737),
            .I(N__47397));
    ClkMux I__10737 (
            .O(N__47736),
            .I(N__47397));
    ClkMux I__10736 (
            .O(N__47735),
            .I(N__47397));
    ClkMux I__10735 (
            .O(N__47734),
            .I(N__47397));
    ClkMux I__10734 (
            .O(N__47733),
            .I(N__47397));
    ClkMux I__10733 (
            .O(N__47732),
            .I(N__47397));
    ClkMux I__10732 (
            .O(N__47731),
            .I(N__47397));
    ClkMux I__10731 (
            .O(N__47730),
            .I(N__47397));
    ClkMux I__10730 (
            .O(N__47729),
            .I(N__47397));
    ClkMux I__10729 (
            .O(N__47728),
            .I(N__47397));
    ClkMux I__10728 (
            .O(N__47727),
            .I(N__47397));
    ClkMux I__10727 (
            .O(N__47726),
            .I(N__47397));
    ClkMux I__10726 (
            .O(N__47725),
            .I(N__47397));
    ClkMux I__10725 (
            .O(N__47724),
            .I(N__47397));
    ClkMux I__10724 (
            .O(N__47723),
            .I(N__47397));
    ClkMux I__10723 (
            .O(N__47722),
            .I(N__47397));
    ClkMux I__10722 (
            .O(N__47721),
            .I(N__47397));
    ClkMux I__10721 (
            .O(N__47720),
            .I(N__47397));
    ClkMux I__10720 (
            .O(N__47719),
            .I(N__47397));
    ClkMux I__10719 (
            .O(N__47718),
            .I(N__47397));
    ClkMux I__10718 (
            .O(N__47717),
            .I(N__47397));
    ClkMux I__10717 (
            .O(N__47716),
            .I(N__47397));
    ClkMux I__10716 (
            .O(N__47715),
            .I(N__47397));
    ClkMux I__10715 (
            .O(N__47714),
            .I(N__47397));
    ClkMux I__10714 (
            .O(N__47713),
            .I(N__47397));
    ClkMux I__10713 (
            .O(N__47712),
            .I(N__47397));
    ClkMux I__10712 (
            .O(N__47711),
            .I(N__47397));
    ClkMux I__10711 (
            .O(N__47710),
            .I(N__47397));
    ClkMux I__10710 (
            .O(N__47709),
            .I(N__47397));
    ClkMux I__10709 (
            .O(N__47708),
            .I(N__47397));
    ClkMux I__10708 (
            .O(N__47707),
            .I(N__47397));
    ClkMux I__10707 (
            .O(N__47706),
            .I(N__47397));
    ClkMux I__10706 (
            .O(N__47705),
            .I(N__47397));
    ClkMux I__10705 (
            .O(N__47704),
            .I(N__47397));
    ClkMux I__10704 (
            .O(N__47703),
            .I(N__47397));
    ClkMux I__10703 (
            .O(N__47702),
            .I(N__47397));
    GlobalMux I__10702 (
            .O(N__47397),
            .I(N__47394));
    gio2CtrlBuf I__10701 (
            .O(N__47394),
            .I(pll_clk128_g));
    CEMux I__10700 (
            .O(N__47391),
            .I(N__47388));
    LocalMux I__10699 (
            .O(N__47388),
            .I(N__47385));
    Span4Mux_v I__10698 (
            .O(N__47385),
            .I(N__47381));
    CEMux I__10697 (
            .O(N__47384),
            .I(N__47378));
    Span4Mux_h I__10696 (
            .O(N__47381),
            .I(N__47372));
    LocalMux I__10695 (
            .O(N__47378),
            .I(N__47369));
    CEMux I__10694 (
            .O(N__47377),
            .I(N__47366));
    CEMux I__10693 (
            .O(N__47376),
            .I(N__47363));
    CEMux I__10692 (
            .O(N__47375),
            .I(N__47360));
    Span4Mux_h I__10691 (
            .O(N__47372),
            .I(N__47353));
    Span4Mux_h I__10690 (
            .O(N__47369),
            .I(N__47353));
    LocalMux I__10689 (
            .O(N__47366),
            .I(N__47353));
    LocalMux I__10688 (
            .O(N__47363),
            .I(N__47350));
    LocalMux I__10687 (
            .O(N__47360),
            .I(N__47347));
    Odrv4 I__10686 (
            .O(N__47353),
            .I(sDAC_mem_12_1_sqmuxa));
    Odrv4 I__10685 (
            .O(N__47350),
            .I(sDAC_mem_12_1_sqmuxa));
    Odrv4 I__10684 (
            .O(N__47347),
            .I(sDAC_mem_12_1_sqmuxa));
    InMux I__10683 (
            .O(N__47340),
            .I(N__47337));
    LocalMux I__10682 (
            .O(N__47337),
            .I(N__47334));
    Span4Mux_h I__10681 (
            .O(N__47334),
            .I(N__47331));
    Span4Mux_h I__10680 (
            .O(N__47331),
            .I(N__47328));
    Odrv4 I__10679 (
            .O(N__47328),
            .I(sDAC_mem_9Z0Z_7));
    CEMux I__10678 (
            .O(N__47325),
            .I(N__47322));
    LocalMux I__10677 (
            .O(N__47322),
            .I(N__47319));
    Span4Mux_v I__10676 (
            .O(N__47319),
            .I(N__47316));
    Odrv4 I__10675 (
            .O(N__47316),
            .I(sDAC_mem_9_1_sqmuxa));
    CascadeMux I__10674 (
            .O(N__47313),
            .I(N_14_3_cascade_));
    CascadeMux I__10673 (
            .O(N__47310),
            .I(N_8_cascade_));
    InMux I__10672 (
            .O(N__47307),
            .I(N__47301));
    InMux I__10671 (
            .O(N__47306),
            .I(N__47301));
    LocalMux I__10670 (
            .O(N__47301),
            .I(N__47297));
    InMux I__10669 (
            .O(N__47300),
            .I(N__47294));
    Span12Mux_h I__10668 (
            .O(N__47297),
            .I(N__47291));
    LocalMux I__10667 (
            .O(N__47294),
            .I(sDAC_spi_startZ0));
    Odrv12 I__10666 (
            .O(N__47291),
            .I(sDAC_spi_startZ0));
    InMux I__10665 (
            .O(N__47286),
            .I(N__47283));
    LocalMux I__10664 (
            .O(N__47283),
            .I(un1_scounterdac8_i_a2_1_2));
    InMux I__10663 (
            .O(N__47280),
            .I(N__47277));
    LocalMux I__10662 (
            .O(N__47277),
            .I(un1_scounterdac8_i_a2_0));
    InMux I__10661 (
            .O(N__47274),
            .I(N__47271));
    LocalMux I__10660 (
            .O(N__47271),
            .I(N__47268));
    Span4Mux_h I__10659 (
            .O(N__47268),
            .I(N__47265));
    Odrv4 I__10658 (
            .O(N__47265),
            .I(sDAC_data_RNO_18Z0Z_10));
    InMux I__10657 (
            .O(N__47262),
            .I(N__47259));
    LocalMux I__10656 (
            .O(N__47259),
            .I(N__47256));
    Span4Mux_h I__10655 (
            .O(N__47256),
            .I(N__47253));
    Odrv4 I__10654 (
            .O(N__47253),
            .I(sEEDACZ0Z_5));
    InMux I__10653 (
            .O(N__47250),
            .I(N__47247));
    LocalMux I__10652 (
            .O(N__47247),
            .I(N__47244));
    Span4Mux_h I__10651 (
            .O(N__47244),
            .I(N__47241));
    Odrv4 I__10650 (
            .O(N__47241),
            .I(sEEDACZ0Z_6));
    CEMux I__10649 (
            .O(N__47238),
            .I(N__47235));
    LocalMux I__10648 (
            .O(N__47235),
            .I(N__47231));
    CEMux I__10647 (
            .O(N__47234),
            .I(N__47228));
    Span4Mux_h I__10646 (
            .O(N__47231),
            .I(N__47225));
    LocalMux I__10645 (
            .O(N__47228),
            .I(N__47222));
    Odrv4 I__10644 (
            .O(N__47225),
            .I(sEEDAC_1_sqmuxa));
    Odrv4 I__10643 (
            .O(N__47222),
            .I(sEEDAC_1_sqmuxa));
    InMux I__10642 (
            .O(N__47217),
            .I(N__47214));
    LocalMux I__10641 (
            .O(N__47214),
            .I(N__47211));
    Span4Mux_h I__10640 (
            .O(N__47211),
            .I(N__47208));
    Odrv4 I__10639 (
            .O(N__47208),
            .I(sDAC_mem_9Z0Z_0));
    InMux I__10638 (
            .O(N__47205),
            .I(N__47202));
    LocalMux I__10637 (
            .O(N__47202),
            .I(N__47199));
    Span4Mux_v I__10636 (
            .O(N__47199),
            .I(N__47196));
    Odrv4 I__10635 (
            .O(N__47196),
            .I(sDAC_mem_9Z0Z_1));
    InMux I__10634 (
            .O(N__47193),
            .I(N__47190));
    LocalMux I__10633 (
            .O(N__47190),
            .I(N__47187));
    Span4Mux_h I__10632 (
            .O(N__47187),
            .I(N__47184));
    Span4Mux_h I__10631 (
            .O(N__47184),
            .I(N__47181));
    Odrv4 I__10630 (
            .O(N__47181),
            .I(sDAC_mem_9Z0Z_2));
    InMux I__10629 (
            .O(N__47178),
            .I(N__47175));
    LocalMux I__10628 (
            .O(N__47175),
            .I(N__47172));
    Span4Mux_h I__10627 (
            .O(N__47172),
            .I(N__47169));
    Odrv4 I__10626 (
            .O(N__47169),
            .I(sDAC_mem_9Z0Z_3));
    InMux I__10625 (
            .O(N__47166),
            .I(N__47163));
    LocalMux I__10624 (
            .O(N__47163),
            .I(N__47160));
    Span4Mux_h I__10623 (
            .O(N__47160),
            .I(N__47157));
    Span4Mux_h I__10622 (
            .O(N__47157),
            .I(N__47154));
    Odrv4 I__10621 (
            .O(N__47154),
            .I(sDAC_mem_9Z0Z_4));
    InMux I__10620 (
            .O(N__47151),
            .I(N__47144));
    InMux I__10619 (
            .O(N__47150),
            .I(N__47141));
    InMux I__10618 (
            .O(N__47149),
            .I(N__47127));
    InMux I__10617 (
            .O(N__47148),
            .I(N__47123));
    InMux I__10616 (
            .O(N__47147),
            .I(N__47120));
    LocalMux I__10615 (
            .O(N__47144),
            .I(N__47112));
    LocalMux I__10614 (
            .O(N__47141),
            .I(N__47112));
    InMux I__10613 (
            .O(N__47140),
            .I(N__47109));
    InMux I__10612 (
            .O(N__47139),
            .I(N__47106));
    InMux I__10611 (
            .O(N__47138),
            .I(N__47103));
    InMux I__10610 (
            .O(N__47137),
            .I(N__47100));
    InMux I__10609 (
            .O(N__47136),
            .I(N__47096));
    InMux I__10608 (
            .O(N__47135),
            .I(N__47093));
    InMux I__10607 (
            .O(N__47134),
            .I(N__47090));
    InMux I__10606 (
            .O(N__47133),
            .I(N__47085));
    InMux I__10605 (
            .O(N__47132),
            .I(N__47082));
    InMux I__10604 (
            .O(N__47131),
            .I(N__47078));
    InMux I__10603 (
            .O(N__47130),
            .I(N__47075));
    LocalMux I__10602 (
            .O(N__47127),
            .I(N__47068));
    InMux I__10601 (
            .O(N__47126),
            .I(N__47065));
    LocalMux I__10600 (
            .O(N__47123),
            .I(N__47057));
    LocalMux I__10599 (
            .O(N__47120),
            .I(N__47057));
    InMux I__10598 (
            .O(N__47119),
            .I(N__47054));
    InMux I__10597 (
            .O(N__47118),
            .I(N__47050));
    InMux I__10596 (
            .O(N__47117),
            .I(N__47047));
    Span4Mux_v I__10595 (
            .O(N__47112),
            .I(N__47034));
    LocalMux I__10594 (
            .O(N__47109),
            .I(N__47034));
    LocalMux I__10593 (
            .O(N__47106),
            .I(N__47034));
    LocalMux I__10592 (
            .O(N__47103),
            .I(N__47034));
    LocalMux I__10591 (
            .O(N__47100),
            .I(N__47034));
    InMux I__10590 (
            .O(N__47099),
            .I(N__47031));
    LocalMux I__10589 (
            .O(N__47096),
            .I(N__47024));
    LocalMux I__10588 (
            .O(N__47093),
            .I(N__47024));
    LocalMux I__10587 (
            .O(N__47090),
            .I(N__47024));
    InMux I__10586 (
            .O(N__47089),
            .I(N__47021));
    InMux I__10585 (
            .O(N__47088),
            .I(N__47018));
    LocalMux I__10584 (
            .O(N__47085),
            .I(N__47013));
    LocalMux I__10583 (
            .O(N__47082),
            .I(N__47010));
    InMux I__10582 (
            .O(N__47081),
            .I(N__47007));
    LocalMux I__10581 (
            .O(N__47078),
            .I(N__47004));
    LocalMux I__10580 (
            .O(N__47075),
            .I(N__47001));
    InMux I__10579 (
            .O(N__47074),
            .I(N__46998));
    InMux I__10578 (
            .O(N__47073),
            .I(N__46995));
    InMux I__10577 (
            .O(N__47072),
            .I(N__46990));
    InMux I__10576 (
            .O(N__47071),
            .I(N__46987));
    Span4Mux_h I__10575 (
            .O(N__47068),
            .I(N__46980));
    LocalMux I__10574 (
            .O(N__47065),
            .I(N__46977));
    InMux I__10573 (
            .O(N__47064),
            .I(N__46974));
    InMux I__10572 (
            .O(N__47063),
            .I(N__46971));
    InMux I__10571 (
            .O(N__47062),
            .I(N__46967));
    Span4Mux_h I__10570 (
            .O(N__47057),
            .I(N__46962));
    LocalMux I__10569 (
            .O(N__47054),
            .I(N__46962));
    InMux I__10568 (
            .O(N__47053),
            .I(N__46959));
    LocalMux I__10567 (
            .O(N__47050),
            .I(N__46953));
    LocalMux I__10566 (
            .O(N__47047),
            .I(N__46950));
    InMux I__10565 (
            .O(N__47046),
            .I(N__46947));
    InMux I__10564 (
            .O(N__47045),
            .I(N__46944));
    Span4Mux_v I__10563 (
            .O(N__47034),
            .I(N__46939));
    LocalMux I__10562 (
            .O(N__47031),
            .I(N__46939));
    Span4Mux_v I__10561 (
            .O(N__47024),
            .I(N__46934));
    LocalMux I__10560 (
            .O(N__47021),
            .I(N__46934));
    LocalMux I__10559 (
            .O(N__47018),
            .I(N__46931));
    InMux I__10558 (
            .O(N__47017),
            .I(N__46928));
    InMux I__10557 (
            .O(N__47016),
            .I(N__46925));
    Span4Mux_v I__10556 (
            .O(N__47013),
            .I(N__46918));
    Span4Mux_h I__10555 (
            .O(N__47010),
            .I(N__46918));
    LocalMux I__10554 (
            .O(N__47007),
            .I(N__46918));
    Span4Mux_h I__10553 (
            .O(N__47004),
            .I(N__46913));
    Span4Mux_h I__10552 (
            .O(N__47001),
            .I(N__46913));
    LocalMux I__10551 (
            .O(N__46998),
            .I(N__46908));
    LocalMux I__10550 (
            .O(N__46995),
            .I(N__46908));
    InMux I__10549 (
            .O(N__46994),
            .I(N__46905));
    InMux I__10548 (
            .O(N__46993),
            .I(N__46902));
    LocalMux I__10547 (
            .O(N__46990),
            .I(N__46899));
    LocalMux I__10546 (
            .O(N__46987),
            .I(N__46894));
    InMux I__10545 (
            .O(N__46986),
            .I(N__46891));
    InMux I__10544 (
            .O(N__46985),
            .I(N__46888));
    InMux I__10543 (
            .O(N__46984),
            .I(N__46885));
    InMux I__10542 (
            .O(N__46983),
            .I(N__46882));
    Span4Mux_v I__10541 (
            .O(N__46980),
            .I(N__46871));
    Span4Mux_h I__10540 (
            .O(N__46977),
            .I(N__46871));
    LocalMux I__10539 (
            .O(N__46974),
            .I(N__46868));
    LocalMux I__10538 (
            .O(N__46971),
            .I(N__46865));
    InMux I__10537 (
            .O(N__46970),
            .I(N__46862));
    LocalMux I__10536 (
            .O(N__46967),
            .I(N__46858));
    Span4Mux_h I__10535 (
            .O(N__46962),
            .I(N__46853));
    LocalMux I__10534 (
            .O(N__46959),
            .I(N__46853));
    InMux I__10533 (
            .O(N__46958),
            .I(N__46850));
    InMux I__10532 (
            .O(N__46957),
            .I(N__46845));
    InMux I__10531 (
            .O(N__46956),
            .I(N__46845));
    Span4Mux_h I__10530 (
            .O(N__46953),
            .I(N__46842));
    Span4Mux_h I__10529 (
            .O(N__46950),
            .I(N__46835));
    LocalMux I__10528 (
            .O(N__46947),
            .I(N__46835));
    LocalMux I__10527 (
            .O(N__46944),
            .I(N__46835));
    Span4Mux_h I__10526 (
            .O(N__46939),
            .I(N__46832));
    Span4Mux_v I__10525 (
            .O(N__46934),
            .I(N__46823));
    Span4Mux_h I__10524 (
            .O(N__46931),
            .I(N__46823));
    LocalMux I__10523 (
            .O(N__46928),
            .I(N__46823));
    LocalMux I__10522 (
            .O(N__46925),
            .I(N__46823));
    Span4Mux_v I__10521 (
            .O(N__46918),
            .I(N__46820));
    Span4Mux_v I__10520 (
            .O(N__46913),
            .I(N__46811));
    Span4Mux_h I__10519 (
            .O(N__46908),
            .I(N__46811));
    LocalMux I__10518 (
            .O(N__46905),
            .I(N__46811));
    LocalMux I__10517 (
            .O(N__46902),
            .I(N__46811));
    Span4Mux_h I__10516 (
            .O(N__46899),
            .I(N__46808));
    InMux I__10515 (
            .O(N__46898),
            .I(N__46805));
    InMux I__10514 (
            .O(N__46897),
            .I(N__46802));
    Span4Mux_h I__10513 (
            .O(N__46894),
            .I(N__46795));
    LocalMux I__10512 (
            .O(N__46891),
            .I(N__46795));
    LocalMux I__10511 (
            .O(N__46888),
            .I(N__46795));
    LocalMux I__10510 (
            .O(N__46885),
            .I(N__46788));
    LocalMux I__10509 (
            .O(N__46882),
            .I(N__46788));
    InMux I__10508 (
            .O(N__46881),
            .I(N__46785));
    InMux I__10507 (
            .O(N__46880),
            .I(N__46782));
    InMux I__10506 (
            .O(N__46879),
            .I(N__46779));
    InMux I__10505 (
            .O(N__46878),
            .I(N__46776));
    InMux I__10504 (
            .O(N__46877),
            .I(N__46773));
    InMux I__10503 (
            .O(N__46876),
            .I(N__46770));
    Span4Mux_v I__10502 (
            .O(N__46871),
            .I(N__46766));
    Span4Mux_v I__10501 (
            .O(N__46868),
            .I(N__46759));
    Span4Mux_v I__10500 (
            .O(N__46865),
            .I(N__46759));
    LocalMux I__10499 (
            .O(N__46862),
            .I(N__46759));
    InMux I__10498 (
            .O(N__46861),
            .I(N__46756));
    Span4Mux_h I__10497 (
            .O(N__46858),
            .I(N__46747));
    Span4Mux_v I__10496 (
            .O(N__46853),
            .I(N__46747));
    LocalMux I__10495 (
            .O(N__46850),
            .I(N__46747));
    LocalMux I__10494 (
            .O(N__46845),
            .I(N__46747));
    Span4Mux_h I__10493 (
            .O(N__46842),
            .I(N__46738));
    Span4Mux_v I__10492 (
            .O(N__46835),
            .I(N__46738));
    Span4Mux_h I__10491 (
            .O(N__46832),
            .I(N__46738));
    Span4Mux_h I__10490 (
            .O(N__46823),
            .I(N__46738));
    Span4Mux_h I__10489 (
            .O(N__46820),
            .I(N__46733));
    Span4Mux_v I__10488 (
            .O(N__46811),
            .I(N__46733));
    Span4Mux_h I__10487 (
            .O(N__46808),
            .I(N__46726));
    LocalMux I__10486 (
            .O(N__46805),
            .I(N__46726));
    LocalMux I__10485 (
            .O(N__46802),
            .I(N__46726));
    Span4Mux_v I__10484 (
            .O(N__46795),
            .I(N__46723));
    InMux I__10483 (
            .O(N__46794),
            .I(N__46720));
    InMux I__10482 (
            .O(N__46793),
            .I(N__46717));
    Span4Mux_h I__10481 (
            .O(N__46788),
            .I(N__46702));
    LocalMux I__10480 (
            .O(N__46785),
            .I(N__46702));
    LocalMux I__10479 (
            .O(N__46782),
            .I(N__46702));
    LocalMux I__10478 (
            .O(N__46779),
            .I(N__46702));
    LocalMux I__10477 (
            .O(N__46776),
            .I(N__46702));
    LocalMux I__10476 (
            .O(N__46773),
            .I(N__46702));
    LocalMux I__10475 (
            .O(N__46770),
            .I(N__46702));
    InMux I__10474 (
            .O(N__46769),
            .I(N__46699));
    Span4Mux_v I__10473 (
            .O(N__46766),
            .I(N__46690));
    Span4Mux_h I__10472 (
            .O(N__46759),
            .I(N__46690));
    LocalMux I__10471 (
            .O(N__46756),
            .I(N__46690));
    Span4Mux_v I__10470 (
            .O(N__46747),
            .I(N__46690));
    Span4Mux_v I__10469 (
            .O(N__46738),
            .I(N__46687));
    Span4Mux_v I__10468 (
            .O(N__46733),
            .I(N__46676));
    Span4Mux_v I__10467 (
            .O(N__46726),
            .I(N__46676));
    Span4Mux_h I__10466 (
            .O(N__46723),
            .I(N__46676));
    LocalMux I__10465 (
            .O(N__46720),
            .I(N__46676));
    LocalMux I__10464 (
            .O(N__46717),
            .I(N__46676));
    Span4Mux_v I__10463 (
            .O(N__46702),
            .I(N__46669));
    LocalMux I__10462 (
            .O(N__46699),
            .I(N__46669));
    Span4Mux_v I__10461 (
            .O(N__46690),
            .I(N__46669));
    Odrv4 I__10460 (
            .O(N__46687),
            .I(spi_data_mosi_5));
    Odrv4 I__10459 (
            .O(N__46676),
            .I(spi_data_mosi_5));
    Odrv4 I__10458 (
            .O(N__46669),
            .I(spi_data_mosi_5));
    InMux I__10457 (
            .O(N__46662),
            .I(N__46659));
    LocalMux I__10456 (
            .O(N__46659),
            .I(N__46656));
    Span4Mux_v I__10455 (
            .O(N__46656),
            .I(N__46653));
    Odrv4 I__10454 (
            .O(N__46653),
            .I(sDAC_mem_9Z0Z_5));
    InMux I__10453 (
            .O(N__46650),
            .I(N__46647));
    LocalMux I__10452 (
            .O(N__46647),
            .I(N__46644));
    Span4Mux_h I__10451 (
            .O(N__46644),
            .I(N__46641));
    Span4Mux_h I__10450 (
            .O(N__46641),
            .I(N__46638));
    Odrv4 I__10449 (
            .O(N__46638),
            .I(sDAC_mem_9Z0Z_6));
    CEMux I__10448 (
            .O(N__46635),
            .I(N__46632));
    LocalMux I__10447 (
            .O(N__46632),
            .I(N__46626));
    CEMux I__10446 (
            .O(N__46631),
            .I(N__46623));
    CEMux I__10445 (
            .O(N__46630),
            .I(N__46620));
    CEMux I__10444 (
            .O(N__46629),
            .I(N__46617));
    Span4Mux_v I__10443 (
            .O(N__46626),
            .I(N__46614));
    LocalMux I__10442 (
            .O(N__46623),
            .I(N__46611));
    LocalMux I__10441 (
            .O(N__46620),
            .I(N__46608));
    LocalMux I__10440 (
            .O(N__46617),
            .I(N__46605));
    Span4Mux_h I__10439 (
            .O(N__46614),
            .I(N__46598));
    Span4Mux_v I__10438 (
            .O(N__46611),
            .I(N__46598));
    Span4Mux_v I__10437 (
            .O(N__46608),
            .I(N__46598));
    Span4Mux_h I__10436 (
            .O(N__46605),
            .I(N__46595));
    Span4Mux_v I__10435 (
            .O(N__46598),
            .I(N__46590));
    Span4Mux_h I__10434 (
            .O(N__46595),
            .I(N__46590));
    Odrv4 I__10433 (
            .O(N__46590),
            .I(sDAC_mem_16_1_sqmuxa));
    InMux I__10432 (
            .O(N__46587),
            .I(N__46584));
    LocalMux I__10431 (
            .O(N__46584),
            .I(N__46581));
    Span12Mux_v I__10430 (
            .O(N__46581),
            .I(N__46578));
    Odrv12 I__10429 (
            .O(N__46578),
            .I(sEEDACZ0Z_7));
    CascadeMux I__10428 (
            .O(N__46575),
            .I(N__46570));
    InMux I__10427 (
            .O(N__46574),
            .I(N__46560));
    InMux I__10426 (
            .O(N__46573),
            .I(N__46556));
    InMux I__10425 (
            .O(N__46570),
            .I(N__46551));
    InMux I__10424 (
            .O(N__46569),
            .I(N__46551));
    InMux I__10423 (
            .O(N__46568),
            .I(N__46538));
    InMux I__10422 (
            .O(N__46567),
            .I(N__46538));
    InMux I__10421 (
            .O(N__46566),
            .I(N__46538));
    InMux I__10420 (
            .O(N__46565),
            .I(N__46538));
    InMux I__10419 (
            .O(N__46564),
            .I(N__46538));
    InMux I__10418 (
            .O(N__46563),
            .I(N__46538));
    LocalMux I__10417 (
            .O(N__46560),
            .I(N__46535));
    InMux I__10416 (
            .O(N__46559),
            .I(N__46532));
    LocalMux I__10415 (
            .O(N__46556),
            .I(N__46529));
    LocalMux I__10414 (
            .O(N__46551),
            .I(N__46525));
    LocalMux I__10413 (
            .O(N__46538),
            .I(N__46522));
    Span4Mux_v I__10412 (
            .O(N__46535),
            .I(N__46519));
    LocalMux I__10411 (
            .O(N__46532),
            .I(N__46514));
    Span4Mux_v I__10410 (
            .O(N__46529),
            .I(N__46514));
    InMux I__10409 (
            .O(N__46528),
            .I(N__46508));
    Span4Mux_h I__10408 (
            .O(N__46525),
            .I(N__46505));
    Span4Mux_h I__10407 (
            .O(N__46522),
            .I(N__46502));
    Span4Mux_v I__10406 (
            .O(N__46519),
            .I(N__46497));
    Span4Mux_h I__10405 (
            .O(N__46514),
            .I(N__46497));
    InMux I__10404 (
            .O(N__46513),
            .I(N__46490));
    InMux I__10403 (
            .O(N__46512),
            .I(N__46490));
    InMux I__10402 (
            .O(N__46511),
            .I(N__46490));
    LocalMux I__10401 (
            .O(N__46508),
            .I(N__46487));
    Span4Mux_h I__10400 (
            .O(N__46505),
            .I(N__46482));
    Span4Mux_h I__10399 (
            .O(N__46502),
            .I(N__46479));
    Span4Mux_h I__10398 (
            .O(N__46497),
            .I(N__46474));
    LocalMux I__10397 (
            .O(N__46490),
            .I(N__46474));
    Span12Mux_v I__10396 (
            .O(N__46487),
            .I(N__46471));
    InMux I__10395 (
            .O(N__46486),
            .I(N__46468));
    InMux I__10394 (
            .O(N__46485),
            .I(N__46465));
    Odrv4 I__10393 (
            .O(N__46482),
            .I(sAddressZ0Z_5));
    Odrv4 I__10392 (
            .O(N__46479),
            .I(sAddressZ0Z_5));
    Odrv4 I__10391 (
            .O(N__46474),
            .I(sAddressZ0Z_5));
    Odrv12 I__10390 (
            .O(N__46471),
            .I(sAddressZ0Z_5));
    LocalMux I__10389 (
            .O(N__46468),
            .I(sAddressZ0Z_5));
    LocalMux I__10388 (
            .O(N__46465),
            .I(sAddressZ0Z_5));
    CascadeMux I__10387 (
            .O(N__46452),
            .I(N__46446));
    InMux I__10386 (
            .O(N__46451),
            .I(N__46442));
    CascadeMux I__10385 (
            .O(N__46450),
            .I(N__46439));
    CascadeMux I__10384 (
            .O(N__46449),
            .I(N__46435));
    InMux I__10383 (
            .O(N__46446),
            .I(N__46432));
    CascadeMux I__10382 (
            .O(N__46445),
            .I(N__46429));
    LocalMux I__10381 (
            .O(N__46442),
            .I(N__46425));
    InMux I__10380 (
            .O(N__46439),
            .I(N__46422));
    InMux I__10379 (
            .O(N__46438),
            .I(N__46419));
    InMux I__10378 (
            .O(N__46435),
            .I(N__46415));
    LocalMux I__10377 (
            .O(N__46432),
            .I(N__46409));
    InMux I__10376 (
            .O(N__46429),
            .I(N__46406));
    InMux I__10375 (
            .O(N__46428),
            .I(N__46403));
    Span4Mux_v I__10374 (
            .O(N__46425),
            .I(N__46398));
    LocalMux I__10373 (
            .O(N__46422),
            .I(N__46398));
    LocalMux I__10372 (
            .O(N__46419),
            .I(N__46395));
    InMux I__10371 (
            .O(N__46418),
            .I(N__46392));
    LocalMux I__10370 (
            .O(N__46415),
            .I(N__46389));
    InMux I__10369 (
            .O(N__46414),
            .I(N__46382));
    InMux I__10368 (
            .O(N__46413),
            .I(N__46382));
    InMux I__10367 (
            .O(N__46412),
            .I(N__46382));
    Span4Mux_h I__10366 (
            .O(N__46409),
            .I(N__46379));
    LocalMux I__10365 (
            .O(N__46406),
            .I(N__46376));
    LocalMux I__10364 (
            .O(N__46403),
            .I(N__46373));
    Span4Mux_h I__10363 (
            .O(N__46398),
            .I(N__46368));
    Span4Mux_v I__10362 (
            .O(N__46395),
            .I(N__46368));
    LocalMux I__10361 (
            .O(N__46392),
            .I(N__46365));
    Span4Mux_h I__10360 (
            .O(N__46389),
            .I(N__46362));
    LocalMux I__10359 (
            .O(N__46382),
            .I(N__46359));
    Span4Mux_v I__10358 (
            .O(N__46379),
            .I(N__46354));
    Span4Mux_h I__10357 (
            .O(N__46376),
            .I(N__46354));
    Span4Mux_v I__10356 (
            .O(N__46373),
            .I(N__46351));
    Span4Mux_v I__10355 (
            .O(N__46368),
            .I(N__46348));
    Span4Mux_h I__10354 (
            .O(N__46365),
            .I(N__46341));
    Span4Mux_v I__10353 (
            .O(N__46362),
            .I(N__46341));
    Span4Mux_h I__10352 (
            .O(N__46359),
            .I(N__46341));
    Span4Mux_v I__10351 (
            .O(N__46354),
            .I(N__46334));
    Span4Mux_h I__10350 (
            .O(N__46351),
            .I(N__46334));
    Span4Mux_h I__10349 (
            .O(N__46348),
            .I(N__46334));
    Odrv4 I__10348 (
            .O(N__46341),
            .I(N_139));
    Odrv4 I__10347 (
            .O(N__46334),
            .I(N_139));
    InMux I__10346 (
            .O(N__46329),
            .I(N__46323));
    InMux I__10345 (
            .O(N__46328),
            .I(N__46323));
    LocalMux I__10344 (
            .O(N__46323),
            .I(N__46316));
    InMux I__10343 (
            .O(N__46322),
            .I(N__46313));
    InMux I__10342 (
            .O(N__46321),
            .I(N__46308));
    InMux I__10341 (
            .O(N__46320),
            .I(N__46308));
    InMux I__10340 (
            .O(N__46319),
            .I(N__46305));
    Span4Mux_h I__10339 (
            .O(N__46316),
            .I(N__46302));
    LocalMux I__10338 (
            .O(N__46313),
            .I(N__46297));
    LocalMux I__10337 (
            .O(N__46308),
            .I(N__46297));
    LocalMux I__10336 (
            .O(N__46305),
            .I(N__46289));
    Span4Mux_h I__10335 (
            .O(N__46302),
            .I(N__46286));
    Span4Mux_h I__10334 (
            .O(N__46297),
            .I(N__46283));
    InMux I__10333 (
            .O(N__46296),
            .I(N__46272));
    InMux I__10332 (
            .O(N__46295),
            .I(N__46272));
    InMux I__10331 (
            .O(N__46294),
            .I(N__46272));
    InMux I__10330 (
            .O(N__46293),
            .I(N__46272));
    InMux I__10329 (
            .O(N__46292),
            .I(N__46272));
    Odrv4 I__10328 (
            .O(N__46289),
            .I(N_278));
    Odrv4 I__10327 (
            .O(N__46286),
            .I(N_278));
    Odrv4 I__10326 (
            .O(N__46283),
            .I(N_278));
    LocalMux I__10325 (
            .O(N__46272),
            .I(N_278));
    CEMux I__10324 (
            .O(N__46263),
            .I(N__46260));
    LocalMux I__10323 (
            .O(N__46260),
            .I(N__46257));
    Span4Mux_v I__10322 (
            .O(N__46257),
            .I(N__46254));
    Odrv4 I__10321 (
            .O(N__46254),
            .I(sDAC_mem_41_1_sqmuxa));
    CascadeMux I__10320 (
            .O(N__46251),
            .I(N__46240));
    InMux I__10319 (
            .O(N__46250),
            .I(N__46237));
    InMux I__10318 (
            .O(N__46249),
            .I(N__46234));
    InMux I__10317 (
            .O(N__46248),
            .I(N__46231));
    CascadeMux I__10316 (
            .O(N__46247),
            .I(N__46228));
    CascadeMux I__10315 (
            .O(N__46246),
            .I(N__46225));
    CascadeMux I__10314 (
            .O(N__46245),
            .I(N__46222));
    InMux I__10313 (
            .O(N__46244),
            .I(N__46217));
    InMux I__10312 (
            .O(N__46243),
            .I(N__46217));
    InMux I__10311 (
            .O(N__46240),
            .I(N__46214));
    LocalMux I__10310 (
            .O(N__46237),
            .I(N__46211));
    LocalMux I__10309 (
            .O(N__46234),
            .I(N__46208));
    LocalMux I__10308 (
            .O(N__46231),
            .I(N__46204));
    InMux I__10307 (
            .O(N__46228),
            .I(N__46201));
    InMux I__10306 (
            .O(N__46225),
            .I(N__46196));
    InMux I__10305 (
            .O(N__46222),
            .I(N__46196));
    LocalMux I__10304 (
            .O(N__46217),
            .I(N__46193));
    LocalMux I__10303 (
            .O(N__46214),
            .I(N__46190));
    Span4Mux_h I__10302 (
            .O(N__46211),
            .I(N__46185));
    Span4Mux_h I__10301 (
            .O(N__46208),
            .I(N__46185));
    CascadeMux I__10300 (
            .O(N__46207),
            .I(N__46181));
    Span4Mux_h I__10299 (
            .O(N__46204),
            .I(N__46176));
    LocalMux I__10298 (
            .O(N__46201),
            .I(N__46176));
    LocalMux I__10297 (
            .O(N__46196),
            .I(N__46173));
    Span4Mux_h I__10296 (
            .O(N__46193),
            .I(N__46170));
    Span4Mux_v I__10295 (
            .O(N__46190),
            .I(N__46165));
    Span4Mux_v I__10294 (
            .O(N__46185),
            .I(N__46165));
    InMux I__10293 (
            .O(N__46184),
            .I(N__46160));
    InMux I__10292 (
            .O(N__46181),
            .I(N__46160));
    Span4Mux_v I__10291 (
            .O(N__46176),
            .I(N__46157));
    Span4Mux_v I__10290 (
            .O(N__46173),
            .I(N__46154));
    Span4Mux_h I__10289 (
            .O(N__46170),
            .I(N__46151));
    Span4Mux_h I__10288 (
            .O(N__46165),
            .I(N__46148));
    LocalMux I__10287 (
            .O(N__46160),
            .I(N__46141));
    Span4Mux_h I__10286 (
            .O(N__46157),
            .I(N__46141));
    Span4Mux_v I__10285 (
            .O(N__46154),
            .I(N__46141));
    Odrv4 I__10284 (
            .O(N__46151),
            .I(N_285));
    Odrv4 I__10283 (
            .O(N__46148),
            .I(N_285));
    Odrv4 I__10282 (
            .O(N__46141),
            .I(N_285));
    InMux I__10281 (
            .O(N__46134),
            .I(N__46129));
    CascadeMux I__10280 (
            .O(N__46133),
            .I(N__46125));
    InMux I__10279 (
            .O(N__46132),
            .I(N__46120));
    LocalMux I__10278 (
            .O(N__46129),
            .I(N__46115));
    InMux I__10277 (
            .O(N__46128),
            .I(N__46112));
    InMux I__10276 (
            .O(N__46125),
            .I(N__46105));
    InMux I__10275 (
            .O(N__46124),
            .I(N__46105));
    InMux I__10274 (
            .O(N__46123),
            .I(N__46105));
    LocalMux I__10273 (
            .O(N__46120),
            .I(N__46102));
    InMux I__10272 (
            .O(N__46119),
            .I(N__46097));
    InMux I__10271 (
            .O(N__46118),
            .I(N__46097));
    Span4Mux_h I__10270 (
            .O(N__46115),
            .I(N__46093));
    LocalMux I__10269 (
            .O(N__46112),
            .I(N__46088));
    LocalMux I__10268 (
            .O(N__46105),
            .I(N__46088));
    Span4Mux_v I__10267 (
            .O(N__46102),
            .I(N__46085));
    LocalMux I__10266 (
            .O(N__46097),
            .I(N__46082));
    InMux I__10265 (
            .O(N__46096),
            .I(N__46079));
    Span4Mux_v I__10264 (
            .O(N__46093),
            .I(N__46074));
    Span4Mux_v I__10263 (
            .O(N__46088),
            .I(N__46074));
    Span4Mux_v I__10262 (
            .O(N__46085),
            .I(N__46069));
    Span4Mux_h I__10261 (
            .O(N__46082),
            .I(N__46069));
    LocalMux I__10260 (
            .O(N__46079),
            .I(N__46062));
    Span4Mux_h I__10259 (
            .O(N__46074),
            .I(N__46062));
    Span4Mux_h I__10258 (
            .O(N__46069),
            .I(N__46059));
    InMux I__10257 (
            .O(N__46068),
            .I(N__46056));
    InMux I__10256 (
            .O(N__46067),
            .I(N__46053));
    Odrv4 I__10255 (
            .O(N__46062),
            .I(N_1480));
    Odrv4 I__10254 (
            .O(N__46059),
            .I(N_1480));
    LocalMux I__10253 (
            .O(N__46056),
            .I(N_1480));
    LocalMux I__10252 (
            .O(N__46053),
            .I(N_1480));
    InMux I__10251 (
            .O(N__46044),
            .I(N__46040));
    InMux I__10250 (
            .O(N__46043),
            .I(N__46037));
    LocalMux I__10249 (
            .O(N__46040),
            .I(N__46034));
    LocalMux I__10248 (
            .O(N__46037),
            .I(N__46031));
    Span4Mux_v I__10247 (
            .O(N__46034),
            .I(N__46028));
    Span4Mux_h I__10246 (
            .O(N__46031),
            .I(N__46025));
    Span4Mux_h I__10245 (
            .O(N__46028),
            .I(N__46020));
    Span4Mux_h I__10244 (
            .O(N__46025),
            .I(N__46020));
    Odrv4 I__10243 (
            .O(N__46020),
            .I(N_360));
    InMux I__10242 (
            .O(N__46017),
            .I(N__46014));
    LocalMux I__10241 (
            .O(N__46014),
            .I(N__46011));
    Span4Mux_v I__10240 (
            .O(N__46011),
            .I(N__46008));
    Span4Mux_h I__10239 (
            .O(N__46008),
            .I(N__46005));
    Odrv4 I__10238 (
            .O(N__46005),
            .I(sEEDACZ0Z_0));
    InMux I__10237 (
            .O(N__46002),
            .I(N__45999));
    LocalMux I__10236 (
            .O(N__45999),
            .I(N__45996));
    Span4Mux_v I__10235 (
            .O(N__45996),
            .I(N__45993));
    Odrv4 I__10234 (
            .O(N__45993),
            .I(sEEDACZ0Z_1));
    InMux I__10233 (
            .O(N__45990),
            .I(N__45987));
    LocalMux I__10232 (
            .O(N__45987),
            .I(N__45984));
    Span4Mux_h I__10231 (
            .O(N__45984),
            .I(N__45981));
    Span4Mux_h I__10230 (
            .O(N__45981),
            .I(N__45978));
    Odrv4 I__10229 (
            .O(N__45978),
            .I(sEEDACZ0Z_2));
    InMux I__10228 (
            .O(N__45975),
            .I(N__45972));
    LocalMux I__10227 (
            .O(N__45972),
            .I(N__45969));
    Span4Mux_v I__10226 (
            .O(N__45969),
            .I(N__45966));
    Sp12to4 I__10225 (
            .O(N__45966),
            .I(N__45963));
    Odrv12 I__10224 (
            .O(N__45963),
            .I(sEEDACZ0Z_3));
    InMux I__10223 (
            .O(N__45960),
            .I(N__45957));
    LocalMux I__10222 (
            .O(N__45957),
            .I(N__45954));
    Span4Mux_h I__10221 (
            .O(N__45954),
            .I(N__45951));
    Span4Mux_h I__10220 (
            .O(N__45951),
            .I(N__45948));
    Odrv4 I__10219 (
            .O(N__45948),
            .I(sEEDACZ0Z_4));
    CascadeMux I__10218 (
            .O(N__45945),
            .I(N__45939));
    CascadeMux I__10217 (
            .O(N__45944),
            .I(N__45935));
    InMux I__10216 (
            .O(N__45943),
            .I(N__45922));
    InMux I__10215 (
            .O(N__45942),
            .I(N__45922));
    InMux I__10214 (
            .O(N__45939),
            .I(N__45922));
    InMux I__10213 (
            .O(N__45938),
            .I(N__45922));
    InMux I__10212 (
            .O(N__45935),
            .I(N__45919));
    InMux I__10211 (
            .O(N__45934),
            .I(N__45912));
    InMux I__10210 (
            .O(N__45933),
            .I(N__45912));
    InMux I__10209 (
            .O(N__45932),
            .I(N__45912));
    InMux I__10208 (
            .O(N__45931),
            .I(N__45905));
    LocalMux I__10207 (
            .O(N__45922),
            .I(N__45902));
    LocalMux I__10206 (
            .O(N__45919),
            .I(N__45897));
    LocalMux I__10205 (
            .O(N__45912),
            .I(N__45897));
    InMux I__10204 (
            .O(N__45911),
            .I(N__45892));
    InMux I__10203 (
            .O(N__45910),
            .I(N__45892));
    CascadeMux I__10202 (
            .O(N__45909),
            .I(N__45884));
    CascadeMux I__10201 (
            .O(N__45908),
            .I(N__45862));
    LocalMux I__10200 (
            .O(N__45905),
            .I(N__45856));
    Span4Mux_h I__10199 (
            .O(N__45902),
            .I(N__45849));
    Span4Mux_v I__10198 (
            .O(N__45897),
            .I(N__45849));
    LocalMux I__10197 (
            .O(N__45892),
            .I(N__45849));
    InMux I__10196 (
            .O(N__45891),
            .I(N__45842));
    InMux I__10195 (
            .O(N__45890),
            .I(N__45842));
    InMux I__10194 (
            .O(N__45889),
            .I(N__45838));
    InMux I__10193 (
            .O(N__45888),
            .I(N__45829));
    InMux I__10192 (
            .O(N__45887),
            .I(N__45829));
    InMux I__10191 (
            .O(N__45884),
            .I(N__45829));
    InMux I__10190 (
            .O(N__45883),
            .I(N__45829));
    CascadeMux I__10189 (
            .O(N__45882),
            .I(N__45825));
    InMux I__10188 (
            .O(N__45881),
            .I(N__45822));
    InMux I__10187 (
            .O(N__45880),
            .I(N__45817));
    InMux I__10186 (
            .O(N__45879),
            .I(N__45817));
    InMux I__10185 (
            .O(N__45878),
            .I(N__45814));
    InMux I__10184 (
            .O(N__45877),
            .I(N__45809));
    InMux I__10183 (
            .O(N__45876),
            .I(N__45809));
    CascadeMux I__10182 (
            .O(N__45875),
            .I(N__45804));
    InMux I__10181 (
            .O(N__45874),
            .I(N__45800));
    InMux I__10180 (
            .O(N__45873),
            .I(N__45796));
    InMux I__10179 (
            .O(N__45872),
            .I(N__45793));
    InMux I__10178 (
            .O(N__45871),
            .I(N__45784));
    InMux I__10177 (
            .O(N__45870),
            .I(N__45784));
    InMux I__10176 (
            .O(N__45869),
            .I(N__45784));
    InMux I__10175 (
            .O(N__45868),
            .I(N__45784));
    InMux I__10174 (
            .O(N__45867),
            .I(N__45780));
    InMux I__10173 (
            .O(N__45866),
            .I(N__45777));
    InMux I__10172 (
            .O(N__45865),
            .I(N__45770));
    InMux I__10171 (
            .O(N__45862),
            .I(N__45770));
    InMux I__10170 (
            .O(N__45861),
            .I(N__45770));
    InMux I__10169 (
            .O(N__45860),
            .I(N__45765));
    InMux I__10168 (
            .O(N__45859),
            .I(N__45765));
    Span4Mux_v I__10167 (
            .O(N__45856),
            .I(N__45760));
    Span4Mux_v I__10166 (
            .O(N__45849),
            .I(N__45760));
    InMux I__10165 (
            .O(N__45848),
            .I(N__45755));
    InMux I__10164 (
            .O(N__45847),
            .I(N__45755));
    LocalMux I__10163 (
            .O(N__45842),
            .I(N__45752));
    CascadeMux I__10162 (
            .O(N__45841),
            .I(N__45747));
    LocalMux I__10161 (
            .O(N__45838),
            .I(N__45741));
    LocalMux I__10160 (
            .O(N__45829),
            .I(N__45741));
    InMux I__10159 (
            .O(N__45828),
            .I(N__45738));
    InMux I__10158 (
            .O(N__45825),
            .I(N__45731));
    LocalMux I__10157 (
            .O(N__45822),
            .I(N__45723));
    LocalMux I__10156 (
            .O(N__45817),
            .I(N__45723));
    LocalMux I__10155 (
            .O(N__45814),
            .I(N__45718));
    LocalMux I__10154 (
            .O(N__45809),
            .I(N__45718));
    CascadeMux I__10153 (
            .O(N__45808),
            .I(N__45713));
    CascadeMux I__10152 (
            .O(N__45807),
            .I(N__45706));
    InMux I__10151 (
            .O(N__45804),
            .I(N__45701));
    InMux I__10150 (
            .O(N__45803),
            .I(N__45701));
    LocalMux I__10149 (
            .O(N__45800),
            .I(N__45698));
    InMux I__10148 (
            .O(N__45799),
            .I(N__45695));
    LocalMux I__10147 (
            .O(N__45796),
            .I(N__45690));
    LocalMux I__10146 (
            .O(N__45793),
            .I(N__45690));
    LocalMux I__10145 (
            .O(N__45784),
            .I(N__45687));
    InMux I__10144 (
            .O(N__45783),
            .I(N__45684));
    LocalMux I__10143 (
            .O(N__45780),
            .I(N__45681));
    LocalMux I__10142 (
            .O(N__45777),
            .I(N__45676));
    LocalMux I__10141 (
            .O(N__45770),
            .I(N__45676));
    LocalMux I__10140 (
            .O(N__45765),
            .I(N__45667));
    Span4Mux_h I__10139 (
            .O(N__45760),
            .I(N__45667));
    LocalMux I__10138 (
            .O(N__45755),
            .I(N__45667));
    Span4Mux_h I__10137 (
            .O(N__45752),
            .I(N__45667));
    InMux I__10136 (
            .O(N__45751),
            .I(N__45664));
    InMux I__10135 (
            .O(N__45750),
            .I(N__45661));
    InMux I__10134 (
            .O(N__45747),
            .I(N__45656));
    InMux I__10133 (
            .O(N__45746),
            .I(N__45656));
    Span4Mux_h I__10132 (
            .O(N__45741),
            .I(N__45651));
    LocalMux I__10131 (
            .O(N__45738),
            .I(N__45651));
    InMux I__10130 (
            .O(N__45737),
            .I(N__45648));
    InMux I__10129 (
            .O(N__45736),
            .I(N__45645));
    InMux I__10128 (
            .O(N__45735),
            .I(N__45640));
    InMux I__10127 (
            .O(N__45734),
            .I(N__45640));
    LocalMux I__10126 (
            .O(N__45731),
            .I(N__45636));
    InMux I__10125 (
            .O(N__45730),
            .I(N__45629));
    InMux I__10124 (
            .O(N__45729),
            .I(N__45629));
    InMux I__10123 (
            .O(N__45728),
            .I(N__45629));
    Span4Mux_h I__10122 (
            .O(N__45723),
            .I(N__45624));
    Span4Mux_v I__10121 (
            .O(N__45718),
            .I(N__45624));
    InMux I__10120 (
            .O(N__45717),
            .I(N__45621));
    InMux I__10119 (
            .O(N__45716),
            .I(N__45618));
    InMux I__10118 (
            .O(N__45713),
            .I(N__45611));
    InMux I__10117 (
            .O(N__45712),
            .I(N__45611));
    InMux I__10116 (
            .O(N__45711),
            .I(N__45611));
    InMux I__10115 (
            .O(N__45710),
            .I(N__45606));
    InMux I__10114 (
            .O(N__45709),
            .I(N__45606));
    InMux I__10113 (
            .O(N__45706),
            .I(N__45603));
    LocalMux I__10112 (
            .O(N__45701),
            .I(N__45596));
    Span4Mux_h I__10111 (
            .O(N__45698),
            .I(N__45596));
    LocalMux I__10110 (
            .O(N__45695),
            .I(N__45596));
    Span4Mux_h I__10109 (
            .O(N__45690),
            .I(N__45591));
    Span4Mux_v I__10108 (
            .O(N__45687),
            .I(N__45591));
    LocalMux I__10107 (
            .O(N__45684),
            .I(N__45582));
    Span4Mux_h I__10106 (
            .O(N__45681),
            .I(N__45582));
    Span4Mux_h I__10105 (
            .O(N__45676),
            .I(N__45582));
    Span4Mux_v I__10104 (
            .O(N__45667),
            .I(N__45582));
    LocalMux I__10103 (
            .O(N__45664),
            .I(N__45567));
    LocalMux I__10102 (
            .O(N__45661),
            .I(N__45567));
    LocalMux I__10101 (
            .O(N__45656),
            .I(N__45567));
    Sp12to4 I__10100 (
            .O(N__45651),
            .I(N__45567));
    LocalMux I__10099 (
            .O(N__45648),
            .I(N__45567));
    LocalMux I__10098 (
            .O(N__45645),
            .I(N__45567));
    LocalMux I__10097 (
            .O(N__45640),
            .I(N__45567));
    InMux I__10096 (
            .O(N__45639),
            .I(N__45564));
    Span4Mux_h I__10095 (
            .O(N__45636),
            .I(N__45557));
    LocalMux I__10094 (
            .O(N__45629),
            .I(N__45557));
    Span4Mux_v I__10093 (
            .O(N__45624),
            .I(N__45557));
    LocalMux I__10092 (
            .O(N__45621),
            .I(sDAC_mem_pointerZ0Z_2));
    LocalMux I__10091 (
            .O(N__45618),
            .I(sDAC_mem_pointerZ0Z_2));
    LocalMux I__10090 (
            .O(N__45611),
            .I(sDAC_mem_pointerZ0Z_2));
    LocalMux I__10089 (
            .O(N__45606),
            .I(sDAC_mem_pointerZ0Z_2));
    LocalMux I__10088 (
            .O(N__45603),
            .I(sDAC_mem_pointerZ0Z_2));
    Odrv4 I__10087 (
            .O(N__45596),
            .I(sDAC_mem_pointerZ0Z_2));
    Odrv4 I__10086 (
            .O(N__45591),
            .I(sDAC_mem_pointerZ0Z_2));
    Odrv4 I__10085 (
            .O(N__45582),
            .I(sDAC_mem_pointerZ0Z_2));
    Odrv12 I__10084 (
            .O(N__45567),
            .I(sDAC_mem_pointerZ0Z_2));
    LocalMux I__10083 (
            .O(N__45564),
            .I(sDAC_mem_pointerZ0Z_2));
    Odrv4 I__10082 (
            .O(N__45557),
            .I(sDAC_mem_pointerZ0Z_2));
    CascadeMux I__10081 (
            .O(N__45534),
            .I(N__45530));
    InMux I__10080 (
            .O(N__45533),
            .I(N__45515));
    InMux I__10079 (
            .O(N__45530),
            .I(N__45512));
    InMux I__10078 (
            .O(N__45529),
            .I(N__45507));
    InMux I__10077 (
            .O(N__45528),
            .I(N__45507));
    InMux I__10076 (
            .O(N__45527),
            .I(N__45502));
    InMux I__10075 (
            .O(N__45526),
            .I(N__45502));
    InMux I__10074 (
            .O(N__45525),
            .I(N__45496));
    InMux I__10073 (
            .O(N__45524),
            .I(N__45496));
    InMux I__10072 (
            .O(N__45523),
            .I(N__45487));
    InMux I__10071 (
            .O(N__45522),
            .I(N__45482));
    InMux I__10070 (
            .O(N__45521),
            .I(N__45482));
    InMux I__10069 (
            .O(N__45520),
            .I(N__45477));
    InMux I__10068 (
            .O(N__45519),
            .I(N__45472));
    InMux I__10067 (
            .O(N__45518),
            .I(N__45472));
    LocalMux I__10066 (
            .O(N__45515),
            .I(N__45465));
    LocalMux I__10065 (
            .O(N__45512),
            .I(N__45465));
    LocalMux I__10064 (
            .O(N__45507),
            .I(N__45465));
    LocalMux I__10063 (
            .O(N__45502),
            .I(N__45462));
    InMux I__10062 (
            .O(N__45501),
            .I(N__45459));
    LocalMux I__10061 (
            .O(N__45496),
            .I(N__45454));
    InMux I__10060 (
            .O(N__45495),
            .I(N__45449));
    InMux I__10059 (
            .O(N__45494),
            .I(N__45449));
    InMux I__10058 (
            .O(N__45493),
            .I(N__45444));
    InMux I__10057 (
            .O(N__45492),
            .I(N__45444));
    CascadeMux I__10056 (
            .O(N__45491),
            .I(N__45441));
    InMux I__10055 (
            .O(N__45490),
            .I(N__45436));
    LocalMux I__10054 (
            .O(N__45487),
            .I(N__45433));
    LocalMux I__10053 (
            .O(N__45482),
            .I(N__45430));
    InMux I__10052 (
            .O(N__45481),
            .I(N__45425));
    InMux I__10051 (
            .O(N__45480),
            .I(N__45425));
    LocalMux I__10050 (
            .O(N__45477),
            .I(N__45416));
    LocalMux I__10049 (
            .O(N__45472),
            .I(N__45416));
    Span4Mux_v I__10048 (
            .O(N__45465),
            .I(N__45411));
    Span4Mux_v I__10047 (
            .O(N__45462),
            .I(N__45406));
    LocalMux I__10046 (
            .O(N__45459),
            .I(N__45406));
    InMux I__10045 (
            .O(N__45458),
            .I(N__45401));
    InMux I__10044 (
            .O(N__45457),
            .I(N__45401));
    Span4Mux_v I__10043 (
            .O(N__45454),
            .I(N__45396));
    LocalMux I__10042 (
            .O(N__45449),
            .I(N__45396));
    LocalMux I__10041 (
            .O(N__45444),
            .I(N__45393));
    InMux I__10040 (
            .O(N__45441),
            .I(N__45390));
    InMux I__10039 (
            .O(N__45440),
            .I(N__45387));
    InMux I__10038 (
            .O(N__45439),
            .I(N__45384));
    LocalMux I__10037 (
            .O(N__45436),
            .I(N__45381));
    Span4Mux_v I__10036 (
            .O(N__45433),
            .I(N__45374));
    Span4Mux_h I__10035 (
            .O(N__45430),
            .I(N__45374));
    LocalMux I__10034 (
            .O(N__45425),
            .I(N__45374));
    InMux I__10033 (
            .O(N__45424),
            .I(N__45369));
    InMux I__10032 (
            .O(N__45423),
            .I(N__45366));
    InMux I__10031 (
            .O(N__45422),
            .I(N__45361));
    InMux I__10030 (
            .O(N__45421),
            .I(N__45361));
    Span4Mux_v I__10029 (
            .O(N__45416),
            .I(N__45358));
    InMux I__10028 (
            .O(N__45415),
            .I(N__45353));
    InMux I__10027 (
            .O(N__45414),
            .I(N__45353));
    Span4Mux_h I__10026 (
            .O(N__45411),
            .I(N__45348));
    Span4Mux_v I__10025 (
            .O(N__45406),
            .I(N__45348));
    LocalMux I__10024 (
            .O(N__45401),
            .I(N__45341));
    Span4Mux_v I__10023 (
            .O(N__45396),
            .I(N__45341));
    Span4Mux_v I__10022 (
            .O(N__45393),
            .I(N__45341));
    LocalMux I__10021 (
            .O(N__45390),
            .I(N__45334));
    LocalMux I__10020 (
            .O(N__45387),
            .I(N__45334));
    LocalMux I__10019 (
            .O(N__45384),
            .I(N__45334));
    Span4Mux_v I__10018 (
            .O(N__45381),
            .I(N__45329));
    Span4Mux_v I__10017 (
            .O(N__45374),
            .I(N__45329));
    InMux I__10016 (
            .O(N__45373),
            .I(N__45324));
    InMux I__10015 (
            .O(N__45372),
            .I(N__45324));
    LocalMux I__10014 (
            .O(N__45369),
            .I(sDAC_mem_pointerZ0Z_1));
    LocalMux I__10013 (
            .O(N__45366),
            .I(sDAC_mem_pointerZ0Z_1));
    LocalMux I__10012 (
            .O(N__45361),
            .I(sDAC_mem_pointerZ0Z_1));
    Odrv4 I__10011 (
            .O(N__45358),
            .I(sDAC_mem_pointerZ0Z_1));
    LocalMux I__10010 (
            .O(N__45353),
            .I(sDAC_mem_pointerZ0Z_1));
    Odrv4 I__10009 (
            .O(N__45348),
            .I(sDAC_mem_pointerZ0Z_1));
    Odrv4 I__10008 (
            .O(N__45341),
            .I(sDAC_mem_pointerZ0Z_1));
    Odrv12 I__10007 (
            .O(N__45334),
            .I(sDAC_mem_pointerZ0Z_1));
    Odrv4 I__10006 (
            .O(N__45329),
            .I(sDAC_mem_pointerZ0Z_1));
    LocalMux I__10005 (
            .O(N__45324),
            .I(sDAC_mem_pointerZ0Z_1));
    CascadeMux I__10004 (
            .O(N__45303),
            .I(sDAC_data_RNO_18Z0Z_4_cascade_));
    InMux I__10003 (
            .O(N__45300),
            .I(N__45297));
    LocalMux I__10002 (
            .O(N__45297),
            .I(sDAC_data_2_24_ns_1_4));
    InMux I__10001 (
            .O(N__45294),
            .I(N__45291));
    LocalMux I__10000 (
            .O(N__45291),
            .I(sDAC_mem_12Z0Z_0));
    InMux I__9999 (
            .O(N__45288),
            .I(N__45285));
    LocalMux I__9998 (
            .O(N__45285),
            .I(N__45282));
    Odrv4 I__9997 (
            .O(N__45282),
            .I(sDAC_mem_15Z0Z_1));
    InMux I__9996 (
            .O(N__45279),
            .I(N__45276));
    LocalMux I__9995 (
            .O(N__45276),
            .I(sDAC_mem_14Z0Z_1));
    InMux I__9994 (
            .O(N__45273),
            .I(N__45270));
    LocalMux I__9993 (
            .O(N__45270),
            .I(sDAC_data_RNO_19Z0Z_4));
    InMux I__9992 (
            .O(N__45267),
            .I(N__45264));
    LocalMux I__9991 (
            .O(N__45264),
            .I(sDAC_mem_12Z0Z_1));
    InMux I__9990 (
            .O(N__45261),
            .I(N__45258));
    LocalMux I__9989 (
            .O(N__45258),
            .I(N__45255));
    Span4Mux_v I__9988 (
            .O(N__45255),
            .I(N__45252));
    Span4Mux_h I__9987 (
            .O(N__45252),
            .I(N__45249));
    Odrv4 I__9986 (
            .O(N__45249),
            .I(sDAC_mem_27Z0Z_0));
    CEMux I__9985 (
            .O(N__45246),
            .I(N__45242));
    CEMux I__9984 (
            .O(N__45245),
            .I(N__45239));
    LocalMux I__9983 (
            .O(N__45242),
            .I(sDAC_mem_27_1_sqmuxa));
    LocalMux I__9982 (
            .O(N__45239),
            .I(sDAC_mem_27_1_sqmuxa));
    InMux I__9981 (
            .O(N__45234),
            .I(N__45231));
    LocalMux I__9980 (
            .O(N__45231),
            .I(N__45228));
    Odrv12 I__9979 (
            .O(N__45228),
            .I(sDAC_mem_13Z0Z_6));
    InMux I__9978 (
            .O(N__45225),
            .I(N__45222));
    LocalMux I__9977 (
            .O(N__45222),
            .I(sDAC_mem_13Z0Z_5));
    InMux I__9976 (
            .O(N__45219),
            .I(N__45216));
    LocalMux I__9975 (
            .O(N__45216),
            .I(N__45213));
    Span4Mux_h I__9974 (
            .O(N__45213),
            .I(N__45210));
    Odrv4 I__9973 (
            .O(N__45210),
            .I(sDAC_mem_16Z0Z_1));
    InMux I__9972 (
            .O(N__45207),
            .I(N__45204));
    LocalMux I__9971 (
            .O(N__45204),
            .I(N__45201));
    Span4Mux_v I__9970 (
            .O(N__45201),
            .I(N__45198));
    Span4Mux_h I__9969 (
            .O(N__45198),
            .I(N__45195));
    Odrv4 I__9968 (
            .O(N__45195),
            .I(sDAC_mem_11Z0Z_2));
    InMux I__9967 (
            .O(N__45192),
            .I(N__45189));
    LocalMux I__9966 (
            .O(N__45189),
            .I(N__45186));
    Span4Mux_v I__9965 (
            .O(N__45186),
            .I(N__45183));
    Odrv4 I__9964 (
            .O(N__45183),
            .I(sDAC_mem_11Z0Z_3));
    InMux I__9963 (
            .O(N__45180),
            .I(N__45177));
    LocalMux I__9962 (
            .O(N__45177),
            .I(N__45174));
    Span4Mux_h I__9961 (
            .O(N__45174),
            .I(N__45171));
    Span4Mux_v I__9960 (
            .O(N__45171),
            .I(N__45168));
    Odrv4 I__9959 (
            .O(N__45168),
            .I(sDAC_mem_11Z0Z_4));
    InMux I__9958 (
            .O(N__45165),
            .I(N__45162));
    LocalMux I__9957 (
            .O(N__45162),
            .I(N__45159));
    Odrv4 I__9956 (
            .O(N__45159),
            .I(sDAC_mem_11Z0Z_5));
    InMux I__9955 (
            .O(N__45156),
            .I(N__45153));
    LocalMux I__9954 (
            .O(N__45153),
            .I(N__45150));
    Span4Mux_h I__9953 (
            .O(N__45150),
            .I(N__45147));
    Span4Mux_v I__9952 (
            .O(N__45147),
            .I(N__45144));
    Odrv4 I__9951 (
            .O(N__45144),
            .I(sDAC_mem_11Z0Z_6));
    InMux I__9950 (
            .O(N__45141),
            .I(N__45138));
    LocalMux I__9949 (
            .O(N__45138),
            .I(N__45135));
    Span4Mux_v I__9948 (
            .O(N__45135),
            .I(N__45132));
    Odrv4 I__9947 (
            .O(N__45132),
            .I(sDAC_mem_11Z0Z_7));
    CEMux I__9946 (
            .O(N__45129),
            .I(N__45126));
    LocalMux I__9945 (
            .O(N__45126),
            .I(sDAC_mem_11_1_sqmuxa));
    InMux I__9944 (
            .O(N__45123),
            .I(N__45120));
    LocalMux I__9943 (
            .O(N__45120),
            .I(N__45117));
    Odrv12 I__9942 (
            .O(N__45117),
            .I(sDAC_mem_15Z0Z_0));
    InMux I__9941 (
            .O(N__45114),
            .I(N__45111));
    LocalMux I__9940 (
            .O(N__45111),
            .I(sDAC_mem_14Z0Z_0));
    CascadeMux I__9939 (
            .O(N__45108),
            .I(sDAC_data_RNO_18Z0Z_3_cascade_));
    InMux I__9938 (
            .O(N__45105),
            .I(N__45102));
    LocalMux I__9937 (
            .O(N__45102),
            .I(sDAC_data_RNO_19Z0Z_3));
    InMux I__9936 (
            .O(N__45099),
            .I(N__45096));
    LocalMux I__9935 (
            .O(N__45096),
            .I(N__45093));
    Odrv4 I__9934 (
            .O(N__45093),
            .I(sDAC_data_2_24_ns_1_3));
    InMux I__9933 (
            .O(N__45090),
            .I(N__45087));
    LocalMux I__9932 (
            .O(N__45087),
            .I(N__45084));
    Span4Mux_v I__9931 (
            .O(N__45084),
            .I(N__45081));
    Span4Mux_h I__9930 (
            .O(N__45081),
            .I(N__45078));
    Odrv4 I__9929 (
            .O(N__45078),
            .I(sDAC_mem_15Z0Z_2));
    InMux I__9928 (
            .O(N__45075),
            .I(N__45072));
    LocalMux I__9927 (
            .O(N__45072),
            .I(N__45069));
    Span4Mux_v I__9926 (
            .O(N__45069),
            .I(N__45066));
    Span4Mux_h I__9925 (
            .O(N__45066),
            .I(N__45063));
    Odrv4 I__9924 (
            .O(N__45063),
            .I(sDAC_mem_15Z0Z_3));
    InMux I__9923 (
            .O(N__45060),
            .I(N__45057));
    LocalMux I__9922 (
            .O(N__45057),
            .I(N__45054));
    Span4Mux_v I__9921 (
            .O(N__45054),
            .I(N__45051));
    Odrv4 I__9920 (
            .O(N__45051),
            .I(sDAC_mem_15Z0Z_4));
    InMux I__9919 (
            .O(N__45048),
            .I(N__45045));
    LocalMux I__9918 (
            .O(N__45045),
            .I(N__45042));
    Span4Mux_v I__9917 (
            .O(N__45042),
            .I(N__45039));
    Odrv4 I__9916 (
            .O(N__45039),
            .I(sDAC_mem_15Z0Z_5));
    InMux I__9915 (
            .O(N__45036),
            .I(N__45033));
    LocalMux I__9914 (
            .O(N__45033),
            .I(N__45030));
    Span4Mux_v I__9913 (
            .O(N__45030),
            .I(N__45027));
    Odrv4 I__9912 (
            .O(N__45027),
            .I(sDAC_mem_15Z0Z_6));
    CEMux I__9911 (
            .O(N__45024),
            .I(N__45021));
    LocalMux I__9910 (
            .O(N__45021),
            .I(N__45018));
    Span4Mux_h I__9909 (
            .O(N__45018),
            .I(N__45015));
    Odrv4 I__9908 (
            .O(N__45015),
            .I(sDAC_mem_15_1_sqmuxa));
    InMux I__9907 (
            .O(N__45012),
            .I(N__45009));
    LocalMux I__9906 (
            .O(N__45009),
            .I(sDAC_mem_11Z0Z_0));
    InMux I__9905 (
            .O(N__45006),
            .I(N__45003));
    LocalMux I__9904 (
            .O(N__45003),
            .I(sDAC_mem_11Z0Z_1));
    CEMux I__9903 (
            .O(N__45000),
            .I(N__44997));
    LocalMux I__9902 (
            .O(N__44997),
            .I(N__44994));
    Span4Mux_h I__9901 (
            .O(N__44994),
            .I(N__44990));
    CEMux I__9900 (
            .O(N__44993),
            .I(N__44987));
    Span4Mux_h I__9899 (
            .O(N__44990),
            .I(N__44984));
    LocalMux I__9898 (
            .O(N__44987),
            .I(N__44981));
    Odrv4 I__9897 (
            .O(N__44984),
            .I(sDAC_mem_10_1_sqmuxa));
    Odrv12 I__9896 (
            .O(N__44981),
            .I(sDAC_mem_10_1_sqmuxa));
    CEMux I__9895 (
            .O(N__44976),
            .I(N__44973));
    LocalMux I__9894 (
            .O(N__44973),
            .I(N__44970));
    Span4Mux_v I__9893 (
            .O(N__44970),
            .I(N__44967));
    Span4Mux_h I__9892 (
            .O(N__44967),
            .I(N__44964));
    Odrv4 I__9891 (
            .O(N__44964),
            .I(sDAC_mem_42_1_sqmuxa));
    CascadeMux I__9890 (
            .O(N__44961),
            .I(N__44954));
    InMux I__9889 (
            .O(N__44960),
            .I(N__44949));
    InMux I__9888 (
            .O(N__44959),
            .I(N__44946));
    InMux I__9887 (
            .O(N__44958),
            .I(N__44943));
    InMux I__9886 (
            .O(N__44957),
            .I(N__44940));
    InMux I__9885 (
            .O(N__44954),
            .I(N__44935));
    InMux I__9884 (
            .O(N__44953),
            .I(N__44935));
    InMux I__9883 (
            .O(N__44952),
            .I(N__44932));
    LocalMux I__9882 (
            .O(N__44949),
            .I(N__44926));
    LocalMux I__9881 (
            .O(N__44946),
            .I(N__44926));
    LocalMux I__9880 (
            .O(N__44943),
            .I(N__44923));
    LocalMux I__9879 (
            .O(N__44940),
            .I(N__44920));
    LocalMux I__9878 (
            .O(N__44935),
            .I(N__44915));
    LocalMux I__9877 (
            .O(N__44932),
            .I(N__44915));
    InMux I__9876 (
            .O(N__44931),
            .I(N__44912));
    Span4Mux_h I__9875 (
            .O(N__44926),
            .I(N__44909));
    Span4Mux_h I__9874 (
            .O(N__44923),
            .I(N__44906));
    Span4Mux_v I__9873 (
            .O(N__44920),
            .I(N__44901));
    Span4Mux_h I__9872 (
            .O(N__44915),
            .I(N__44901));
    LocalMux I__9871 (
            .O(N__44912),
            .I(N__44898));
    Span4Mux_h I__9870 (
            .O(N__44909),
            .I(N__44893));
    Span4Mux_h I__9869 (
            .O(N__44906),
            .I(N__44890));
    Span4Mux_h I__9868 (
            .O(N__44901),
            .I(N__44885));
    Span4Mux_h I__9867 (
            .O(N__44898),
            .I(N__44885));
    InMux I__9866 (
            .O(N__44897),
            .I(N__44880));
    InMux I__9865 (
            .O(N__44896),
            .I(N__44880));
    Odrv4 I__9864 (
            .O(N__44893),
            .I(sAddressZ0Z_2));
    Odrv4 I__9863 (
            .O(N__44890),
            .I(sAddressZ0Z_2));
    Odrv4 I__9862 (
            .O(N__44885),
            .I(sAddressZ0Z_2));
    LocalMux I__9861 (
            .O(N__44880),
            .I(sAddressZ0Z_2));
    InMux I__9860 (
            .O(N__44871),
            .I(N__44865));
    InMux I__9859 (
            .O(N__44870),
            .I(N__44862));
    InMux I__9858 (
            .O(N__44869),
            .I(N__44859));
    InMux I__9857 (
            .O(N__44868),
            .I(N__44856));
    LocalMux I__9856 (
            .O(N__44865),
            .I(N__44848));
    LocalMux I__9855 (
            .O(N__44862),
            .I(N__44848));
    LocalMux I__9854 (
            .O(N__44859),
            .I(N__44848));
    LocalMux I__9853 (
            .O(N__44856),
            .I(N__44845));
    InMux I__9852 (
            .O(N__44855),
            .I(N__44842));
    Span4Mux_v I__9851 (
            .O(N__44848),
            .I(N__44839));
    Span4Mux_h I__9850 (
            .O(N__44845),
            .I(N__44836));
    LocalMux I__9849 (
            .O(N__44842),
            .I(N__44833));
    Span4Mux_h I__9848 (
            .O(N__44839),
            .I(N__44828));
    Span4Mux_h I__9847 (
            .O(N__44836),
            .I(N__44825));
    Span4Mux_v I__9846 (
            .O(N__44833),
            .I(N__44822));
    InMux I__9845 (
            .O(N__44832),
            .I(N__44817));
    InMux I__9844 (
            .O(N__44831),
            .I(N__44817));
    Odrv4 I__9843 (
            .O(N__44828),
            .I(sAddressZ0Z_1));
    Odrv4 I__9842 (
            .O(N__44825),
            .I(sAddressZ0Z_1));
    Odrv4 I__9841 (
            .O(N__44822),
            .I(sAddressZ0Z_1));
    LocalMux I__9840 (
            .O(N__44817),
            .I(sAddressZ0Z_1));
    CascadeMux I__9839 (
            .O(N__44808),
            .I(N__44804));
    CascadeMux I__9838 (
            .O(N__44807),
            .I(N__44801));
    InMux I__9837 (
            .O(N__44804),
            .I(N__44798));
    InMux I__9836 (
            .O(N__44801),
            .I(N__44794));
    LocalMux I__9835 (
            .O(N__44798),
            .I(N__44791));
    CascadeMux I__9834 (
            .O(N__44797),
            .I(N__44788));
    LocalMux I__9833 (
            .O(N__44794),
            .I(N__44785));
    Span4Mux_h I__9832 (
            .O(N__44791),
            .I(N__44782));
    InMux I__9831 (
            .O(N__44788),
            .I(N__44779));
    Span4Mux_v I__9830 (
            .O(N__44785),
            .I(N__44775));
    Span4Mux_v I__9829 (
            .O(N__44782),
            .I(N__44770));
    LocalMux I__9828 (
            .O(N__44779),
            .I(N__44770));
    InMux I__9827 (
            .O(N__44778),
            .I(N__44767));
    Span4Mux_v I__9826 (
            .O(N__44775),
            .I(N__44762));
    Span4Mux_v I__9825 (
            .O(N__44770),
            .I(N__44762));
    LocalMux I__9824 (
            .O(N__44767),
            .I(N__44759));
    Sp12to4 I__9823 (
            .O(N__44762),
            .I(N__44754));
    Sp12to4 I__9822 (
            .O(N__44759),
            .I(N__44754));
    Odrv12 I__9821 (
            .O(N__44754),
            .I(sDAC_mem_30_1_sqmuxa_0_a2_1_0));
    InMux I__9820 (
            .O(N__44751),
            .I(N__44746));
    InMux I__9819 (
            .O(N__44750),
            .I(N__44742));
    InMux I__9818 (
            .O(N__44749),
            .I(N__44738));
    LocalMux I__9817 (
            .O(N__44746),
            .I(N__44735));
    InMux I__9816 (
            .O(N__44745),
            .I(N__44732));
    LocalMux I__9815 (
            .O(N__44742),
            .I(N__44727));
    InMux I__9814 (
            .O(N__44741),
            .I(N__44724));
    LocalMux I__9813 (
            .O(N__44738),
            .I(N__44719));
    Span4Mux_v I__9812 (
            .O(N__44735),
            .I(N__44711));
    LocalMux I__9811 (
            .O(N__44732),
            .I(N__44711));
    InMux I__9810 (
            .O(N__44731),
            .I(N__44706));
    InMux I__9809 (
            .O(N__44730),
            .I(N__44706));
    Span4Mux_v I__9808 (
            .O(N__44727),
            .I(N__44701));
    LocalMux I__9807 (
            .O(N__44724),
            .I(N__44701));
    InMux I__9806 (
            .O(N__44723),
            .I(N__44698));
    InMux I__9805 (
            .O(N__44722),
            .I(N__44695));
    Span4Mux_h I__9804 (
            .O(N__44719),
            .I(N__44690));
    InMux I__9803 (
            .O(N__44718),
            .I(N__44687));
    InMux I__9802 (
            .O(N__44717),
            .I(N__44682));
    InMux I__9801 (
            .O(N__44716),
            .I(N__44682));
    Span4Mux_h I__9800 (
            .O(N__44711),
            .I(N__44679));
    LocalMux I__9799 (
            .O(N__44706),
            .I(N__44674));
    Span4Mux_h I__9798 (
            .O(N__44701),
            .I(N__44674));
    LocalMux I__9797 (
            .O(N__44698),
            .I(N__44669));
    LocalMux I__9796 (
            .O(N__44695),
            .I(N__44669));
    InMux I__9795 (
            .O(N__44694),
            .I(N__44664));
    InMux I__9794 (
            .O(N__44693),
            .I(N__44664));
    Odrv4 I__9793 (
            .O(N__44690),
            .I(N_275));
    LocalMux I__9792 (
            .O(N__44687),
            .I(N_275));
    LocalMux I__9791 (
            .O(N__44682),
            .I(N_275));
    Odrv4 I__9790 (
            .O(N__44679),
            .I(N_275));
    Odrv4 I__9789 (
            .O(N__44674),
            .I(N_275));
    Odrv12 I__9788 (
            .O(N__44669),
            .I(N_275));
    LocalMux I__9787 (
            .O(N__44664),
            .I(N_275));
    InMux I__9786 (
            .O(N__44649),
            .I(N__44646));
    LocalMux I__9785 (
            .O(N__44646),
            .I(N__44641));
    InMux I__9784 (
            .O(N__44645),
            .I(N__44638));
    InMux I__9783 (
            .O(N__44644),
            .I(N__44633));
    Span4Mux_v I__9782 (
            .O(N__44641),
            .I(N__44628));
    LocalMux I__9781 (
            .O(N__44638),
            .I(N__44628));
    InMux I__9780 (
            .O(N__44637),
            .I(N__44625));
    InMux I__9779 (
            .O(N__44636),
            .I(N__44622));
    LocalMux I__9778 (
            .O(N__44633),
            .I(N__44617));
    Span4Mux_h I__9777 (
            .O(N__44628),
            .I(N__44617));
    LocalMux I__9776 (
            .O(N__44625),
            .I(N__44614));
    LocalMux I__9775 (
            .O(N__44622),
            .I(N__44610));
    Span4Mux_v I__9774 (
            .O(N__44617),
            .I(N__44605));
    Span4Mux_v I__9773 (
            .O(N__44614),
            .I(N__44605));
    InMux I__9772 (
            .O(N__44613),
            .I(N__44602));
    Odrv12 I__9771 (
            .O(N__44610),
            .I(sAddressZ0Z_4));
    Odrv4 I__9770 (
            .O(N__44605),
            .I(sAddressZ0Z_4));
    LocalMux I__9769 (
            .O(N__44602),
            .I(sAddressZ0Z_4));
    CascadeMux I__9768 (
            .O(N__44595),
            .I(N__44589));
    CascadeMux I__9767 (
            .O(N__44594),
            .I(N__44583));
    CascadeMux I__9766 (
            .O(N__44593),
            .I(N__44580));
    InMux I__9765 (
            .O(N__44592),
            .I(N__44577));
    InMux I__9764 (
            .O(N__44589),
            .I(N__44572));
    InMux I__9763 (
            .O(N__44588),
            .I(N__44572));
    CascadeMux I__9762 (
            .O(N__44587),
            .I(N__44568));
    CascadeMux I__9761 (
            .O(N__44586),
            .I(N__44565));
    InMux I__9760 (
            .O(N__44583),
            .I(N__44560));
    InMux I__9759 (
            .O(N__44580),
            .I(N__44560));
    LocalMux I__9758 (
            .O(N__44577),
            .I(N__44555));
    LocalMux I__9757 (
            .O(N__44572),
            .I(N__44555));
    CascadeMux I__9756 (
            .O(N__44571),
            .I(N__44550));
    InMux I__9755 (
            .O(N__44568),
            .I(N__44546));
    InMux I__9754 (
            .O(N__44565),
            .I(N__44543));
    LocalMux I__9753 (
            .O(N__44560),
            .I(N__44540));
    Span4Mux_h I__9752 (
            .O(N__44555),
            .I(N__44536));
    CascadeMux I__9751 (
            .O(N__44554),
            .I(N__44533));
    InMux I__9750 (
            .O(N__44553),
            .I(N__44528));
    InMux I__9749 (
            .O(N__44550),
            .I(N__44528));
    InMux I__9748 (
            .O(N__44549),
            .I(N__44525));
    LocalMux I__9747 (
            .O(N__44546),
            .I(N__44520));
    LocalMux I__9746 (
            .O(N__44543),
            .I(N__44520));
    Span4Mux_h I__9745 (
            .O(N__44540),
            .I(N__44517));
    InMux I__9744 (
            .O(N__44539),
            .I(N__44514));
    Span4Mux_h I__9743 (
            .O(N__44536),
            .I(N__44511));
    InMux I__9742 (
            .O(N__44533),
            .I(N__44508));
    LocalMux I__9741 (
            .O(N__44528),
            .I(N__44503));
    LocalMux I__9740 (
            .O(N__44525),
            .I(N__44503));
    Span4Mux_h I__9739 (
            .O(N__44520),
            .I(N__44500));
    Span4Mux_v I__9738 (
            .O(N__44517),
            .I(N__44497));
    LocalMux I__9737 (
            .O(N__44514),
            .I(N__44492));
    Span4Mux_h I__9736 (
            .O(N__44511),
            .I(N__44492));
    LocalMux I__9735 (
            .O(N__44508),
            .I(N_286));
    Odrv12 I__9734 (
            .O(N__44503),
            .I(N_286));
    Odrv4 I__9733 (
            .O(N__44500),
            .I(N_286));
    Odrv4 I__9732 (
            .O(N__44497),
            .I(N_286));
    Odrv4 I__9731 (
            .O(N__44492),
            .I(N_286));
    CascadeMux I__9730 (
            .O(N__44481),
            .I(N_278_cascade_));
    CascadeMux I__9729 (
            .O(N__44478),
            .I(N__44475));
    InMux I__9728 (
            .O(N__44475),
            .I(N__44472));
    LocalMux I__9727 (
            .O(N__44472),
            .I(N__44466));
    CascadeMux I__9726 (
            .O(N__44471),
            .I(N__44463));
    CascadeMux I__9725 (
            .O(N__44470),
            .I(N__44460));
    CascadeMux I__9724 (
            .O(N__44469),
            .I(N__44456));
    Span4Mux_h I__9723 (
            .O(N__44466),
            .I(N__44453));
    InMux I__9722 (
            .O(N__44463),
            .I(N__44446));
    InMux I__9721 (
            .O(N__44460),
            .I(N__44446));
    InMux I__9720 (
            .O(N__44459),
            .I(N__44446));
    InMux I__9719 (
            .O(N__44456),
            .I(N__44440));
    Span4Mux_v I__9718 (
            .O(N__44453),
            .I(N__44437));
    LocalMux I__9717 (
            .O(N__44446),
            .I(N__44434));
    InMux I__9716 (
            .O(N__44445),
            .I(N__44431));
    InMux I__9715 (
            .O(N__44444),
            .I(N__44425));
    InMux I__9714 (
            .O(N__44443),
            .I(N__44425));
    LocalMux I__9713 (
            .O(N__44440),
            .I(N__44422));
    Span4Mux_h I__9712 (
            .O(N__44437),
            .I(N__44415));
    Span4Mux_v I__9711 (
            .O(N__44434),
            .I(N__44415));
    LocalMux I__9710 (
            .O(N__44431),
            .I(N__44415));
    InMux I__9709 (
            .O(N__44430),
            .I(N__44412));
    LocalMux I__9708 (
            .O(N__44425),
            .I(N__44406));
    Span12Mux_v I__9707 (
            .O(N__44422),
            .I(N__44403));
    Span4Mux_h I__9706 (
            .O(N__44415),
            .I(N__44400));
    LocalMux I__9705 (
            .O(N__44412),
            .I(N__44397));
    InMux I__9704 (
            .O(N__44411),
            .I(N__44390));
    InMux I__9703 (
            .O(N__44410),
            .I(N__44390));
    InMux I__9702 (
            .O(N__44409),
            .I(N__44390));
    Span4Mux_h I__9701 (
            .O(N__44406),
            .I(N__44387));
    Odrv12 I__9700 (
            .O(N__44403),
            .I(N_142));
    Odrv4 I__9699 (
            .O(N__44400),
            .I(N_142));
    Odrv4 I__9698 (
            .O(N__44397),
            .I(N_142));
    LocalMux I__9697 (
            .O(N__44390),
            .I(N_142));
    Odrv4 I__9696 (
            .O(N__44387),
            .I(N_142));
    InMux I__9695 (
            .O(N__44376),
            .I(N__44373));
    LocalMux I__9694 (
            .O(N__44373),
            .I(N__44370));
    Odrv4 I__9693 (
            .O(N__44370),
            .I(sDAC_mem_42Z0Z_5));
    InMux I__9692 (
            .O(N__44367),
            .I(N__44364));
    LocalMux I__9691 (
            .O(N__44364),
            .I(N__44361));
    Span4Mux_h I__9690 (
            .O(N__44361),
            .I(N__44358));
    Odrv4 I__9689 (
            .O(N__44358),
            .I(sDAC_mem_42Z0Z_6));
    InMux I__9688 (
            .O(N__44355),
            .I(N__44352));
    LocalMux I__9687 (
            .O(N__44352),
            .I(N__44349));
    Span4Mux_h I__9686 (
            .O(N__44349),
            .I(N__44346));
    Span4Mux_h I__9685 (
            .O(N__44346),
            .I(N__44343));
    Odrv4 I__9684 (
            .O(N__44343),
            .I(sDAC_mem_42Z0Z_7));
    InMux I__9683 (
            .O(N__44340),
            .I(N__44337));
    LocalMux I__9682 (
            .O(N__44337),
            .I(N__44334));
    Odrv4 I__9681 (
            .O(N__44334),
            .I(sDAC_mem_10Z0Z_0));
    InMux I__9680 (
            .O(N__44331),
            .I(N__44328));
    LocalMux I__9679 (
            .O(N__44328),
            .I(N__44325));
    Span4Mux_v I__9678 (
            .O(N__44325),
            .I(N__44322));
    Odrv4 I__9677 (
            .O(N__44322),
            .I(sDAC_mem_10Z0Z_1));
    InMux I__9676 (
            .O(N__44319),
            .I(N__44316));
    LocalMux I__9675 (
            .O(N__44316),
            .I(N__44313));
    Span4Mux_h I__9674 (
            .O(N__44313),
            .I(N__44310));
    Span4Mux_h I__9673 (
            .O(N__44310),
            .I(N__44307));
    Odrv4 I__9672 (
            .O(N__44307),
            .I(sDAC_mem_10Z0Z_2));
    InMux I__9671 (
            .O(N__44304),
            .I(N__44301));
    LocalMux I__9670 (
            .O(N__44301),
            .I(N__44298));
    Span4Mux_h I__9669 (
            .O(N__44298),
            .I(N__44295));
    Odrv4 I__9668 (
            .O(N__44295),
            .I(sDAC_mem_10Z0Z_3));
    InMux I__9667 (
            .O(N__44292),
            .I(N__44289));
    LocalMux I__9666 (
            .O(N__44289),
            .I(N__44286));
    Span4Mux_h I__9665 (
            .O(N__44286),
            .I(N__44283));
    Span4Mux_h I__9664 (
            .O(N__44283),
            .I(N__44280));
    Odrv4 I__9663 (
            .O(N__44280),
            .I(sDAC_mem_10Z0Z_4));
    InMux I__9662 (
            .O(N__44277),
            .I(N__44274));
    LocalMux I__9661 (
            .O(N__44274),
            .I(sDAC_mem_10Z0Z_5));
    InMux I__9660 (
            .O(N__44271),
            .I(N__44268));
    LocalMux I__9659 (
            .O(N__44268),
            .I(N__44265));
    Span4Mux_h I__9658 (
            .O(N__44265),
            .I(N__44262));
    Odrv4 I__9657 (
            .O(N__44262),
            .I(sDAC_mem_10Z0Z_6));
    InMux I__9656 (
            .O(N__44259),
            .I(N__44256));
    LocalMux I__9655 (
            .O(N__44256),
            .I(N__44253));
    Span4Mux_v I__9654 (
            .O(N__44253),
            .I(N__44250));
    Span4Mux_h I__9653 (
            .O(N__44250),
            .I(N__44247));
    Odrv4 I__9652 (
            .O(N__44247),
            .I(sDAC_mem_41Z0Z_4));
    InMux I__9651 (
            .O(N__44244),
            .I(N__44241));
    LocalMux I__9650 (
            .O(N__44241),
            .I(N__44238));
    Span4Mux_h I__9649 (
            .O(N__44238),
            .I(N__44235));
    Odrv4 I__9648 (
            .O(N__44235),
            .I(sDAC_mem_41Z0Z_5));
    InMux I__9647 (
            .O(N__44232),
            .I(N__44229));
    LocalMux I__9646 (
            .O(N__44229),
            .I(N__44226));
    Span4Mux_h I__9645 (
            .O(N__44226),
            .I(N__44223));
    Odrv4 I__9644 (
            .O(N__44223),
            .I(sDAC_mem_41Z0Z_6));
    InMux I__9643 (
            .O(N__44220),
            .I(N__44217));
    LocalMux I__9642 (
            .O(N__44217),
            .I(N__44214));
    Span4Mux_v I__9641 (
            .O(N__44214),
            .I(N__44211));
    Odrv4 I__9640 (
            .O(N__44211),
            .I(sDAC_mem_41Z0Z_7));
    InMux I__9639 (
            .O(N__44208),
            .I(N__44205));
    LocalMux I__9638 (
            .O(N__44205),
            .I(N__44202));
    Span4Mux_v I__9637 (
            .O(N__44202),
            .I(N__44199));
    Odrv4 I__9636 (
            .O(N__44199),
            .I(sDAC_mem_42Z0Z_0));
    InMux I__9635 (
            .O(N__44196),
            .I(N__44193));
    LocalMux I__9634 (
            .O(N__44193),
            .I(N__44190));
    Span4Mux_v I__9633 (
            .O(N__44190),
            .I(N__44187));
    Odrv4 I__9632 (
            .O(N__44187),
            .I(sDAC_mem_42Z0Z_1));
    InMux I__9631 (
            .O(N__44184),
            .I(N__44181));
    LocalMux I__9630 (
            .O(N__44181),
            .I(N__44178));
    Span12Mux_h I__9629 (
            .O(N__44178),
            .I(N__44175));
    Odrv12 I__9628 (
            .O(N__44175),
            .I(sDAC_mem_42Z0Z_2));
    InMux I__9627 (
            .O(N__44172),
            .I(N__44169));
    LocalMux I__9626 (
            .O(N__44169),
            .I(N__44166));
    Span4Mux_v I__9625 (
            .O(N__44166),
            .I(N__44163));
    Span4Mux_h I__9624 (
            .O(N__44163),
            .I(N__44160));
    Odrv4 I__9623 (
            .O(N__44160),
            .I(sDAC_mem_42Z0Z_3));
    InMux I__9622 (
            .O(N__44157),
            .I(N__44154));
    LocalMux I__9621 (
            .O(N__44154),
            .I(N__44151));
    Odrv12 I__9620 (
            .O(N__44151),
            .I(sDAC_mem_42Z0Z_4));
    InMux I__9619 (
            .O(N__44148),
            .I(N__44145));
    LocalMux I__9618 (
            .O(N__44145),
            .I(sDAC_mem_12Z0Z_5));
    CascadeMux I__9617 (
            .O(N__44142),
            .I(N__44139));
    InMux I__9616 (
            .O(N__44139),
            .I(N__44136));
    LocalMux I__9615 (
            .O(N__44136),
            .I(N__44133));
    Span4Mux_h I__9614 (
            .O(N__44133),
            .I(N__44130));
    Odrv4 I__9613 (
            .O(N__44130),
            .I(sEEADC_freqZ0Z_1));
    CEMux I__9612 (
            .O(N__44127),
            .I(N__44123));
    CEMux I__9611 (
            .O(N__44126),
            .I(N__44119));
    LocalMux I__9610 (
            .O(N__44123),
            .I(N__44116));
    CEMux I__9609 (
            .O(N__44122),
            .I(N__44113));
    LocalMux I__9608 (
            .O(N__44119),
            .I(N__44110));
    Span4Mux_h I__9607 (
            .O(N__44116),
            .I(N__44105));
    LocalMux I__9606 (
            .O(N__44113),
            .I(N__44105));
    Span4Mux_h I__9605 (
            .O(N__44110),
            .I(N__44102));
    Span4Mux_h I__9604 (
            .O(N__44105),
            .I(N__44099));
    Odrv4 I__9603 (
            .O(N__44102),
            .I(sEEADC_freq_1_sqmuxa));
    Odrv4 I__9602 (
            .O(N__44099),
            .I(sEEADC_freq_1_sqmuxa));
    InMux I__9601 (
            .O(N__44094),
            .I(N__44091));
    LocalMux I__9600 (
            .O(N__44091),
            .I(N__44088));
    Span12Mux_h I__9599 (
            .O(N__44088),
            .I(N__44085));
    Odrv12 I__9598 (
            .O(N__44085),
            .I(sDAC_mem_17Z0Z_0));
    InMux I__9597 (
            .O(N__44082),
            .I(N__44079));
    LocalMux I__9596 (
            .O(N__44079),
            .I(N__44076));
    Span4Mux_h I__9595 (
            .O(N__44076),
            .I(N__44073));
    Odrv4 I__9594 (
            .O(N__44073),
            .I(sDAC_mem_16Z0Z_0));
    CascadeMux I__9593 (
            .O(N__44070),
            .I(N__44067));
    InMux I__9592 (
            .O(N__44067),
            .I(N__44064));
    LocalMux I__9591 (
            .O(N__44064),
            .I(N__44061));
    Span4Mux_v I__9590 (
            .O(N__44061),
            .I(N__44058));
    Odrv4 I__9589 (
            .O(N__44058),
            .I(sDAC_data_RNO_29Z0Z_3));
    InMux I__9588 (
            .O(N__44055),
            .I(N__44052));
    LocalMux I__9587 (
            .O(N__44052),
            .I(N__44049));
    Odrv12 I__9586 (
            .O(N__44049),
            .I(sDAC_mem_16Z0Z_3));
    InMux I__9585 (
            .O(N__44046),
            .I(N__44043));
    LocalMux I__9584 (
            .O(N__44043),
            .I(N__44040));
    Span4Mux_v I__9583 (
            .O(N__44040),
            .I(N__44037));
    Span4Mux_v I__9582 (
            .O(N__44037),
            .I(N__44034));
    Odrv4 I__9581 (
            .O(N__44034),
            .I(sDAC_mem_20Z0Z_7));
    CEMux I__9580 (
            .O(N__44031),
            .I(N__44026));
    CEMux I__9579 (
            .O(N__44030),
            .I(N__44023));
    CEMux I__9578 (
            .O(N__44029),
            .I(N__44020));
    LocalMux I__9577 (
            .O(N__44026),
            .I(N__44017));
    LocalMux I__9576 (
            .O(N__44023),
            .I(N__44014));
    LocalMux I__9575 (
            .O(N__44020),
            .I(N__44011));
    Span4Mux_h I__9574 (
            .O(N__44017),
            .I(N__44008));
    Span4Mux_h I__9573 (
            .O(N__44014),
            .I(N__44003));
    Span4Mux_h I__9572 (
            .O(N__44011),
            .I(N__44003));
    Odrv4 I__9571 (
            .O(N__44008),
            .I(sDAC_mem_20_1_sqmuxa));
    Odrv4 I__9570 (
            .O(N__44003),
            .I(sDAC_mem_20_1_sqmuxa));
    InMux I__9569 (
            .O(N__43998),
            .I(N__43995));
    LocalMux I__9568 (
            .O(N__43995),
            .I(N__43992));
    Span4Mux_v I__9567 (
            .O(N__43992),
            .I(N__43989));
    Odrv4 I__9566 (
            .O(N__43989),
            .I(sDAC_mem_41Z0Z_0));
    InMux I__9565 (
            .O(N__43986),
            .I(N__43983));
    LocalMux I__9564 (
            .O(N__43983),
            .I(N__43980));
    Span4Mux_v I__9563 (
            .O(N__43980),
            .I(N__43977));
    Odrv4 I__9562 (
            .O(N__43977),
            .I(sDAC_mem_41Z0Z_1));
    InMux I__9561 (
            .O(N__43974),
            .I(N__43971));
    LocalMux I__9560 (
            .O(N__43971),
            .I(N__43968));
    Span4Mux_h I__9559 (
            .O(N__43968),
            .I(N__43965));
    Span4Mux_h I__9558 (
            .O(N__43965),
            .I(N__43962));
    Odrv4 I__9557 (
            .O(N__43962),
            .I(sDAC_mem_41Z0Z_2));
    InMux I__9556 (
            .O(N__43959),
            .I(N__43956));
    LocalMux I__9555 (
            .O(N__43956),
            .I(N__43953));
    Span4Mux_h I__9554 (
            .O(N__43953),
            .I(N__43950));
    Odrv4 I__9553 (
            .O(N__43950),
            .I(sDAC_mem_41Z0Z_3));
    InMux I__9552 (
            .O(N__43947),
            .I(N__43944));
    LocalMux I__9551 (
            .O(N__43944),
            .I(N__43941));
    Span4Mux_h I__9550 (
            .O(N__43941),
            .I(N__43938));
    Odrv4 I__9549 (
            .O(N__43938),
            .I(sDAC_mem_14Z0Z_6));
    CEMux I__9548 (
            .O(N__43935),
            .I(N__43932));
    LocalMux I__9547 (
            .O(N__43932),
            .I(sDAC_mem_14_1_sqmuxa));
    InMux I__9546 (
            .O(N__43929),
            .I(N__43926));
    LocalMux I__9545 (
            .O(N__43926),
            .I(sDAC_mem_14Z0Z_4));
    CascadeMux I__9544 (
            .O(N__43923),
            .I(sDAC_data_RNO_18Z0Z_7_cascade_));
    InMux I__9543 (
            .O(N__43920),
            .I(N__43917));
    LocalMux I__9542 (
            .O(N__43917),
            .I(sDAC_data_RNO_19Z0Z_7));
    InMux I__9541 (
            .O(N__43914),
            .I(N__43911));
    LocalMux I__9540 (
            .O(N__43911),
            .I(N__43908));
    Span4Mux_h I__9539 (
            .O(N__43908),
            .I(N__43905));
    Span4Mux_v I__9538 (
            .O(N__43905),
            .I(N__43902));
    Odrv4 I__9537 (
            .O(N__43902),
            .I(sDAC_data_2_24_ns_1_7));
    CascadeMux I__9536 (
            .O(N__43899),
            .I(sDAC_data_RNO_18Z0Z_8_cascade_));
    InMux I__9535 (
            .O(N__43896),
            .I(N__43893));
    LocalMux I__9534 (
            .O(N__43893),
            .I(N__43890));
    Odrv12 I__9533 (
            .O(N__43890),
            .I(sDAC_data_2_24_ns_1_8));
    InMux I__9532 (
            .O(N__43887),
            .I(N__43884));
    LocalMux I__9531 (
            .O(N__43884),
            .I(sDAC_mem_12Z0Z_4));
    InMux I__9530 (
            .O(N__43881),
            .I(N__43878));
    LocalMux I__9529 (
            .O(N__43878),
            .I(sDAC_mem_14Z0Z_5));
    InMux I__9528 (
            .O(N__43875),
            .I(N__43872));
    LocalMux I__9527 (
            .O(N__43872),
            .I(sDAC_data_RNO_19Z0Z_8));
    InMux I__9526 (
            .O(N__43869),
            .I(N__43863));
    InMux I__9525 (
            .O(N__43868),
            .I(N__43863));
    LocalMux I__9524 (
            .O(N__43863),
            .I(N__43857));
    InMux I__9523 (
            .O(N__43862),
            .I(N__43848));
    InMux I__9522 (
            .O(N__43861),
            .I(N__43848));
    InMux I__9521 (
            .O(N__43860),
            .I(N__43848));
    Span4Mux_v I__9520 (
            .O(N__43857),
            .I(N__43840));
    InMux I__9519 (
            .O(N__43856),
            .I(N__43837));
    InMux I__9518 (
            .O(N__43855),
            .I(N__43834));
    LocalMux I__9517 (
            .O(N__43848),
            .I(N__43829));
    InMux I__9516 (
            .O(N__43847),
            .I(N__43824));
    InMux I__9515 (
            .O(N__43846),
            .I(N__43824));
    InMux I__9514 (
            .O(N__43845),
            .I(N__43817));
    InMux I__9513 (
            .O(N__43844),
            .I(N__43817));
    InMux I__9512 (
            .O(N__43843),
            .I(N__43817));
    Span4Mux_h I__9511 (
            .O(N__43840),
            .I(N__43812));
    LocalMux I__9510 (
            .O(N__43837),
            .I(N__43812));
    LocalMux I__9509 (
            .O(N__43834),
            .I(N__43809));
    InMux I__9508 (
            .O(N__43833),
            .I(N__43806));
    InMux I__9507 (
            .O(N__43832),
            .I(N__43803));
    Span4Mux_v I__9506 (
            .O(N__43829),
            .I(N__43800));
    LocalMux I__9505 (
            .O(N__43824),
            .I(N__43797));
    LocalMux I__9504 (
            .O(N__43817),
            .I(N__43792));
    Span4Mux_h I__9503 (
            .O(N__43812),
            .I(N__43792));
    Odrv12 I__9502 (
            .O(N__43809),
            .I(sPointerZ0Z_1));
    LocalMux I__9501 (
            .O(N__43806),
            .I(sPointerZ0Z_1));
    LocalMux I__9500 (
            .O(N__43803),
            .I(sPointerZ0Z_1));
    Odrv4 I__9499 (
            .O(N__43800),
            .I(sPointerZ0Z_1));
    Odrv12 I__9498 (
            .O(N__43797),
            .I(sPointerZ0Z_1));
    Odrv4 I__9497 (
            .O(N__43792),
            .I(sPointerZ0Z_1));
    CEMux I__9496 (
            .O(N__43779),
            .I(N__43776));
    LocalMux I__9495 (
            .O(N__43776),
            .I(N__43772));
    CEMux I__9494 (
            .O(N__43775),
            .I(N__43768));
    Span4Mux_v I__9493 (
            .O(N__43772),
            .I(N__43765));
    CEMux I__9492 (
            .O(N__43771),
            .I(N__43762));
    LocalMux I__9491 (
            .O(N__43768),
            .I(N__43759));
    Span4Mux_h I__9490 (
            .O(N__43765),
            .I(N__43754));
    LocalMux I__9489 (
            .O(N__43762),
            .I(N__43754));
    Span4Mux_v I__9488 (
            .O(N__43759),
            .I(N__43751));
    Sp12to4 I__9487 (
            .O(N__43754),
            .I(N__43748));
    Span4Mux_h I__9486 (
            .O(N__43751),
            .I(N__43745));
    Odrv12 I__9485 (
            .O(N__43748),
            .I(un1_spointer11_0));
    Odrv4 I__9484 (
            .O(N__43745),
            .I(un1_spointer11_0));
    InMux I__9483 (
            .O(N__43740),
            .I(N__43737));
    LocalMux I__9482 (
            .O(N__43737),
            .I(N__43734));
    Span4Mux_v I__9481 (
            .O(N__43734),
            .I(N__43731));
    Odrv4 I__9480 (
            .O(N__43731),
            .I(sDAC_mem_14Z0Z_2));
    InMux I__9479 (
            .O(N__43728),
            .I(N__43725));
    LocalMux I__9478 (
            .O(N__43725),
            .I(N__43722));
    Span4Mux_h I__9477 (
            .O(N__43722),
            .I(N__43719));
    Odrv4 I__9476 (
            .O(N__43719),
            .I(sDAC_mem_14Z0Z_3));
    InMux I__9475 (
            .O(N__43716),
            .I(N__43713));
    LocalMux I__9474 (
            .O(N__43713),
            .I(N__43710));
    Odrv12 I__9473 (
            .O(N__43710),
            .I(sDAC_mem_40Z0Z_1));
    InMux I__9472 (
            .O(N__43707),
            .I(N__43704));
    LocalMux I__9471 (
            .O(N__43704),
            .I(N__43701));
    Span4Mux_h I__9470 (
            .O(N__43701),
            .I(N__43698));
    Span4Mux_v I__9469 (
            .O(N__43698),
            .I(N__43695));
    Odrv4 I__9468 (
            .O(N__43695),
            .I(sDAC_mem_8Z0Z_1));
    CascadeMux I__9467 (
            .O(N__43692),
            .I(sDAC_data_2_20_am_1_4_cascade_));
    CascadeMux I__9466 (
            .O(N__43689),
            .I(N__43683));
    CascadeMux I__9465 (
            .O(N__43688),
            .I(N__43679));
    CascadeMux I__9464 (
            .O(N__43687),
            .I(N__43675));
    CascadeMux I__9463 (
            .O(N__43686),
            .I(N__43662));
    InMux I__9462 (
            .O(N__43683),
            .I(N__43659));
    InMux I__9461 (
            .O(N__43682),
            .I(N__43654));
    InMux I__9460 (
            .O(N__43679),
            .I(N__43654));
    InMux I__9459 (
            .O(N__43678),
            .I(N__43647));
    InMux I__9458 (
            .O(N__43675),
            .I(N__43647));
    InMux I__9457 (
            .O(N__43674),
            .I(N__43647));
    CascadeMux I__9456 (
            .O(N__43673),
            .I(N__43644));
    CascadeMux I__9455 (
            .O(N__43672),
            .I(N__43641));
    CascadeMux I__9454 (
            .O(N__43671),
            .I(N__43638));
    CascadeMux I__9453 (
            .O(N__43670),
            .I(N__43630));
    CascadeMux I__9452 (
            .O(N__43669),
            .I(N__43625));
    CascadeMux I__9451 (
            .O(N__43668),
            .I(N__43617));
    CascadeMux I__9450 (
            .O(N__43667),
            .I(N__43614));
    CascadeMux I__9449 (
            .O(N__43666),
            .I(N__43611));
    CascadeMux I__9448 (
            .O(N__43665),
            .I(N__43608));
    InMux I__9447 (
            .O(N__43662),
            .I(N__43603));
    LocalMux I__9446 (
            .O(N__43659),
            .I(N__43596));
    LocalMux I__9445 (
            .O(N__43654),
            .I(N__43596));
    LocalMux I__9444 (
            .O(N__43647),
            .I(N__43596));
    InMux I__9443 (
            .O(N__43644),
            .I(N__43591));
    InMux I__9442 (
            .O(N__43641),
            .I(N__43591));
    InMux I__9441 (
            .O(N__43638),
            .I(N__43588));
    CascadeMux I__9440 (
            .O(N__43637),
            .I(N__43585));
    CascadeMux I__9439 (
            .O(N__43636),
            .I(N__43582));
    CascadeMux I__9438 (
            .O(N__43635),
            .I(N__43572));
    CascadeMux I__9437 (
            .O(N__43634),
            .I(N__43569));
    CascadeMux I__9436 (
            .O(N__43633),
            .I(N__43566));
    InMux I__9435 (
            .O(N__43630),
            .I(N__43559));
    InMux I__9434 (
            .O(N__43629),
            .I(N__43559));
    InMux I__9433 (
            .O(N__43628),
            .I(N__43556));
    InMux I__9432 (
            .O(N__43625),
            .I(N__43551));
    InMux I__9431 (
            .O(N__43624),
            .I(N__43551));
    CascadeMux I__9430 (
            .O(N__43623),
            .I(N__43547));
    CascadeMux I__9429 (
            .O(N__43622),
            .I(N__43544));
    CascadeMux I__9428 (
            .O(N__43621),
            .I(N__43539));
    CascadeMux I__9427 (
            .O(N__43620),
            .I(N__43536));
    InMux I__9426 (
            .O(N__43617),
            .I(N__43533));
    InMux I__9425 (
            .O(N__43614),
            .I(N__43528));
    InMux I__9424 (
            .O(N__43611),
            .I(N__43528));
    InMux I__9423 (
            .O(N__43608),
            .I(N__43521));
    InMux I__9422 (
            .O(N__43607),
            .I(N__43521));
    InMux I__9421 (
            .O(N__43606),
            .I(N__43521));
    LocalMux I__9420 (
            .O(N__43603),
            .I(N__43508));
    Span4Mux_v I__9419 (
            .O(N__43596),
            .I(N__43508));
    LocalMux I__9418 (
            .O(N__43591),
            .I(N__43503));
    LocalMux I__9417 (
            .O(N__43588),
            .I(N__43503));
    InMux I__9416 (
            .O(N__43585),
            .I(N__43495));
    InMux I__9415 (
            .O(N__43582),
            .I(N__43495));
    InMux I__9414 (
            .O(N__43581),
            .I(N__43492));
    InMux I__9413 (
            .O(N__43580),
            .I(N__43489));
    InMux I__9412 (
            .O(N__43579),
            .I(N__43480));
    InMux I__9411 (
            .O(N__43578),
            .I(N__43480));
    InMux I__9410 (
            .O(N__43577),
            .I(N__43480));
    InMux I__9409 (
            .O(N__43576),
            .I(N__43480));
    CascadeMux I__9408 (
            .O(N__43575),
            .I(N__43476));
    InMux I__9407 (
            .O(N__43572),
            .I(N__43473));
    InMux I__9406 (
            .O(N__43569),
            .I(N__43468));
    InMux I__9405 (
            .O(N__43566),
            .I(N__43468));
    CascadeMux I__9404 (
            .O(N__43565),
            .I(N__43465));
    CascadeMux I__9403 (
            .O(N__43564),
            .I(N__43462));
    LocalMux I__9402 (
            .O(N__43559),
            .I(N__43455));
    LocalMux I__9401 (
            .O(N__43556),
            .I(N__43455));
    LocalMux I__9400 (
            .O(N__43551),
            .I(N__43455));
    CascadeMux I__9399 (
            .O(N__43550),
            .I(N__43452));
    InMux I__9398 (
            .O(N__43547),
            .I(N__43441));
    InMux I__9397 (
            .O(N__43544),
            .I(N__43441));
    InMux I__9396 (
            .O(N__43543),
            .I(N__43441));
    InMux I__9395 (
            .O(N__43542),
            .I(N__43434));
    InMux I__9394 (
            .O(N__43539),
            .I(N__43434));
    InMux I__9393 (
            .O(N__43536),
            .I(N__43434));
    LocalMux I__9392 (
            .O(N__43533),
            .I(N__43429));
    LocalMux I__9391 (
            .O(N__43528),
            .I(N__43429));
    LocalMux I__9390 (
            .O(N__43521),
            .I(N__43426));
    InMux I__9389 (
            .O(N__43520),
            .I(N__43417));
    InMux I__9388 (
            .O(N__43519),
            .I(N__43417));
    InMux I__9387 (
            .O(N__43518),
            .I(N__43417));
    InMux I__9386 (
            .O(N__43517),
            .I(N__43417));
    InMux I__9385 (
            .O(N__43516),
            .I(N__43408));
    InMux I__9384 (
            .O(N__43515),
            .I(N__43408));
    InMux I__9383 (
            .O(N__43514),
            .I(N__43408));
    InMux I__9382 (
            .O(N__43513),
            .I(N__43408));
    Span4Mux_h I__9381 (
            .O(N__43508),
            .I(N__43403));
    Span4Mux_h I__9380 (
            .O(N__43503),
            .I(N__43403));
    InMux I__9379 (
            .O(N__43502),
            .I(N__43396));
    InMux I__9378 (
            .O(N__43501),
            .I(N__43396));
    InMux I__9377 (
            .O(N__43500),
            .I(N__43396));
    LocalMux I__9376 (
            .O(N__43495),
            .I(N__43387));
    LocalMux I__9375 (
            .O(N__43492),
            .I(N__43387));
    LocalMux I__9374 (
            .O(N__43489),
            .I(N__43387));
    LocalMux I__9373 (
            .O(N__43480),
            .I(N__43387));
    InMux I__9372 (
            .O(N__43479),
            .I(N__43384));
    InMux I__9371 (
            .O(N__43476),
            .I(N__43381));
    LocalMux I__9370 (
            .O(N__43473),
            .I(N__43376));
    LocalMux I__9369 (
            .O(N__43468),
            .I(N__43376));
    InMux I__9368 (
            .O(N__43465),
            .I(N__43371));
    InMux I__9367 (
            .O(N__43462),
            .I(N__43371));
    Span4Mux_v I__9366 (
            .O(N__43455),
            .I(N__43368));
    InMux I__9365 (
            .O(N__43452),
            .I(N__43365));
    InMux I__9364 (
            .O(N__43451),
            .I(N__43356));
    InMux I__9363 (
            .O(N__43450),
            .I(N__43356));
    InMux I__9362 (
            .O(N__43449),
            .I(N__43356));
    InMux I__9361 (
            .O(N__43448),
            .I(N__43356));
    LocalMux I__9360 (
            .O(N__43441),
            .I(N__43353));
    LocalMux I__9359 (
            .O(N__43434),
            .I(N__43344));
    Span4Mux_v I__9358 (
            .O(N__43429),
            .I(N__43344));
    Span4Mux_h I__9357 (
            .O(N__43426),
            .I(N__43344));
    LocalMux I__9356 (
            .O(N__43417),
            .I(N__43344));
    LocalMux I__9355 (
            .O(N__43408),
            .I(N__43337));
    Span4Mux_v I__9354 (
            .O(N__43403),
            .I(N__43337));
    LocalMux I__9353 (
            .O(N__43396),
            .I(N__43337));
    Span4Mux_h I__9352 (
            .O(N__43387),
            .I(N__43334));
    LocalMux I__9351 (
            .O(N__43384),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9350 (
            .O(N__43381),
            .I(sDAC_mem_pointerZ0Z_5));
    Odrv4 I__9349 (
            .O(N__43376),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9348 (
            .O(N__43371),
            .I(sDAC_mem_pointerZ0Z_5));
    Odrv4 I__9347 (
            .O(N__43368),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9346 (
            .O(N__43365),
            .I(sDAC_mem_pointerZ0Z_5));
    LocalMux I__9345 (
            .O(N__43356),
            .I(sDAC_mem_pointerZ0Z_5));
    Odrv12 I__9344 (
            .O(N__43353),
            .I(sDAC_mem_pointerZ0Z_5));
    Odrv4 I__9343 (
            .O(N__43344),
            .I(sDAC_mem_pointerZ0Z_5));
    Odrv4 I__9342 (
            .O(N__43337),
            .I(sDAC_mem_pointerZ0Z_5));
    Odrv4 I__9341 (
            .O(N__43334),
            .I(sDAC_mem_pointerZ0Z_5));
    CascadeMux I__9340 (
            .O(N__43311),
            .I(sDAC_data_RNO_17Z0Z_4_cascade_));
    CascadeMux I__9339 (
            .O(N__43308),
            .I(sDAC_data_RNO_8Z0Z_4_cascade_));
    InMux I__9338 (
            .O(N__43305),
            .I(N__43302));
    LocalMux I__9337 (
            .O(N__43302),
            .I(sDAC_data_RNO_7Z0Z_4));
    InMux I__9336 (
            .O(N__43299),
            .I(N__43296));
    LocalMux I__9335 (
            .O(N__43296),
            .I(N__43293));
    Odrv4 I__9334 (
            .O(N__43293),
            .I(sDAC_data_RNO_2Z0Z_4));
    CascadeMux I__9333 (
            .O(N__43290),
            .I(N_284_cascade_));
    InMux I__9332 (
            .O(N__43287),
            .I(N__43284));
    LocalMux I__9331 (
            .O(N__43284),
            .I(N__43278));
    InMux I__9330 (
            .O(N__43283),
            .I(N__43273));
    InMux I__9329 (
            .O(N__43282),
            .I(N__43273));
    InMux I__9328 (
            .O(N__43281),
            .I(N__43270));
    Span4Mux_v I__9327 (
            .O(N__43278),
            .I(N__43266));
    LocalMux I__9326 (
            .O(N__43273),
            .I(N__43261));
    LocalMux I__9325 (
            .O(N__43270),
            .I(N__43261));
    InMux I__9324 (
            .O(N__43269),
            .I(N__43257));
    Span4Mux_h I__9323 (
            .O(N__43266),
            .I(N__43249));
    Span4Mux_v I__9322 (
            .O(N__43261),
            .I(N__43249));
    InMux I__9321 (
            .O(N__43260),
            .I(N__43246));
    LocalMux I__9320 (
            .O(N__43257),
            .I(N__43243));
    InMux I__9319 (
            .O(N__43256),
            .I(N__43238));
    InMux I__9318 (
            .O(N__43255),
            .I(N__43238));
    InMux I__9317 (
            .O(N__43254),
            .I(N__43235));
    Span4Mux_h I__9316 (
            .O(N__43249),
            .I(N__43230));
    LocalMux I__9315 (
            .O(N__43246),
            .I(N__43230));
    Span4Mux_h I__9314 (
            .O(N__43243),
            .I(N__43227));
    LocalMux I__9313 (
            .O(N__43238),
            .I(N__43222));
    LocalMux I__9312 (
            .O(N__43235),
            .I(N__43219));
    Span4Mux_v I__9311 (
            .O(N__43230),
            .I(N__43216));
    Span4Mux_h I__9310 (
            .O(N__43227),
            .I(N__43213));
    InMux I__9309 (
            .O(N__43226),
            .I(N__43208));
    InMux I__9308 (
            .O(N__43225),
            .I(N__43208));
    Sp12to4 I__9307 (
            .O(N__43222),
            .I(N__43205));
    Span4Mux_v I__9306 (
            .O(N__43219),
            .I(N__43200));
    Span4Mux_h I__9305 (
            .O(N__43216),
            .I(N__43200));
    Odrv4 I__9304 (
            .O(N__43213),
            .I(N_284));
    LocalMux I__9303 (
            .O(N__43208),
            .I(N_284));
    Odrv12 I__9302 (
            .O(N__43205),
            .I(N_284));
    Odrv4 I__9301 (
            .O(N__43200),
            .I(N_284));
    InMux I__9300 (
            .O(N__43191),
            .I(N__43186));
    InMux I__9299 (
            .O(N__43190),
            .I(N__43183));
    InMux I__9298 (
            .O(N__43189),
            .I(N__43180));
    LocalMux I__9297 (
            .O(N__43186),
            .I(N__43174));
    LocalMux I__9296 (
            .O(N__43183),
            .I(N__43171));
    LocalMux I__9295 (
            .O(N__43180),
            .I(N__43168));
    InMux I__9294 (
            .O(N__43179),
            .I(N__43161));
    InMux I__9293 (
            .O(N__43178),
            .I(N__43161));
    InMux I__9292 (
            .O(N__43177),
            .I(N__43161));
    Span4Mux_h I__9291 (
            .O(N__43174),
            .I(N__43157));
    Span4Mux_v I__9290 (
            .O(N__43171),
            .I(N__43154));
    Span4Mux_v I__9289 (
            .O(N__43168),
            .I(N__43149));
    LocalMux I__9288 (
            .O(N__43161),
            .I(N__43149));
    InMux I__9287 (
            .O(N__43160),
            .I(N__43146));
    Span4Mux_h I__9286 (
            .O(N__43157),
            .I(N__43135));
    Span4Mux_h I__9285 (
            .O(N__43154),
            .I(N__43130));
    Span4Mux_h I__9284 (
            .O(N__43149),
            .I(N__43130));
    LocalMux I__9283 (
            .O(N__43146),
            .I(N__43127));
    InMux I__9282 (
            .O(N__43145),
            .I(N__43120));
    InMux I__9281 (
            .O(N__43144),
            .I(N__43120));
    InMux I__9280 (
            .O(N__43143),
            .I(N__43120));
    InMux I__9279 (
            .O(N__43142),
            .I(N__43115));
    InMux I__9278 (
            .O(N__43141),
            .I(N__43115));
    InMux I__9277 (
            .O(N__43140),
            .I(N__43108));
    InMux I__9276 (
            .O(N__43139),
            .I(N__43108));
    InMux I__9275 (
            .O(N__43138),
            .I(N__43108));
    Odrv4 I__9274 (
            .O(N__43135),
            .I(N_280));
    Odrv4 I__9273 (
            .O(N__43130),
            .I(N_280));
    Odrv4 I__9272 (
            .O(N__43127),
            .I(N_280));
    LocalMux I__9271 (
            .O(N__43120),
            .I(N_280));
    LocalMux I__9270 (
            .O(N__43115),
            .I(N_280));
    LocalMux I__9269 (
            .O(N__43108),
            .I(N_280));
    InMux I__9268 (
            .O(N__43095),
            .I(N__43092));
    LocalMux I__9267 (
            .O(N__43092),
            .I(sDAC_mem_6Z0Z_6));
    CEMux I__9266 (
            .O(N__43089),
            .I(N__43086));
    LocalMux I__9265 (
            .O(N__43086),
            .I(N__43082));
    CEMux I__9264 (
            .O(N__43085),
            .I(N__43079));
    Span4Mux_v I__9263 (
            .O(N__43082),
            .I(N__43075));
    LocalMux I__9262 (
            .O(N__43079),
            .I(N__43072));
    CEMux I__9261 (
            .O(N__43078),
            .I(N__43068));
    Span4Mux_v I__9260 (
            .O(N__43075),
            .I(N__43063));
    Span4Mux_v I__9259 (
            .O(N__43072),
            .I(N__43063));
    CEMux I__9258 (
            .O(N__43071),
            .I(N__43060));
    LocalMux I__9257 (
            .O(N__43068),
            .I(N__43057));
    Sp12to4 I__9256 (
            .O(N__43063),
            .I(N__43054));
    LocalMux I__9255 (
            .O(N__43060),
            .I(N__43051));
    Span4Mux_h I__9254 (
            .O(N__43057),
            .I(N__43048));
    Odrv12 I__9253 (
            .O(N__43054),
            .I(sDAC_mem_6_1_sqmuxa));
    Odrv4 I__9252 (
            .O(N__43051),
            .I(sDAC_mem_6_1_sqmuxa));
    Odrv4 I__9251 (
            .O(N__43048),
            .I(sDAC_mem_6_1_sqmuxa));
    InMux I__9250 (
            .O(N__43041),
            .I(N__43038));
    LocalMux I__9249 (
            .O(N__43038),
            .I(N__43035));
    Odrv12 I__9248 (
            .O(N__43035),
            .I(sDAC_mem_40Z0Z_0));
    InMux I__9247 (
            .O(N__43032),
            .I(N__43029));
    LocalMux I__9246 (
            .O(N__43029),
            .I(N__43026));
    Span4Mux_h I__9245 (
            .O(N__43026),
            .I(N__43023));
    Span4Mux_v I__9244 (
            .O(N__43023),
            .I(N__43020));
    Odrv4 I__9243 (
            .O(N__43020),
            .I(sDAC_mem_8Z0Z_0));
    CascadeMux I__9242 (
            .O(N__43017),
            .I(sDAC_data_2_20_am_1_3_cascade_));
    CascadeMux I__9241 (
            .O(N__43014),
            .I(sDAC_data_RNO_17Z0Z_3_cascade_));
    CascadeMux I__9240 (
            .O(N__43011),
            .I(sDAC_data_RNO_8Z0Z_3_cascade_));
    InMux I__9239 (
            .O(N__43008),
            .I(N__43005));
    LocalMux I__9238 (
            .O(N__43005),
            .I(sDAC_data_RNO_7Z0Z_3));
    InMux I__9237 (
            .O(N__43002),
            .I(N__42999));
    LocalMux I__9236 (
            .O(N__42999),
            .I(sDAC_data_RNO_2Z0Z_3));
    CEMux I__9235 (
            .O(N__42996),
            .I(N__42993));
    LocalMux I__9234 (
            .O(N__42993),
            .I(N__42989));
    CEMux I__9233 (
            .O(N__42992),
            .I(N__42986));
    Span4Mux_h I__9232 (
            .O(N__42989),
            .I(N__42979));
    LocalMux I__9231 (
            .O(N__42986),
            .I(N__42979));
    CEMux I__9230 (
            .O(N__42985),
            .I(N__42974));
    CEMux I__9229 (
            .O(N__42984),
            .I(N__42971));
    Span4Mux_v I__9228 (
            .O(N__42979),
            .I(N__42968));
    CEMux I__9227 (
            .O(N__42978),
            .I(N__42965));
    CEMux I__9226 (
            .O(N__42977),
            .I(N__42962));
    LocalMux I__9225 (
            .O(N__42974),
            .I(N__42957));
    LocalMux I__9224 (
            .O(N__42971),
            .I(N__42954));
    Span4Mux_h I__9223 (
            .O(N__42968),
            .I(N__42951));
    LocalMux I__9222 (
            .O(N__42965),
            .I(N__42948));
    LocalMux I__9221 (
            .O(N__42962),
            .I(N__42945));
    CEMux I__9220 (
            .O(N__42961),
            .I(N__42942));
    CEMux I__9219 (
            .O(N__42960),
            .I(N__42939));
    Span4Mux_h I__9218 (
            .O(N__42957),
            .I(N__42936));
    Span4Mux_v I__9217 (
            .O(N__42954),
            .I(N__42933));
    Span4Mux_h I__9216 (
            .O(N__42951),
            .I(N__42922));
    Span4Mux_v I__9215 (
            .O(N__42948),
            .I(N__42922));
    Span4Mux_h I__9214 (
            .O(N__42945),
            .I(N__42922));
    LocalMux I__9213 (
            .O(N__42942),
            .I(N__42922));
    LocalMux I__9212 (
            .O(N__42939),
            .I(N__42922));
    Span4Mux_v I__9211 (
            .O(N__42936),
            .I(N__42919));
    Span4Mux_h I__9210 (
            .O(N__42933),
            .I(N__42916));
    Sp12to4 I__9209 (
            .O(N__42922),
            .I(N__42913));
    Odrv4 I__9208 (
            .O(N__42919),
            .I(sDAC_mem_3_1_sqmuxa));
    Odrv4 I__9207 (
            .O(N__42916),
            .I(sDAC_mem_3_1_sqmuxa));
    Odrv12 I__9206 (
            .O(N__42913),
            .I(sDAC_mem_3_1_sqmuxa));
    CascadeMux I__9205 (
            .O(N__42906),
            .I(N__42903));
    InMux I__9204 (
            .O(N__42903),
            .I(N__42900));
    LocalMux I__9203 (
            .O(N__42900),
            .I(N__42897));
    Span4Mux_v I__9202 (
            .O(N__42897),
            .I(N__42894));
    Span4Mux_h I__9201 (
            .O(N__42894),
            .I(N__42891));
    Span4Mux_v I__9200 (
            .O(N__42891),
            .I(N__42888));
    Odrv4 I__9199 (
            .O(N__42888),
            .I(sDAC_mem_34Z0Z_7));
    InMux I__9198 (
            .O(N__42885),
            .I(N__42882));
    LocalMux I__9197 (
            .O(N__42882),
            .I(N__42879));
    Span4Mux_v I__9196 (
            .O(N__42879),
            .I(N__42876));
    Span4Mux_h I__9195 (
            .O(N__42876),
            .I(N__42873));
    Odrv4 I__9194 (
            .O(N__42873),
            .I(sDAC_mem_2Z0Z_7));
    InMux I__9193 (
            .O(N__42870),
            .I(N__42867));
    LocalMux I__9192 (
            .O(N__42867),
            .I(N__42864));
    Span4Mux_v I__9191 (
            .O(N__42864),
            .I(N__42861));
    Odrv4 I__9190 (
            .O(N__42861),
            .I(sDAC_mem_35Z0Z_7));
    CascadeMux I__9189 (
            .O(N__42858),
            .I(sDAC_data_2_6_bm_1_10_cascade_));
    InMux I__9188 (
            .O(N__42855),
            .I(N__42852));
    LocalMux I__9187 (
            .O(N__42852),
            .I(sDAC_mem_3Z0Z_7));
    CascadeMux I__9186 (
            .O(N__42849),
            .I(N__42846));
    InMux I__9185 (
            .O(N__42846),
            .I(N__42843));
    LocalMux I__9184 (
            .O(N__42843),
            .I(N__42840));
    Odrv4 I__9183 (
            .O(N__42840),
            .I(sDAC_data_RNO_15Z0Z_10));
    InMux I__9182 (
            .O(N__42837),
            .I(N__42834));
    LocalMux I__9181 (
            .O(N__42834),
            .I(N__42831));
    Span4Mux_v I__9180 (
            .O(N__42831),
            .I(N__42828));
    Odrv4 I__9179 (
            .O(N__42828),
            .I(sDAC_mem_35Z0Z_3));
    CascadeMux I__9178 (
            .O(N__42825),
            .I(sDAC_data_2_6_bm_1_6_cascade_));
    InMux I__9177 (
            .O(N__42822),
            .I(N__42819));
    LocalMux I__9176 (
            .O(N__42819),
            .I(sDAC_mem_3Z0Z_3));
    CascadeMux I__9175 (
            .O(N__42816),
            .I(N__42813));
    InMux I__9174 (
            .O(N__42813),
            .I(N__42810));
    LocalMux I__9173 (
            .O(N__42810),
            .I(sDAC_data_RNO_15Z0Z_6));
    CascadeMux I__9172 (
            .O(N__42807),
            .I(sDAC_data_RNO_17Z0Z_8_cascade_));
    InMux I__9171 (
            .O(N__42804),
            .I(N__42801));
    LocalMux I__9170 (
            .O(N__42801),
            .I(N__42798));
    Odrv12 I__9169 (
            .O(N__42798),
            .I(sDAC_mem_40Z0Z_5));
    InMux I__9168 (
            .O(N__42795),
            .I(N__42792));
    LocalMux I__9167 (
            .O(N__42792),
            .I(N__42789));
    Span4Mux_v I__9166 (
            .O(N__42789),
            .I(N__42786));
    Odrv4 I__9165 (
            .O(N__42786),
            .I(sDAC_mem_8Z0Z_5));
    CascadeMux I__9164 (
            .O(N__42783),
            .I(sDAC_data_2_20_am_1_8_cascade_));
    CascadeMux I__9163 (
            .O(N__42780),
            .I(sDAC_data_RNO_7Z0Z_8_cascade_));
    InMux I__9162 (
            .O(N__42777),
            .I(N__42774));
    LocalMux I__9161 (
            .O(N__42774),
            .I(sDAC_data_RNO_8Z0Z_8));
    InMux I__9160 (
            .O(N__42771),
            .I(N__42768));
    LocalMux I__9159 (
            .O(N__42768),
            .I(sDAC_data_RNO_2Z0Z_8));
    InMux I__9158 (
            .O(N__42765),
            .I(N__42762));
    LocalMux I__9157 (
            .O(N__42762),
            .I(N__42759));
    Odrv12 I__9156 (
            .O(N__42759),
            .I(sDAC_mem_38Z0Z_6));
    InMux I__9155 (
            .O(N__42756),
            .I(N__42753));
    LocalMux I__9154 (
            .O(N__42753),
            .I(N__42750));
    Span4Mux_v I__9153 (
            .O(N__42750),
            .I(N__42747));
    Odrv4 I__9152 (
            .O(N__42747),
            .I(sDAC_mem_39Z0Z_6));
    CascadeMux I__9151 (
            .O(N__42744),
            .I(sDAC_data_2_13_bm_1_9_cascade_));
    InMux I__9150 (
            .O(N__42741),
            .I(N__42738));
    LocalMux I__9149 (
            .O(N__42738),
            .I(N__42735));
    Span4Mux_h I__9148 (
            .O(N__42735),
            .I(N__42732));
    Span4Mux_v I__9147 (
            .O(N__42732),
            .I(N__42729));
    Odrv4 I__9146 (
            .O(N__42729),
            .I(sDAC_mem_7Z0Z_6));
    InMux I__9145 (
            .O(N__42726),
            .I(N__42723));
    LocalMux I__9144 (
            .O(N__42723),
            .I(N__42720));
    Span4Mux_v I__9143 (
            .O(N__42720),
            .I(N__42717));
    Odrv4 I__9142 (
            .O(N__42717),
            .I(sDAC_data_RNO_5Z0Z_9));
    InMux I__9141 (
            .O(N__42714),
            .I(N__42711));
    LocalMux I__9140 (
            .O(N__42711),
            .I(sDAC_data_RNO_14Z0Z_6));
    InMux I__9139 (
            .O(N__42708),
            .I(N__42705));
    LocalMux I__9138 (
            .O(N__42705),
            .I(sDAC_data_2_14_ns_1_6));
    CascadeMux I__9137 (
            .O(N__42702),
            .I(N__42699));
    InMux I__9136 (
            .O(N__42699),
            .I(N__42696));
    LocalMux I__9135 (
            .O(N__42696),
            .I(N__42693));
    Span4Mux_h I__9134 (
            .O(N__42693),
            .I(N__42690));
    Span4Mux_v I__9133 (
            .O(N__42690),
            .I(N__42687));
    Span4Mux_v I__9132 (
            .O(N__42687),
            .I(N__42684));
    Odrv4 I__9131 (
            .O(N__42684),
            .I(sDAC_data_RNO_29Z0Z_6));
    InMux I__9130 (
            .O(N__42681),
            .I(N__42678));
    LocalMux I__9129 (
            .O(N__42678),
            .I(N__42675));
    Span4Mux_h I__9128 (
            .O(N__42675),
            .I(N__42672));
    Odrv4 I__9127 (
            .O(N__42672),
            .I(sDAC_data_RNO_30Z0Z_6));
    InMux I__9126 (
            .O(N__42669),
            .I(N__42666));
    LocalMux I__9125 (
            .O(N__42666),
            .I(N__42663));
    Span4Mux_h I__9124 (
            .O(N__42663),
            .I(N__42660));
    Span4Mux_h I__9123 (
            .O(N__42660),
            .I(N__42657));
    Odrv4 I__9122 (
            .O(N__42657),
            .I(sDAC_data_RNO_21Z0Z_6));
    CascadeMux I__9121 (
            .O(N__42654),
            .I(sDAC_data_2_32_ns_1_6_cascade_));
    InMux I__9120 (
            .O(N__42651),
            .I(N__42648));
    LocalMux I__9119 (
            .O(N__42648),
            .I(N__42645));
    Odrv4 I__9118 (
            .O(N__42645),
            .I(sDAC_data_RNO_20Z0Z_6));
    InMux I__9117 (
            .O(N__42642),
            .I(N__42635));
    InMux I__9116 (
            .O(N__42641),
            .I(N__42632));
    InMux I__9115 (
            .O(N__42640),
            .I(N__42627));
    InMux I__9114 (
            .O(N__42639),
            .I(N__42624));
    InMux I__9113 (
            .O(N__42638),
            .I(N__42620));
    LocalMux I__9112 (
            .O(N__42635),
            .I(N__42615));
    LocalMux I__9111 (
            .O(N__42632),
            .I(N__42615));
    InMux I__9110 (
            .O(N__42631),
            .I(N__42611));
    InMux I__9109 (
            .O(N__42630),
            .I(N__42607));
    LocalMux I__9108 (
            .O(N__42627),
            .I(N__42604));
    LocalMux I__9107 (
            .O(N__42624),
            .I(N__42601));
    InMux I__9106 (
            .O(N__42623),
            .I(N__42598));
    LocalMux I__9105 (
            .O(N__42620),
            .I(N__42595));
    Span4Mux_v I__9104 (
            .O(N__42615),
            .I(N__42592));
    CascadeMux I__9103 (
            .O(N__42614),
            .I(N__42589));
    LocalMux I__9102 (
            .O(N__42611),
            .I(N__42586));
    InMux I__9101 (
            .O(N__42610),
            .I(N__42583));
    LocalMux I__9100 (
            .O(N__42607),
            .I(N__42576));
    Span4Mux_h I__9099 (
            .O(N__42604),
            .I(N__42576));
    Span4Mux_h I__9098 (
            .O(N__42601),
            .I(N__42576));
    LocalMux I__9097 (
            .O(N__42598),
            .I(N__42569));
    Span4Mux_v I__9096 (
            .O(N__42595),
            .I(N__42569));
    Span4Mux_h I__9095 (
            .O(N__42592),
            .I(N__42569));
    InMux I__9094 (
            .O(N__42589),
            .I(N__42566));
    Odrv12 I__9093 (
            .O(N__42586),
            .I(sDAC_mem_pointerZ0Z_3));
    LocalMux I__9092 (
            .O(N__42583),
            .I(sDAC_mem_pointerZ0Z_3));
    Odrv4 I__9091 (
            .O(N__42576),
            .I(sDAC_mem_pointerZ0Z_3));
    Odrv4 I__9090 (
            .O(N__42569),
            .I(sDAC_mem_pointerZ0Z_3));
    LocalMux I__9089 (
            .O(N__42566),
            .I(sDAC_mem_pointerZ0Z_3));
    CascadeMux I__9088 (
            .O(N__42555),
            .I(sDAC_data_RNO_10Z0Z_6_cascade_));
    InMux I__9087 (
            .O(N__42552),
            .I(N__42549));
    LocalMux I__9086 (
            .O(N__42549),
            .I(N__42546));
    Span4Mux_h I__9085 (
            .O(N__42546),
            .I(N__42543));
    Span4Mux_v I__9084 (
            .O(N__42543),
            .I(N__42540));
    Span4Mux_h I__9083 (
            .O(N__42540),
            .I(N__42537));
    Odrv4 I__9082 (
            .O(N__42537),
            .I(sDAC_data_RNO_11Z0Z_6));
    CascadeMux I__9081 (
            .O(N__42534),
            .I(N__42519));
    InMux I__9080 (
            .O(N__42533),
            .I(N__42514));
    InMux I__9079 (
            .O(N__42532),
            .I(N__42511));
    InMux I__9078 (
            .O(N__42531),
            .I(N__42508));
    InMux I__9077 (
            .O(N__42530),
            .I(N__42505));
    InMux I__9076 (
            .O(N__42529),
            .I(N__42500));
    InMux I__9075 (
            .O(N__42528),
            .I(N__42500));
    InMux I__9074 (
            .O(N__42527),
            .I(N__42497));
    InMux I__9073 (
            .O(N__42526),
            .I(N__42492));
    InMux I__9072 (
            .O(N__42525),
            .I(N__42492));
    InMux I__9071 (
            .O(N__42524),
            .I(N__42489));
    InMux I__9070 (
            .O(N__42523),
            .I(N__42484));
    InMux I__9069 (
            .O(N__42522),
            .I(N__42484));
    InMux I__9068 (
            .O(N__42519),
            .I(N__42480));
    InMux I__9067 (
            .O(N__42518),
            .I(N__42476));
    InMux I__9066 (
            .O(N__42517),
            .I(N__42473));
    LocalMux I__9065 (
            .O(N__42514),
            .I(N__42470));
    LocalMux I__9064 (
            .O(N__42511),
            .I(N__42467));
    LocalMux I__9063 (
            .O(N__42508),
            .I(N__42464));
    LocalMux I__9062 (
            .O(N__42505),
            .I(N__42461));
    LocalMux I__9061 (
            .O(N__42500),
            .I(N__42458));
    LocalMux I__9060 (
            .O(N__42497),
            .I(N__42451));
    LocalMux I__9059 (
            .O(N__42492),
            .I(N__42451));
    LocalMux I__9058 (
            .O(N__42489),
            .I(N__42451));
    LocalMux I__9057 (
            .O(N__42484),
            .I(N__42448));
    InMux I__9056 (
            .O(N__42483),
            .I(N__42444));
    LocalMux I__9055 (
            .O(N__42480),
            .I(N__42441));
    InMux I__9054 (
            .O(N__42479),
            .I(N__42438));
    LocalMux I__9053 (
            .O(N__42476),
            .I(N__42429));
    LocalMux I__9052 (
            .O(N__42473),
            .I(N__42429));
    Span4Mux_v I__9051 (
            .O(N__42470),
            .I(N__42429));
    Span4Mux_v I__9050 (
            .O(N__42467),
            .I(N__42429));
    Span4Mux_h I__9049 (
            .O(N__42464),
            .I(N__42426));
    Span4Mux_v I__9048 (
            .O(N__42461),
            .I(N__42417));
    Span4Mux_v I__9047 (
            .O(N__42458),
            .I(N__42417));
    Span4Mux_v I__9046 (
            .O(N__42451),
            .I(N__42417));
    Span4Mux_v I__9045 (
            .O(N__42448),
            .I(N__42417));
    InMux I__9044 (
            .O(N__42447),
            .I(N__42414));
    LocalMux I__9043 (
            .O(N__42444),
            .I(sDAC_mem_pointerZ0Z_4));
    Odrv12 I__9042 (
            .O(N__42441),
            .I(sDAC_mem_pointerZ0Z_4));
    LocalMux I__9041 (
            .O(N__42438),
            .I(sDAC_mem_pointerZ0Z_4));
    Odrv4 I__9040 (
            .O(N__42429),
            .I(sDAC_mem_pointerZ0Z_4));
    Odrv4 I__9039 (
            .O(N__42426),
            .I(sDAC_mem_pointerZ0Z_4));
    Odrv4 I__9038 (
            .O(N__42417),
            .I(sDAC_mem_pointerZ0Z_4));
    LocalMux I__9037 (
            .O(N__42414),
            .I(sDAC_mem_pointerZ0Z_4));
    InMux I__9036 (
            .O(N__42399),
            .I(N__42396));
    LocalMux I__9035 (
            .O(N__42396),
            .I(sDAC_data_RNO_2Z0Z_6));
    CascadeMux I__9034 (
            .O(N__42393),
            .I(sDAC_data_2_41_ns_1_6_cascade_));
    InMux I__9033 (
            .O(N__42390),
            .I(N__42387));
    LocalMux I__9032 (
            .O(N__42387),
            .I(sDAC_data_RNO_1Z0Z_6));
    InMux I__9031 (
            .O(N__42384),
            .I(N__42370));
    InMux I__9030 (
            .O(N__42383),
            .I(N__42367));
    InMux I__9029 (
            .O(N__42382),
            .I(N__42363));
    InMux I__9028 (
            .O(N__42381),
            .I(N__42360));
    InMux I__9027 (
            .O(N__42380),
            .I(N__42357));
    InMux I__9026 (
            .O(N__42379),
            .I(N__42354));
    InMux I__9025 (
            .O(N__42378),
            .I(N__42351));
    InMux I__9024 (
            .O(N__42377),
            .I(N__42348));
    InMux I__9023 (
            .O(N__42376),
            .I(N__42345));
    InMux I__9022 (
            .O(N__42375),
            .I(N__42338));
    InMux I__9021 (
            .O(N__42374),
            .I(N__42338));
    InMux I__9020 (
            .O(N__42373),
            .I(N__42338));
    LocalMux I__9019 (
            .O(N__42370),
            .I(N__42333));
    LocalMux I__9018 (
            .O(N__42367),
            .I(N__42333));
    InMux I__9017 (
            .O(N__42366),
            .I(N__42330));
    LocalMux I__9016 (
            .O(N__42363),
            .I(N__42325));
    LocalMux I__9015 (
            .O(N__42360),
            .I(N__42325));
    LocalMux I__9014 (
            .O(N__42357),
            .I(N__42322));
    LocalMux I__9013 (
            .O(N__42354),
            .I(N__42315));
    LocalMux I__9012 (
            .O(N__42351),
            .I(N__42315));
    LocalMux I__9011 (
            .O(N__42348),
            .I(N__42315));
    LocalMux I__9010 (
            .O(N__42345),
            .I(N__42308));
    LocalMux I__9009 (
            .O(N__42338),
            .I(N__42308));
    Span4Mux_h I__9008 (
            .O(N__42333),
            .I(N__42308));
    LocalMux I__9007 (
            .O(N__42330),
            .I(N__42305));
    Span4Mux_h I__9006 (
            .O(N__42325),
            .I(N__42302));
    Span4Mux_v I__9005 (
            .O(N__42322),
            .I(N__42299));
    Span4Mux_h I__9004 (
            .O(N__42315),
            .I(N__42295));
    Span4Mux_v I__9003 (
            .O(N__42308),
            .I(N__42292));
    Span4Mux_h I__9002 (
            .O(N__42305),
            .I(N__42289));
    Span4Mux_v I__9001 (
            .O(N__42302),
            .I(N__42286));
    Span4Mux_v I__9000 (
            .O(N__42299),
            .I(N__42283));
    InMux I__8999 (
            .O(N__42298),
            .I(N__42280));
    Span4Mux_v I__8998 (
            .O(N__42295),
            .I(N__42277));
    Span4Mux_v I__8997 (
            .O(N__42292),
            .I(N__42274));
    Span4Mux_v I__8996 (
            .O(N__42289),
            .I(N__42269));
    Span4Mux_v I__8995 (
            .O(N__42286),
            .I(N__42269));
    Span4Mux_v I__8994 (
            .O(N__42283),
            .I(N__42266));
    LocalMux I__8993 (
            .O(N__42280),
            .I(un5_sdacdyn_cry_23_c_RNIELGZ0Z28));
    Odrv4 I__8992 (
            .O(N__42277),
            .I(un5_sdacdyn_cry_23_c_RNIELGZ0Z28));
    Odrv4 I__8991 (
            .O(N__42274),
            .I(un5_sdacdyn_cry_23_c_RNIELGZ0Z28));
    Odrv4 I__8990 (
            .O(N__42269),
            .I(un5_sdacdyn_cry_23_c_RNIELGZ0Z28));
    Odrv4 I__8989 (
            .O(N__42266),
            .I(un5_sdacdyn_cry_23_c_RNIELGZ0Z28));
    CascadeMux I__8988 (
            .O(N__42255),
            .I(sDAC_data_2_6_cascade_));
    InMux I__8987 (
            .O(N__42252),
            .I(N__42249));
    LocalMux I__8986 (
            .O(N__42249),
            .I(N__42246));
    Span4Mux_h I__8985 (
            .O(N__42246),
            .I(N__42243));
    Span4Mux_v I__8984 (
            .O(N__42243),
            .I(N__42240));
    Span4Mux_h I__8983 (
            .O(N__42240),
            .I(N__42237));
    Odrv4 I__8982 (
            .O(N__42237),
            .I(sDAC_dataZ0Z_6));
    CEMux I__8981 (
            .O(N__42234),
            .I(N__42192));
    CEMux I__8980 (
            .O(N__42233),
            .I(N__42192));
    CEMux I__8979 (
            .O(N__42232),
            .I(N__42192));
    CEMux I__8978 (
            .O(N__42231),
            .I(N__42192));
    CEMux I__8977 (
            .O(N__42230),
            .I(N__42192));
    CEMux I__8976 (
            .O(N__42229),
            .I(N__42192));
    CEMux I__8975 (
            .O(N__42228),
            .I(N__42192));
    CEMux I__8974 (
            .O(N__42227),
            .I(N__42192));
    CEMux I__8973 (
            .O(N__42226),
            .I(N__42192));
    CEMux I__8972 (
            .O(N__42225),
            .I(N__42192));
    CEMux I__8971 (
            .O(N__42224),
            .I(N__42192));
    CEMux I__8970 (
            .O(N__42223),
            .I(N__42192));
    CEMux I__8969 (
            .O(N__42222),
            .I(N__42192));
    CEMux I__8968 (
            .O(N__42221),
            .I(N__42192));
    GlobalMux I__8967 (
            .O(N__42192),
            .I(N__42189));
    gio2CtrlBuf I__8966 (
            .O(N__42189),
            .I(op_eq_scounterdac10_g));
    CascadeMux I__8965 (
            .O(N__42186),
            .I(N__42183));
    InMux I__8964 (
            .O(N__42183),
            .I(N__42180));
    LocalMux I__8963 (
            .O(N__42180),
            .I(N__42177));
    Span12Mux_v I__8962 (
            .O(N__42177),
            .I(N__42174));
    Odrv12 I__8961 (
            .O(N__42174),
            .I(sDAC_mem_2Z0Z_3));
    InMux I__8960 (
            .O(N__42171),
            .I(N__42168));
    LocalMux I__8959 (
            .O(N__42168),
            .I(N__42165));
    Span4Mux_v I__8958 (
            .O(N__42165),
            .I(N__42162));
    Odrv4 I__8957 (
            .O(N__42162),
            .I(sDAC_mem_34Z0Z_3));
    InMux I__8956 (
            .O(N__42159),
            .I(N__42156));
    LocalMux I__8955 (
            .O(N__42156),
            .I(N__42153));
    Span4Mux_h I__8954 (
            .O(N__42153),
            .I(N__42150));
    Odrv4 I__8953 (
            .O(N__42150),
            .I(sDAC_mem_33Z0Z_3));
    CascadeMux I__8952 (
            .O(N__42147),
            .I(sDAC_data_RNO_26Z0Z_6_cascade_));
    CascadeMux I__8951 (
            .O(N__42144),
            .I(N__42140));
    CascadeMux I__8950 (
            .O(N__42143),
            .I(N__42137));
    InMux I__8949 (
            .O(N__42140),
            .I(N__42132));
    InMux I__8948 (
            .O(N__42137),
            .I(N__42132));
    LocalMux I__8947 (
            .O(N__42132),
            .I(N__42129));
    Span4Mux_v I__8946 (
            .O(N__42129),
            .I(N__42126));
    Span4Mux_h I__8945 (
            .O(N__42126),
            .I(N__42123));
    Odrv4 I__8944 (
            .O(N__42123),
            .I(sDAC_mem_32Z0Z_3));
    InMux I__8943 (
            .O(N__42120),
            .I(N__42117));
    LocalMux I__8942 (
            .O(N__42117),
            .I(sDAC_data_RNO_27Z0Z_6));
    InMux I__8941 (
            .O(N__42114),
            .I(N__42108));
    InMux I__8940 (
            .O(N__42113),
            .I(N__42108));
    LocalMux I__8939 (
            .O(N__42108),
            .I(sDAC_mem_1Z0Z_3));
    InMux I__8938 (
            .O(N__42105),
            .I(N__42102));
    LocalMux I__8937 (
            .O(N__42102),
            .I(N__42099));
    Odrv12 I__8936 (
            .O(N__42099),
            .I(sDAC_mem_33Z0Z_4));
    CascadeMux I__8935 (
            .O(N__42096),
            .I(sDAC_data_RNO_26Z0Z_7_cascade_));
    CascadeMux I__8934 (
            .O(N__42093),
            .I(N__42090));
    InMux I__8933 (
            .O(N__42090),
            .I(N__42087));
    LocalMux I__8932 (
            .O(N__42087),
            .I(N__42084));
    Span4Mux_h I__8931 (
            .O(N__42084),
            .I(N__42081));
    Odrv4 I__8930 (
            .O(N__42081),
            .I(sDAC_data_RNO_14Z0Z_7));
    CascadeMux I__8929 (
            .O(N__42078),
            .I(N__42074));
    CascadeMux I__8928 (
            .O(N__42077),
            .I(N__42071));
    InMux I__8927 (
            .O(N__42074),
            .I(N__42066));
    InMux I__8926 (
            .O(N__42071),
            .I(N__42066));
    LocalMux I__8925 (
            .O(N__42066),
            .I(N__42063));
    Span4Mux_h I__8924 (
            .O(N__42063),
            .I(N__42060));
    Span4Mux_h I__8923 (
            .O(N__42060),
            .I(N__42057));
    Odrv4 I__8922 (
            .O(N__42057),
            .I(sDAC_mem_32Z0Z_4));
    InMux I__8921 (
            .O(N__42054),
            .I(N__42051));
    LocalMux I__8920 (
            .O(N__42051),
            .I(sDAC_data_RNO_27Z0Z_7));
    InMux I__8919 (
            .O(N__42048),
            .I(N__42042));
    InMux I__8918 (
            .O(N__42047),
            .I(N__42042));
    LocalMux I__8917 (
            .O(N__42042),
            .I(sDAC_mem_1Z0Z_4));
    CEMux I__8916 (
            .O(N__42039),
            .I(N__42036));
    LocalMux I__8915 (
            .O(N__42036),
            .I(N__42033));
    Span4Mux_h I__8914 (
            .O(N__42033),
            .I(N__42028));
    CEMux I__8913 (
            .O(N__42032),
            .I(N__42025));
    CEMux I__8912 (
            .O(N__42031),
            .I(N__42022));
    Odrv4 I__8911 (
            .O(N__42028),
            .I(sDAC_mem_1_1_sqmuxa));
    LocalMux I__8910 (
            .O(N__42025),
            .I(sDAC_mem_1_1_sqmuxa));
    LocalMux I__8909 (
            .O(N__42022),
            .I(sDAC_mem_1_1_sqmuxa));
    InMux I__8908 (
            .O(N__42015),
            .I(N__42012));
    LocalMux I__8907 (
            .O(N__42012),
            .I(sDAC_data_RNO_5Z0Z_6));
    InMux I__8906 (
            .O(N__42009),
            .I(N__42006));
    LocalMux I__8905 (
            .O(N__42006),
            .I(N__42003));
    Span4Mux_v I__8904 (
            .O(N__42003),
            .I(N__42000));
    Odrv4 I__8903 (
            .O(N__42000),
            .I(sDAC_data_RNO_4Z0Z_6));
    InMux I__8902 (
            .O(N__41997),
            .I(N__41994));
    LocalMux I__8901 (
            .O(N__41994),
            .I(N__41991));
    Span12Mux_v I__8900 (
            .O(N__41991),
            .I(N__41988));
    Odrv12 I__8899 (
            .O(N__41988),
            .I(sDAC_mem_40Z0Z_7));
    CEMux I__8898 (
            .O(N__41985),
            .I(N__41982));
    LocalMux I__8897 (
            .O(N__41982),
            .I(N__41979));
    Span4Mux_h I__8896 (
            .O(N__41979),
            .I(N__41976));
    Odrv4 I__8895 (
            .O(N__41976),
            .I(sDAC_mem_40_1_sqmuxa));
    InMux I__8894 (
            .O(N__41973),
            .I(N__41970));
    LocalMux I__8893 (
            .O(N__41970),
            .I(sDAC_mem_21Z0Z_0));
    InMux I__8892 (
            .O(N__41967),
            .I(N__41964));
    LocalMux I__8891 (
            .O(N__41964),
            .I(N__41961));
    Span4Mux_v I__8890 (
            .O(N__41961),
            .I(N__41958));
    Odrv4 I__8889 (
            .O(N__41958),
            .I(sDAC_data_RNO_20Z0Z_3));
    InMux I__8888 (
            .O(N__41955),
            .I(N__41952));
    LocalMux I__8887 (
            .O(N__41952),
            .I(sDAC_mem_20Z0Z_0));
    InMux I__8886 (
            .O(N__41949),
            .I(N__41946));
    LocalMux I__8885 (
            .O(N__41946),
            .I(sDAC_mem_21Z0Z_1));
    InMux I__8884 (
            .O(N__41943),
            .I(N__41940));
    LocalMux I__8883 (
            .O(N__41940),
            .I(N__41937));
    Span4Mux_v I__8882 (
            .O(N__41937),
            .I(N__41934));
    Odrv4 I__8881 (
            .O(N__41934),
            .I(sDAC_data_RNO_20Z0Z_4));
    InMux I__8880 (
            .O(N__41931),
            .I(N__41928));
    LocalMux I__8879 (
            .O(N__41928),
            .I(sDAC_mem_20Z0Z_1));
    InMux I__8878 (
            .O(N__41925),
            .I(N__41922));
    LocalMux I__8877 (
            .O(N__41922),
            .I(sDAC_mem_21Z0Z_2));
    InMux I__8876 (
            .O(N__41919),
            .I(N__41916));
    LocalMux I__8875 (
            .O(N__41916),
            .I(N__41913));
    Odrv12 I__8874 (
            .O(N__41913),
            .I(sDAC_data_RNO_20Z0Z_5));
    InMux I__8873 (
            .O(N__41910),
            .I(N__41907));
    LocalMux I__8872 (
            .O(N__41907),
            .I(sDAC_mem_20Z0Z_2));
    InMux I__8871 (
            .O(N__41904),
            .I(N__41901));
    LocalMux I__8870 (
            .O(N__41901),
            .I(N__41898));
    Odrv4 I__8869 (
            .O(N__41898),
            .I(sDAC_mem_21Z0Z_3));
    InMux I__8868 (
            .O(N__41895),
            .I(N__41892));
    LocalMux I__8867 (
            .O(N__41892),
            .I(sDAC_mem_20Z0Z_3));
    InMux I__8866 (
            .O(N__41889),
            .I(N__41886));
    LocalMux I__8865 (
            .O(N__41886),
            .I(N__41883));
    Odrv4 I__8864 (
            .O(N__41883),
            .I(sDAC_mem_38Z0Z_5));
    InMux I__8863 (
            .O(N__41880),
            .I(N__41877));
    LocalMux I__8862 (
            .O(N__41877),
            .I(N__41874));
    Span4Mux_v I__8861 (
            .O(N__41874),
            .I(N__41871));
    Odrv4 I__8860 (
            .O(N__41871),
            .I(sDAC_mem_38Z0Z_7));
    CEMux I__8859 (
            .O(N__41868),
            .I(N__41863));
    CEMux I__8858 (
            .O(N__41867),
            .I(N__41860));
    CEMux I__8857 (
            .O(N__41866),
            .I(N__41857));
    LocalMux I__8856 (
            .O(N__41863),
            .I(N__41854));
    LocalMux I__8855 (
            .O(N__41860),
            .I(N__41851));
    LocalMux I__8854 (
            .O(N__41857),
            .I(N__41848));
    Span4Mux_h I__8853 (
            .O(N__41854),
            .I(N__41845));
    Span4Mux_v I__8852 (
            .O(N__41851),
            .I(N__41842));
    Span4Mux_v I__8851 (
            .O(N__41848),
            .I(N__41839));
    Odrv4 I__8850 (
            .O(N__41845),
            .I(sDAC_mem_38_1_sqmuxa));
    Odrv4 I__8849 (
            .O(N__41842),
            .I(sDAC_mem_38_1_sqmuxa));
    Odrv4 I__8848 (
            .O(N__41839),
            .I(sDAC_mem_38_1_sqmuxa));
    InMux I__8847 (
            .O(N__41832),
            .I(N__41829));
    LocalMux I__8846 (
            .O(N__41829),
            .I(N__41826));
    Span4Mux_h I__8845 (
            .O(N__41826),
            .I(N__41823));
    Odrv4 I__8844 (
            .O(N__41823),
            .I(sDAC_mem_40Z0Z_2));
    InMux I__8843 (
            .O(N__41820),
            .I(N__41817));
    LocalMux I__8842 (
            .O(N__41817),
            .I(N__41814));
    Span4Mux_v I__8841 (
            .O(N__41814),
            .I(N__41811));
    Odrv4 I__8840 (
            .O(N__41811),
            .I(sDAC_mem_40Z0Z_3));
    InMux I__8839 (
            .O(N__41808),
            .I(N__41805));
    LocalMux I__8838 (
            .O(N__41805),
            .I(N__41802));
    Span4Mux_h I__8837 (
            .O(N__41802),
            .I(N__41799));
    Odrv4 I__8836 (
            .O(N__41799),
            .I(sDAC_mem_40Z0Z_4));
    InMux I__8835 (
            .O(N__41796),
            .I(N__41793));
    LocalMux I__8834 (
            .O(N__41793),
            .I(N__41790));
    Span4Mux_h I__8833 (
            .O(N__41790),
            .I(N__41787));
    Odrv4 I__8832 (
            .O(N__41787),
            .I(sDAC_mem_40Z0Z_6));
    InMux I__8831 (
            .O(N__41784),
            .I(N__41781));
    LocalMux I__8830 (
            .O(N__41781),
            .I(sDAC_mem_28Z0Z_7));
    CEMux I__8829 (
            .O(N__41778),
            .I(N__41773));
    CEMux I__8828 (
            .O(N__41777),
            .I(N__41769));
    CEMux I__8827 (
            .O(N__41776),
            .I(N__41766));
    LocalMux I__8826 (
            .O(N__41773),
            .I(N__41763));
    CEMux I__8825 (
            .O(N__41772),
            .I(N__41760));
    LocalMux I__8824 (
            .O(N__41769),
            .I(N__41757));
    LocalMux I__8823 (
            .O(N__41766),
            .I(N__41754));
    Span4Mux_v I__8822 (
            .O(N__41763),
            .I(N__41751));
    LocalMux I__8821 (
            .O(N__41760),
            .I(N__41748));
    Span4Mux_v I__8820 (
            .O(N__41757),
            .I(N__41745));
    Odrv4 I__8819 (
            .O(N__41754),
            .I(sDAC_mem_28_1_sqmuxa));
    Odrv4 I__8818 (
            .O(N__41751),
            .I(sDAC_mem_28_1_sqmuxa));
    Odrv4 I__8817 (
            .O(N__41748),
            .I(sDAC_mem_28_1_sqmuxa));
    Odrv4 I__8816 (
            .O(N__41745),
            .I(sDAC_mem_28_1_sqmuxa));
    InMux I__8815 (
            .O(N__41736),
            .I(N__41733));
    LocalMux I__8814 (
            .O(N__41733),
            .I(N__41730));
    Odrv4 I__8813 (
            .O(N__41730),
            .I(sDAC_mem_25Z0Z_1));
    CEMux I__8812 (
            .O(N__41727),
            .I(N__41724));
    LocalMux I__8811 (
            .O(N__41724),
            .I(N__41720));
    CEMux I__8810 (
            .O(N__41723),
            .I(N__41717));
    Span4Mux_v I__8809 (
            .O(N__41720),
            .I(N__41713));
    LocalMux I__8808 (
            .O(N__41717),
            .I(N__41710));
    CEMux I__8807 (
            .O(N__41716),
            .I(N__41707));
    Span4Mux_h I__8806 (
            .O(N__41713),
            .I(N__41702));
    Span4Mux_v I__8805 (
            .O(N__41710),
            .I(N__41702));
    LocalMux I__8804 (
            .O(N__41707),
            .I(N__41699));
    Odrv4 I__8803 (
            .O(N__41702),
            .I(sDAC_mem_25_1_sqmuxa));
    Odrv4 I__8802 (
            .O(N__41699),
            .I(sDAC_mem_25_1_sqmuxa));
    InMux I__8801 (
            .O(N__41694),
            .I(N__41691));
    LocalMux I__8800 (
            .O(N__41691),
            .I(N__41688));
    Span4Mux_v I__8799 (
            .O(N__41688),
            .I(N__41685));
    Span4Mux_h I__8798 (
            .O(N__41685),
            .I(N__41682));
    Span4Mux_v I__8797 (
            .O(N__41682),
            .I(N__41679));
    Odrv4 I__8796 (
            .O(N__41679),
            .I(sDAC_mem_17Z0Z_1));
    CascadeMux I__8795 (
            .O(N__41676),
            .I(N__41673));
    InMux I__8794 (
            .O(N__41673),
            .I(N__41670));
    LocalMux I__8793 (
            .O(N__41670),
            .I(N__41667));
    Span12Mux_s11_h I__8792 (
            .O(N__41667),
            .I(N__41664));
    Odrv12 I__8791 (
            .O(N__41664),
            .I(sDAC_data_RNO_29Z0Z_4));
    InMux I__8790 (
            .O(N__41661),
            .I(N__41658));
    LocalMux I__8789 (
            .O(N__41658),
            .I(N__41655));
    Span4Mux_v I__8788 (
            .O(N__41655),
            .I(N__41652));
    Span4Mux_h I__8787 (
            .O(N__41652),
            .I(N__41649));
    Odrv4 I__8786 (
            .O(N__41649),
            .I(sDAC_mem_38Z0Z_0));
    InMux I__8785 (
            .O(N__41646),
            .I(N__41643));
    LocalMux I__8784 (
            .O(N__41643),
            .I(N__41640));
    Span4Mux_h I__8783 (
            .O(N__41640),
            .I(N__41637));
    Odrv4 I__8782 (
            .O(N__41637),
            .I(sDAC_mem_38Z0Z_2));
    InMux I__8781 (
            .O(N__41634),
            .I(N__41631));
    LocalMux I__8780 (
            .O(N__41631),
            .I(N__41628));
    Odrv4 I__8779 (
            .O(N__41628),
            .I(sDAC_mem_38Z0Z_3));
    InMux I__8778 (
            .O(N__41625),
            .I(N__41622));
    LocalMux I__8777 (
            .O(N__41622),
            .I(N__41619));
    Span4Mux_h I__8776 (
            .O(N__41619),
            .I(N__41616));
    Odrv4 I__8775 (
            .O(N__41616),
            .I(sDAC_mem_38Z0Z_4));
    InMux I__8774 (
            .O(N__41613),
            .I(N__41610));
    LocalMux I__8773 (
            .O(N__41610),
            .I(sDAC_mem_28Z0Z_0));
    InMux I__8772 (
            .O(N__41607),
            .I(N__41604));
    LocalMux I__8771 (
            .O(N__41604),
            .I(N__41601));
    Span4Mux_h I__8770 (
            .O(N__41601),
            .I(N__41598));
    Odrv4 I__8769 (
            .O(N__41598),
            .I(sDAC_mem_24Z0Z_1));
    CascadeMux I__8768 (
            .O(N__41595),
            .I(sDAC_data_RNO_31Z0Z_4_cascade_));
    InMux I__8767 (
            .O(N__41592),
            .I(N__41589));
    LocalMux I__8766 (
            .O(N__41589),
            .I(sDAC_data_RNO_24Z0Z_4));
    CascadeMux I__8765 (
            .O(N__41586),
            .I(sDAC_data_2_39_ns_1_4_cascade_));
    InMux I__8764 (
            .O(N__41583),
            .I(N__41580));
    LocalMux I__8763 (
            .O(N__41580),
            .I(sDAC_data_RNO_23Z0Z_4));
    InMux I__8762 (
            .O(N__41577),
            .I(N__41574));
    LocalMux I__8761 (
            .O(N__41574),
            .I(N__41571));
    Odrv12 I__8760 (
            .O(N__41571),
            .I(sDAC_data_RNO_11Z0Z_4));
    InMux I__8759 (
            .O(N__41568),
            .I(N__41565));
    LocalMux I__8758 (
            .O(N__41565),
            .I(N__41562));
    Span4Mux_v I__8757 (
            .O(N__41562),
            .I(N__41559));
    Odrv4 I__8756 (
            .O(N__41559),
            .I(sDAC_mem_26Z0Z_1));
    InMux I__8755 (
            .O(N__41556),
            .I(N__41553));
    LocalMux I__8754 (
            .O(N__41553),
            .I(N__41550));
    Odrv4 I__8753 (
            .O(N__41550),
            .I(sDAC_mem_27Z0Z_1));
    InMux I__8752 (
            .O(N__41547),
            .I(N__41544));
    LocalMux I__8751 (
            .O(N__41544),
            .I(sDAC_data_RNO_32Z0Z_4));
    InMux I__8750 (
            .O(N__41541),
            .I(N__41538));
    LocalMux I__8749 (
            .O(N__41538),
            .I(sDAC_mem_28Z0Z_1));
    InMux I__8748 (
            .O(N__41535),
            .I(N__41532));
    LocalMux I__8747 (
            .O(N__41532),
            .I(N__41529));
    Span4Mux_h I__8746 (
            .O(N__41529),
            .I(N__41526));
    Odrv4 I__8745 (
            .O(N__41526),
            .I(sDAC_mem_28Z0Z_2));
    InMux I__8744 (
            .O(N__41523),
            .I(N__41520));
    LocalMux I__8743 (
            .O(N__41520),
            .I(N__41517));
    Span4Mux_v I__8742 (
            .O(N__41517),
            .I(N__41514));
    Odrv4 I__8741 (
            .O(N__41514),
            .I(sDAC_mem_28Z0Z_4));
    InMux I__8740 (
            .O(N__41511),
            .I(N__41508));
    LocalMux I__8739 (
            .O(N__41508),
            .I(N__41505));
    Span4Mux_h I__8738 (
            .O(N__41505),
            .I(N__41502));
    Odrv4 I__8737 (
            .O(N__41502),
            .I(sDAC_mem_28Z0Z_5));
    InMux I__8736 (
            .O(N__41499),
            .I(N__41496));
    LocalMux I__8735 (
            .O(N__41496),
            .I(N__41493));
    Span4Mux_h I__8734 (
            .O(N__41493),
            .I(N__41490));
    Odrv4 I__8733 (
            .O(N__41490),
            .I(sDAC_mem_27Z0Z_5));
    InMux I__8732 (
            .O(N__41487),
            .I(N__41484));
    LocalMux I__8731 (
            .O(N__41484),
            .I(N__41481));
    Span4Mux_v I__8730 (
            .O(N__41481),
            .I(N__41478));
    Span4Mux_h I__8729 (
            .O(N__41478),
            .I(N__41475));
    Odrv4 I__8728 (
            .O(N__41475),
            .I(sDAC_mem_27Z0Z_6));
    CascadeMux I__8727 (
            .O(N__41472),
            .I(N__41469));
    InMux I__8726 (
            .O(N__41469),
            .I(N__41466));
    LocalMux I__8725 (
            .O(N__41466),
            .I(N__41463));
    Odrv4 I__8724 (
            .O(N__41463),
            .I(sDAC_mem_27Z0Z_7));
    InMux I__8723 (
            .O(N__41460),
            .I(N__41457));
    LocalMux I__8722 (
            .O(N__41457),
            .I(N__41454));
    Odrv12 I__8721 (
            .O(N__41454),
            .I(sEEADC_freqZ0Z_0));
    InMux I__8720 (
            .O(N__41451),
            .I(N__41448));
    LocalMux I__8719 (
            .O(N__41448),
            .I(N__41445));
    Odrv12 I__8718 (
            .O(N__41445),
            .I(sEEADC_freqZ0Z_6));
    CascadeMux I__8717 (
            .O(N__41442),
            .I(N__41439));
    InMux I__8716 (
            .O(N__41439),
            .I(N__41436));
    LocalMux I__8715 (
            .O(N__41436),
            .I(N__41433));
    Span4Mux_h I__8714 (
            .O(N__41433),
            .I(N__41430));
    Odrv4 I__8713 (
            .O(N__41430),
            .I(sEEADC_freqZ0Z_7));
    InMux I__8712 (
            .O(N__41427),
            .I(N__41424));
    LocalMux I__8711 (
            .O(N__41424),
            .I(N__41421));
    Span4Mux_h I__8710 (
            .O(N__41421),
            .I(N__41418));
    Odrv4 I__8709 (
            .O(N__41418),
            .I(sDAC_mem_31Z0Z_0));
    InMux I__8708 (
            .O(N__41415),
            .I(N__41412));
    LocalMux I__8707 (
            .O(N__41412),
            .I(sDAC_mem_30Z0Z_0));
    InMux I__8706 (
            .O(N__41409),
            .I(N__41406));
    LocalMux I__8705 (
            .O(N__41406),
            .I(N__41403));
    Odrv4 I__8704 (
            .O(N__41403),
            .I(sDAC_mem_29Z0Z_0));
    InMux I__8703 (
            .O(N__41400),
            .I(N__41397));
    LocalMux I__8702 (
            .O(N__41397),
            .I(sDAC_data_RNO_24Z0Z_3));
    CascadeMux I__8701 (
            .O(N__41394),
            .I(sDAC_data_RNO_23Z0Z_3_cascade_));
    InMux I__8700 (
            .O(N__41391),
            .I(N__41388));
    LocalMux I__8699 (
            .O(N__41388),
            .I(sDAC_data_2_39_ns_1_3));
    InMux I__8698 (
            .O(N__41385),
            .I(N__41382));
    LocalMux I__8697 (
            .O(N__41382),
            .I(N__41379));
    Span4Mux_h I__8696 (
            .O(N__41379),
            .I(N__41376));
    Odrv4 I__8695 (
            .O(N__41376),
            .I(sDAC_data_RNO_11Z0Z_3));
    CascadeMux I__8694 (
            .O(N__41373),
            .I(sDAC_data_2_3_cascade_));
    InMux I__8693 (
            .O(N__41370),
            .I(N__41367));
    LocalMux I__8692 (
            .O(N__41367),
            .I(N__41364));
    Span4Mux_v I__8691 (
            .O(N__41364),
            .I(N__41361));
    Span4Mux_h I__8690 (
            .O(N__41361),
            .I(N__41358));
    Span4Mux_v I__8689 (
            .O(N__41358),
            .I(N__41355));
    Odrv4 I__8688 (
            .O(N__41355),
            .I(sDAC_dataZ0Z_3));
    InMux I__8687 (
            .O(N__41352),
            .I(N__41349));
    LocalMux I__8686 (
            .O(N__41349),
            .I(N__41346));
    Span4Mux_v I__8685 (
            .O(N__41346),
            .I(N__41343));
    Span4Mux_h I__8684 (
            .O(N__41343),
            .I(N__41340));
    Odrv4 I__8683 (
            .O(N__41340),
            .I(sDAC_mem_16Z0Z_7));
    InMux I__8682 (
            .O(N__41337),
            .I(N__41334));
    LocalMux I__8681 (
            .O(N__41334),
            .I(N__41331));
    Span4Mux_h I__8680 (
            .O(N__41331),
            .I(N__41328));
    Span4Mux_v I__8679 (
            .O(N__41328),
            .I(N__41325));
    Odrv4 I__8678 (
            .O(N__41325),
            .I(sDAC_mem_17Z0Z_7));
    InMux I__8677 (
            .O(N__41322),
            .I(N__41319));
    LocalMux I__8676 (
            .O(N__41319),
            .I(sDAC_data_RNO_29Z0Z_10));
    InMux I__8675 (
            .O(N__41316),
            .I(N__41313));
    LocalMux I__8674 (
            .O(N__41313),
            .I(N__41310));
    Span4Mux_h I__8673 (
            .O(N__41310),
            .I(N__41307));
    Odrv4 I__8672 (
            .O(N__41307),
            .I(sDAC_mem_19Z0Z_3));
    InMux I__8671 (
            .O(N__41304),
            .I(N__41301));
    LocalMux I__8670 (
            .O(N__41301),
            .I(N__41298));
    Odrv12 I__8669 (
            .O(N__41298),
            .I(sDAC_mem_18Z0Z_3));
    InMux I__8668 (
            .O(N__41295),
            .I(N__41292));
    LocalMux I__8667 (
            .O(N__41292),
            .I(N__41289));
    Span4Mux_v I__8666 (
            .O(N__41289),
            .I(N__41286));
    Span4Mux_h I__8665 (
            .O(N__41286),
            .I(N__41283));
    Odrv4 I__8664 (
            .O(N__41283),
            .I(sDAC_mem_23Z0Z_1));
    InMux I__8663 (
            .O(N__41280),
            .I(N__41277));
    LocalMux I__8662 (
            .O(N__41277),
            .I(N__41274));
    Span4Mux_h I__8661 (
            .O(N__41274),
            .I(N__41271));
    Span4Mux_v I__8660 (
            .O(N__41271),
            .I(N__41268));
    Odrv4 I__8659 (
            .O(N__41268),
            .I(sDAC_mem_22Z0Z_1));
    InMux I__8658 (
            .O(N__41265),
            .I(N__41262));
    LocalMux I__8657 (
            .O(N__41262),
            .I(N__41259));
    Odrv12 I__8656 (
            .O(N__41259),
            .I(sDAC_data_RNO_21Z0Z_4));
    InMux I__8655 (
            .O(N__41256),
            .I(N__41253));
    LocalMux I__8654 (
            .O(N__41253),
            .I(N__41250));
    Span4Mux_v I__8653 (
            .O(N__41250),
            .I(N__41247));
    Span4Mux_h I__8652 (
            .O(N__41247),
            .I(N__41244));
    Odrv4 I__8651 (
            .O(N__41244),
            .I(sDAC_mem_27Z0Z_2));
    InMux I__8650 (
            .O(N__41241),
            .I(N__41238));
    LocalMux I__8649 (
            .O(N__41238),
            .I(N__41235));
    Span4Mux_h I__8648 (
            .O(N__41235),
            .I(N__41232));
    Span4Mux_v I__8647 (
            .O(N__41232),
            .I(N__41229));
    Odrv4 I__8646 (
            .O(N__41229),
            .I(sDAC_mem_27Z0Z_3));
    InMux I__8645 (
            .O(N__41226),
            .I(N__41223));
    LocalMux I__8644 (
            .O(N__41223),
            .I(N__41220));
    Span4Mux_h I__8643 (
            .O(N__41220),
            .I(N__41217));
    Odrv4 I__8642 (
            .O(N__41217),
            .I(sDAC_mem_27Z0Z_4));
    CascadeMux I__8641 (
            .O(N__41214),
            .I(sDAC_data_RNO_1Z0Z_4_cascade_));
    InMux I__8640 (
            .O(N__41211),
            .I(N__41208));
    LocalMux I__8639 (
            .O(N__41208),
            .I(sDAC_data_2_41_ns_1_4));
    CascadeMux I__8638 (
            .O(N__41205),
            .I(sDAC_data_2_4_cascade_));
    InMux I__8637 (
            .O(N__41202),
            .I(N__41199));
    LocalMux I__8636 (
            .O(N__41199),
            .I(N__41196));
    Span12Mux_h I__8635 (
            .O(N__41196),
            .I(N__41193));
    Odrv12 I__8634 (
            .O(N__41193),
            .I(sDAC_dataZ0Z_4));
    InMux I__8633 (
            .O(N__41190),
            .I(N__41187));
    LocalMux I__8632 (
            .O(N__41187),
            .I(N__41184));
    Span4Mux_v I__8631 (
            .O(N__41184),
            .I(N__41181));
    Odrv4 I__8630 (
            .O(N__41181),
            .I(sDAC_data_RNO_21Z0Z_3));
    CascadeMux I__8629 (
            .O(N__41178),
            .I(sDAC_data_RNO_10Z0Z_3_cascade_));
    InMux I__8628 (
            .O(N__41175),
            .I(N__41172));
    LocalMux I__8627 (
            .O(N__41172),
            .I(N__41169));
    Odrv4 I__8626 (
            .O(N__41169),
            .I(sDAC_data_RNO_30Z0Z_3));
    InMux I__8625 (
            .O(N__41166),
            .I(N__41163));
    LocalMux I__8624 (
            .O(N__41163),
            .I(sDAC_data_2_32_ns_1_3));
    CascadeMux I__8623 (
            .O(N__41160),
            .I(N__41157));
    InMux I__8622 (
            .O(N__41157),
            .I(N__41154));
    LocalMux I__8621 (
            .O(N__41154),
            .I(N__41151));
    Span4Mux_h I__8620 (
            .O(N__41151),
            .I(N__41148));
    Sp12to4 I__8619 (
            .O(N__41148),
            .I(N__41145));
    Odrv12 I__8618 (
            .O(N__41145),
            .I(sDAC_data_RNO_15Z0Z_3));
    InMux I__8617 (
            .O(N__41142),
            .I(N__41139));
    LocalMux I__8616 (
            .O(N__41139),
            .I(sDAC_data_RNO_14Z0Z_3));
    InMux I__8615 (
            .O(N__41136),
            .I(N__41133));
    LocalMux I__8614 (
            .O(N__41133),
            .I(N__41130));
    Span4Mux_v I__8613 (
            .O(N__41130),
            .I(N__41127));
    Span4Mux_v I__8612 (
            .O(N__41127),
            .I(N__41124));
    Odrv4 I__8611 (
            .O(N__41124),
            .I(sDAC_data_RNO_5Z0Z_3));
    CascadeMux I__8610 (
            .O(N__41121),
            .I(sDAC_data_2_14_ns_1_3_cascade_));
    InMux I__8609 (
            .O(N__41118),
            .I(N__41115));
    LocalMux I__8608 (
            .O(N__41115),
            .I(sDAC_data_RNO_4Z0Z_3));
    CascadeMux I__8607 (
            .O(N__41112),
            .I(sDAC_data_RNO_1Z0Z_3_cascade_));
    InMux I__8606 (
            .O(N__41109),
            .I(N__41106));
    LocalMux I__8605 (
            .O(N__41106),
            .I(sDAC_data_2_41_ns_1_3));
    CascadeMux I__8604 (
            .O(N__41103),
            .I(sDAC_data_RNO_17Z0Z_6_cascade_));
    InMux I__8603 (
            .O(N__41100),
            .I(N__41097));
    LocalMux I__8602 (
            .O(N__41097),
            .I(N__41094));
    Span4Mux_v I__8601 (
            .O(N__41094),
            .I(N__41091));
    Odrv4 I__8600 (
            .O(N__41091),
            .I(sDAC_mem_8Z0Z_3));
    CascadeMux I__8599 (
            .O(N__41088),
            .I(sDAC_data_2_20_am_1_6_cascade_));
    InMux I__8598 (
            .O(N__41085),
            .I(N__41082));
    LocalMux I__8597 (
            .O(N__41082),
            .I(N__41079));
    Span4Mux_v I__8596 (
            .O(N__41079),
            .I(N__41076));
    Odrv4 I__8595 (
            .O(N__41076),
            .I(sDAC_data_2_24_ns_1_6));
    CascadeMux I__8594 (
            .O(N__41073),
            .I(sDAC_data_RNO_7Z0Z_6_cascade_));
    InMux I__8593 (
            .O(N__41070),
            .I(N__41067));
    LocalMux I__8592 (
            .O(N__41067),
            .I(sDAC_data_RNO_8Z0Z_6));
    CascadeMux I__8591 (
            .O(N__41064),
            .I(sDAC_data_RNO_10Z0Z_4_cascade_));
    InMux I__8590 (
            .O(N__41061),
            .I(N__41058));
    LocalMux I__8589 (
            .O(N__41058),
            .I(N__41055));
    Span4Mux_h I__8588 (
            .O(N__41055),
            .I(N__41052));
    Odrv4 I__8587 (
            .O(N__41052),
            .I(sDAC_data_RNO_30Z0Z_4));
    InMux I__8586 (
            .O(N__41049),
            .I(N__41046));
    LocalMux I__8585 (
            .O(N__41046),
            .I(sDAC_data_2_32_ns_1_4));
    CascadeMux I__8584 (
            .O(N__41043),
            .I(N__41040));
    InMux I__8583 (
            .O(N__41040),
            .I(N__41037));
    LocalMux I__8582 (
            .O(N__41037),
            .I(N__41034));
    Odrv12 I__8581 (
            .O(N__41034),
            .I(sDAC_data_RNO_15Z0Z_4));
    InMux I__8580 (
            .O(N__41031),
            .I(N__41028));
    LocalMux I__8579 (
            .O(N__41028),
            .I(N__41025));
    Span4Mux_v I__8578 (
            .O(N__41025),
            .I(N__41022));
    Odrv4 I__8577 (
            .O(N__41022),
            .I(sDAC_data_RNO_14Z0Z_4));
    InMux I__8576 (
            .O(N__41019),
            .I(N__41016));
    LocalMux I__8575 (
            .O(N__41016),
            .I(N__41013));
    Span4Mux_h I__8574 (
            .O(N__41013),
            .I(N__41010));
    Span4Mux_v I__8573 (
            .O(N__41010),
            .I(N__41007));
    Odrv4 I__8572 (
            .O(N__41007),
            .I(sDAC_data_RNO_5Z0Z_4));
    CascadeMux I__8571 (
            .O(N__41004),
            .I(sDAC_data_2_14_ns_1_4_cascade_));
    InMux I__8570 (
            .O(N__41001),
            .I(N__40998));
    LocalMux I__8569 (
            .O(N__40998),
            .I(N__40995));
    Span4Mux_h I__8568 (
            .O(N__40995),
            .I(N__40992));
    Odrv4 I__8567 (
            .O(N__40992),
            .I(sDAC_data_RNO_4Z0Z_4));
    CascadeMux I__8566 (
            .O(N__40989),
            .I(N__40986));
    InMux I__8565 (
            .O(N__40986),
            .I(N__40983));
    LocalMux I__8564 (
            .O(N__40983),
            .I(N__40980));
    Odrv4 I__8563 (
            .O(N__40980),
            .I(sDAC_data_RNO_15Z0Z_8));
    InMux I__8562 (
            .O(N__40977),
            .I(N__40974));
    LocalMux I__8561 (
            .O(N__40974),
            .I(N__40971));
    Odrv4 I__8560 (
            .O(N__40971),
            .I(sDAC_data_RNO_14Z0Z_8));
    InMux I__8559 (
            .O(N__40968),
            .I(N__40965));
    LocalMux I__8558 (
            .O(N__40965),
            .I(sDAC_data_RNO_5Z0Z_8));
    CascadeMux I__8557 (
            .O(N__40962),
            .I(sDAC_data_2_14_ns_1_8_cascade_));
    InMux I__8556 (
            .O(N__40959),
            .I(N__40956));
    LocalMux I__8555 (
            .O(N__40956),
            .I(sDAC_data_RNO_4Z0Z_8));
    InMux I__8554 (
            .O(N__40953),
            .I(N__40950));
    LocalMux I__8553 (
            .O(N__40950),
            .I(sDAC_data_RNO_10Z0Z_8));
    CascadeMux I__8552 (
            .O(N__40947),
            .I(N__40944));
    InMux I__8551 (
            .O(N__40944),
            .I(N__40941));
    LocalMux I__8550 (
            .O(N__40941),
            .I(N__40938));
    Span4Mux_h I__8549 (
            .O(N__40938),
            .I(N__40935));
    Span4Mux_h I__8548 (
            .O(N__40935),
            .I(N__40932));
    Odrv4 I__8547 (
            .O(N__40932),
            .I(sDAC_data_RNO_11Z0Z_8));
    CascadeMux I__8546 (
            .O(N__40929),
            .I(sDAC_data_2_41_ns_1_8_cascade_));
    InMux I__8545 (
            .O(N__40926),
            .I(N__40923));
    LocalMux I__8544 (
            .O(N__40923),
            .I(sDAC_data_RNO_1Z0Z_8));
    CascadeMux I__8543 (
            .O(N__40920),
            .I(sDAC_data_2_8_cascade_));
    InMux I__8542 (
            .O(N__40917),
            .I(N__40914));
    LocalMux I__8541 (
            .O(N__40914),
            .I(N__40911));
    Span4Mux_h I__8540 (
            .O(N__40911),
            .I(N__40908));
    Span4Mux_h I__8539 (
            .O(N__40908),
            .I(N__40905));
    Sp12to4 I__8538 (
            .O(N__40905),
            .I(N__40902));
    Odrv12 I__8537 (
            .O(N__40902),
            .I(sDAC_dataZ0Z_8));
    CascadeMux I__8536 (
            .O(N__40899),
            .I(N__40896));
    InMux I__8535 (
            .O(N__40896),
            .I(N__40893));
    LocalMux I__8534 (
            .O(N__40893),
            .I(N__40890));
    Span4Mux_v I__8533 (
            .O(N__40890),
            .I(N__40887));
    Odrv4 I__8532 (
            .O(N__40887),
            .I(sDAC_mem_2Z0Z_1));
    InMux I__8531 (
            .O(N__40884),
            .I(N__40881));
    LocalMux I__8530 (
            .O(N__40881),
            .I(N__40878));
    Odrv12 I__8529 (
            .O(N__40878),
            .I(sDAC_mem_34Z0Z_1));
    InMux I__8528 (
            .O(N__40875),
            .I(N__40872));
    LocalMux I__8527 (
            .O(N__40872),
            .I(N__40869));
    Odrv12 I__8526 (
            .O(N__40869),
            .I(sDAC_mem_35Z0Z_1));
    CascadeMux I__8525 (
            .O(N__40866),
            .I(sDAC_data_2_6_bm_1_4_cascade_));
    InMux I__8524 (
            .O(N__40863),
            .I(N__40860));
    LocalMux I__8523 (
            .O(N__40860),
            .I(sDAC_mem_3Z0Z_1));
    InMux I__8522 (
            .O(N__40857),
            .I(N__40854));
    LocalMux I__8521 (
            .O(N__40854),
            .I(N__40851));
    Span4Mux_v I__8520 (
            .O(N__40851),
            .I(N__40848));
    Odrv4 I__8519 (
            .O(N__40848),
            .I(sDAC_mem_7Z0Z_3));
    CascadeMux I__8518 (
            .O(N__40845),
            .I(sDAC_data_2_13_bm_1_6_cascade_));
    InMux I__8517 (
            .O(N__40842),
            .I(N__40839));
    LocalMux I__8516 (
            .O(N__40839),
            .I(N__40836));
    Span4Mux_v I__8515 (
            .O(N__40836),
            .I(N__40833));
    Odrv4 I__8514 (
            .O(N__40833),
            .I(sDAC_mem_39Z0Z_3));
    InMux I__8513 (
            .O(N__40830),
            .I(N__40827));
    LocalMux I__8512 (
            .O(N__40827),
            .I(sDAC_mem_6Z0Z_3));
    InMux I__8511 (
            .O(N__40824),
            .I(N__40821));
    LocalMux I__8510 (
            .O(N__40821),
            .I(sDAC_mem_6Z0Z_4));
    InMux I__8509 (
            .O(N__40818),
            .I(N__40815));
    LocalMux I__8508 (
            .O(N__40815),
            .I(N__40812));
    Span4Mux_v I__8507 (
            .O(N__40812),
            .I(N__40809));
    Odrv4 I__8506 (
            .O(N__40809),
            .I(sDAC_mem_6Z0Z_5));
    InMux I__8505 (
            .O(N__40806),
            .I(N__40803));
    LocalMux I__8504 (
            .O(N__40803),
            .I(N__40800));
    Span4Mux_v I__8503 (
            .O(N__40800),
            .I(N__40797));
    Odrv4 I__8502 (
            .O(N__40797),
            .I(sDAC_mem_7Z0Z_5));
    CascadeMux I__8501 (
            .O(N__40794),
            .I(sDAC_data_2_13_bm_1_8_cascade_));
    InMux I__8500 (
            .O(N__40791),
            .I(N__40788));
    LocalMux I__8499 (
            .O(N__40788),
            .I(N__40785));
    Span4Mux_v I__8498 (
            .O(N__40785),
            .I(N__40782));
    Odrv4 I__8497 (
            .O(N__40782),
            .I(sDAC_mem_39Z0Z_5));
    InMux I__8496 (
            .O(N__40779),
            .I(N__40776));
    LocalMux I__8495 (
            .O(N__40776),
            .I(N__40773));
    Span4Mux_v I__8494 (
            .O(N__40773),
            .I(N__40770));
    Odrv4 I__8493 (
            .O(N__40770),
            .I(sDAC_data_RNO_21Z0Z_8));
    InMux I__8492 (
            .O(N__40767),
            .I(N__40764));
    LocalMux I__8491 (
            .O(N__40764),
            .I(N__40761));
    Odrv4 I__8490 (
            .O(N__40761),
            .I(sDAC_data_RNO_20Z0Z_8));
    CascadeMux I__8489 (
            .O(N__40758),
            .I(N__40755));
    InMux I__8488 (
            .O(N__40755),
            .I(N__40752));
    LocalMux I__8487 (
            .O(N__40752),
            .I(N__40749));
    Odrv12 I__8486 (
            .O(N__40749),
            .I(sDAC_data_RNO_29Z0Z_8));
    InMux I__8485 (
            .O(N__40746),
            .I(N__40743));
    LocalMux I__8484 (
            .O(N__40743),
            .I(N__40740));
    Span4Mux_h I__8483 (
            .O(N__40740),
            .I(N__40737));
    Odrv4 I__8482 (
            .O(N__40737),
            .I(sDAC_data_RNO_30Z0Z_8));
    CascadeMux I__8481 (
            .O(N__40734),
            .I(N__40731));
    InMux I__8480 (
            .O(N__40731),
            .I(N__40728));
    LocalMux I__8479 (
            .O(N__40728),
            .I(N__40725));
    Odrv4 I__8478 (
            .O(N__40725),
            .I(sDAC_data_2_32_ns_1_8));
    InMux I__8477 (
            .O(N__40722),
            .I(N__40719));
    LocalMux I__8476 (
            .O(N__40719),
            .I(N__40716));
    Span4Mux_v I__8475 (
            .O(N__40716),
            .I(N__40713));
    Odrv4 I__8474 (
            .O(N__40713),
            .I(sDAC_mem_35Z0Z_6));
    CEMux I__8473 (
            .O(N__40710),
            .I(N__40707));
    LocalMux I__8472 (
            .O(N__40707),
            .I(sDAC_mem_35_1_sqmuxa));
    InMux I__8471 (
            .O(N__40704),
            .I(N__40701));
    LocalMux I__8470 (
            .O(N__40701),
            .I(sDAC_mem_21Z0Z_4));
    InMux I__8469 (
            .O(N__40698),
            .I(N__40695));
    LocalMux I__8468 (
            .O(N__40695),
            .I(sDAC_mem_21Z0Z_5));
    InMux I__8467 (
            .O(N__40692),
            .I(N__40689));
    LocalMux I__8466 (
            .O(N__40689),
            .I(sDAC_mem_21Z0Z_6));
    InMux I__8465 (
            .O(N__40686),
            .I(N__40683));
    LocalMux I__8464 (
            .O(N__40683),
            .I(N__40680));
    Span4Mux_v I__8463 (
            .O(N__40680),
            .I(N__40677));
    Odrv4 I__8462 (
            .O(N__40677),
            .I(sDAC_mem_21Z0Z_7));
    CEMux I__8461 (
            .O(N__40674),
            .I(N__40671));
    LocalMux I__8460 (
            .O(N__40671),
            .I(N__40668));
    Span4Mux_h I__8459 (
            .O(N__40668),
            .I(N__40665));
    Span4Mux_v I__8458 (
            .O(N__40665),
            .I(N__40662));
    Span4Mux_h I__8457 (
            .O(N__40662),
            .I(N__40659));
    Odrv4 I__8456 (
            .O(N__40659),
            .I(sDAC_mem_21_1_sqmuxa));
    CEMux I__8455 (
            .O(N__40656),
            .I(N__40653));
    LocalMux I__8454 (
            .O(N__40653),
            .I(N__40650));
    Span4Mux_h I__8453 (
            .O(N__40650),
            .I(N__40647));
    Span4Mux_h I__8452 (
            .O(N__40647),
            .I(N__40644));
    Odrv4 I__8451 (
            .O(N__40644),
            .I(sDAC_mem_36_1_sqmuxa));
    InMux I__8450 (
            .O(N__40641),
            .I(N__40638));
    LocalMux I__8449 (
            .O(N__40638),
            .I(N__40630));
    InMux I__8448 (
            .O(N__40637),
            .I(N__40619));
    InMux I__8447 (
            .O(N__40636),
            .I(N__40619));
    InMux I__8446 (
            .O(N__40635),
            .I(N__40619));
    InMux I__8445 (
            .O(N__40634),
            .I(N__40619));
    InMux I__8444 (
            .O(N__40633),
            .I(N__40619));
    Odrv4 I__8443 (
            .O(N__40630),
            .I(N_288));
    LocalMux I__8442 (
            .O(N__40619),
            .I(N_288));
    CascadeMux I__8441 (
            .O(N__40614),
            .I(N__40605));
    InMux I__8440 (
            .O(N__40613),
            .I(N__40600));
    InMux I__8439 (
            .O(N__40612),
            .I(N__40587));
    InMux I__8438 (
            .O(N__40611),
            .I(N__40587));
    InMux I__8437 (
            .O(N__40610),
            .I(N__40587));
    InMux I__8436 (
            .O(N__40609),
            .I(N__40587));
    InMux I__8435 (
            .O(N__40608),
            .I(N__40587));
    InMux I__8434 (
            .O(N__40605),
            .I(N__40587));
    CascadeMux I__8433 (
            .O(N__40604),
            .I(N__40579));
    CascadeMux I__8432 (
            .O(N__40603),
            .I(N__40576));
    LocalMux I__8431 (
            .O(N__40600),
            .I(N__40572));
    LocalMux I__8430 (
            .O(N__40587),
            .I(N__40569));
    InMux I__8429 (
            .O(N__40586),
            .I(N__40556));
    InMux I__8428 (
            .O(N__40585),
            .I(N__40556));
    InMux I__8427 (
            .O(N__40584),
            .I(N__40556));
    InMux I__8426 (
            .O(N__40583),
            .I(N__40556));
    InMux I__8425 (
            .O(N__40582),
            .I(N__40556));
    InMux I__8424 (
            .O(N__40579),
            .I(N__40556));
    InMux I__8423 (
            .O(N__40576),
            .I(N__40552));
    InMux I__8422 (
            .O(N__40575),
            .I(N__40549));
    Span4Mux_v I__8421 (
            .O(N__40572),
            .I(N__40542));
    Span4Mux_h I__8420 (
            .O(N__40569),
            .I(N__40542));
    LocalMux I__8419 (
            .O(N__40556),
            .I(N__40542));
    CascadeMux I__8418 (
            .O(N__40555),
            .I(N__40535));
    LocalMux I__8417 (
            .O(N__40552),
            .I(N__40526));
    LocalMux I__8416 (
            .O(N__40549),
            .I(N__40526));
    Span4Mux_v I__8415 (
            .O(N__40542),
            .I(N__40523));
    InMux I__8414 (
            .O(N__40541),
            .I(N__40520));
    CascadeMux I__8413 (
            .O(N__40540),
            .I(N__40513));
    CascadeMux I__8412 (
            .O(N__40539),
            .I(N__40508));
    CascadeMux I__8411 (
            .O(N__40538),
            .I(N__40505));
    InMux I__8410 (
            .O(N__40535),
            .I(N__40502));
    InMux I__8409 (
            .O(N__40534),
            .I(N__40499));
    CascadeMux I__8408 (
            .O(N__40533),
            .I(N__40496));
    InMux I__8407 (
            .O(N__40532),
            .I(N__40490));
    InMux I__8406 (
            .O(N__40531),
            .I(N__40490));
    Span4Mux_v I__8405 (
            .O(N__40526),
            .I(N__40485));
    Span4Mux_h I__8404 (
            .O(N__40523),
            .I(N__40485));
    LocalMux I__8403 (
            .O(N__40520),
            .I(N__40482));
    InMux I__8402 (
            .O(N__40519),
            .I(N__40479));
    InMux I__8401 (
            .O(N__40518),
            .I(N__40472));
    InMux I__8400 (
            .O(N__40517),
            .I(N__40472));
    InMux I__8399 (
            .O(N__40516),
            .I(N__40472));
    InMux I__8398 (
            .O(N__40513),
            .I(N__40465));
    InMux I__8397 (
            .O(N__40512),
            .I(N__40465));
    InMux I__8396 (
            .O(N__40511),
            .I(N__40465));
    InMux I__8395 (
            .O(N__40508),
            .I(N__40462));
    InMux I__8394 (
            .O(N__40505),
            .I(N__40459));
    LocalMux I__8393 (
            .O(N__40502),
            .I(N__40454));
    LocalMux I__8392 (
            .O(N__40499),
            .I(N__40454));
    InMux I__8391 (
            .O(N__40496),
            .I(N__40449));
    InMux I__8390 (
            .O(N__40495),
            .I(N__40449));
    LocalMux I__8389 (
            .O(N__40490),
            .I(N__40444));
    Span4Mux_h I__8388 (
            .O(N__40485),
            .I(N__40444));
    Span4Mux_h I__8387 (
            .O(N__40482),
            .I(N__40441));
    LocalMux I__8386 (
            .O(N__40479),
            .I(sAddressZ0Z_3));
    LocalMux I__8385 (
            .O(N__40472),
            .I(sAddressZ0Z_3));
    LocalMux I__8384 (
            .O(N__40465),
            .I(sAddressZ0Z_3));
    LocalMux I__8383 (
            .O(N__40462),
            .I(sAddressZ0Z_3));
    LocalMux I__8382 (
            .O(N__40459),
            .I(sAddressZ0Z_3));
    Odrv4 I__8381 (
            .O(N__40454),
            .I(sAddressZ0Z_3));
    LocalMux I__8380 (
            .O(N__40449),
            .I(sAddressZ0Z_3));
    Odrv4 I__8379 (
            .O(N__40444),
            .I(sAddressZ0Z_3));
    Odrv4 I__8378 (
            .O(N__40441),
            .I(sAddressZ0Z_3));
    CascadeMux I__8377 (
            .O(N__40422),
            .I(N_288_cascade_));
    CascadeMux I__8376 (
            .O(N__40419),
            .I(N__40413));
    CascadeMux I__8375 (
            .O(N__40418),
            .I(N__40409));
    InMux I__8374 (
            .O(N__40417),
            .I(N__40403));
    InMux I__8373 (
            .O(N__40416),
            .I(N__40392));
    InMux I__8372 (
            .O(N__40413),
            .I(N__40379));
    InMux I__8371 (
            .O(N__40412),
            .I(N__40379));
    InMux I__8370 (
            .O(N__40409),
            .I(N__40379));
    InMux I__8369 (
            .O(N__40408),
            .I(N__40379));
    InMux I__8368 (
            .O(N__40407),
            .I(N__40379));
    InMux I__8367 (
            .O(N__40406),
            .I(N__40379));
    LocalMux I__8366 (
            .O(N__40403),
            .I(N__40376));
    InMux I__8365 (
            .O(N__40402),
            .I(N__40367));
    InMux I__8364 (
            .O(N__40401),
            .I(N__40367));
    InMux I__8363 (
            .O(N__40400),
            .I(N__40367));
    InMux I__8362 (
            .O(N__40399),
            .I(N__40367));
    InMux I__8361 (
            .O(N__40398),
            .I(N__40360));
    InMux I__8360 (
            .O(N__40397),
            .I(N__40360));
    InMux I__8359 (
            .O(N__40396),
            .I(N__40360));
    InMux I__8358 (
            .O(N__40395),
            .I(N__40356));
    LocalMux I__8357 (
            .O(N__40392),
            .I(N__40352));
    LocalMux I__8356 (
            .O(N__40379),
            .I(N__40349));
    Span4Mux_v I__8355 (
            .O(N__40376),
            .I(N__40340));
    LocalMux I__8354 (
            .O(N__40367),
            .I(N__40340));
    LocalMux I__8353 (
            .O(N__40360),
            .I(N__40340));
    InMux I__8352 (
            .O(N__40359),
            .I(N__40337));
    LocalMux I__8351 (
            .O(N__40356),
            .I(N__40330));
    CascadeMux I__8350 (
            .O(N__40355),
            .I(N__40320));
    Span4Mux_v I__8349 (
            .O(N__40352),
            .I(N__40315));
    Span4Mux_v I__8348 (
            .O(N__40349),
            .I(N__40315));
    InMux I__8347 (
            .O(N__40348),
            .I(N__40310));
    InMux I__8346 (
            .O(N__40347),
            .I(N__40310));
    Span4Mux_h I__8345 (
            .O(N__40340),
            .I(N__40307));
    LocalMux I__8344 (
            .O(N__40337),
            .I(N__40301));
    InMux I__8343 (
            .O(N__40336),
            .I(N__40296));
    InMux I__8342 (
            .O(N__40335),
            .I(N__40296));
    InMux I__8341 (
            .O(N__40334),
            .I(N__40291));
    InMux I__8340 (
            .O(N__40333),
            .I(N__40291));
    Span4Mux_h I__8339 (
            .O(N__40330),
            .I(N__40288));
    InMux I__8338 (
            .O(N__40329),
            .I(N__40283));
    InMux I__8337 (
            .O(N__40328),
            .I(N__40283));
    InMux I__8336 (
            .O(N__40327),
            .I(N__40278));
    InMux I__8335 (
            .O(N__40326),
            .I(N__40278));
    InMux I__8334 (
            .O(N__40325),
            .I(N__40269));
    InMux I__8333 (
            .O(N__40324),
            .I(N__40269));
    InMux I__8332 (
            .O(N__40323),
            .I(N__40269));
    InMux I__8331 (
            .O(N__40320),
            .I(N__40269));
    Span4Mux_h I__8330 (
            .O(N__40315),
            .I(N__40264));
    LocalMux I__8329 (
            .O(N__40310),
            .I(N__40264));
    Span4Mux_v I__8328 (
            .O(N__40307),
            .I(N__40261));
    InMux I__8327 (
            .O(N__40306),
            .I(N__40254));
    InMux I__8326 (
            .O(N__40305),
            .I(N__40254));
    InMux I__8325 (
            .O(N__40304),
            .I(N__40254));
    Span12Mux_h I__8324 (
            .O(N__40301),
            .I(N__40251));
    LocalMux I__8323 (
            .O(N__40296),
            .I(sAddressZ0Z_0));
    LocalMux I__8322 (
            .O(N__40291),
            .I(sAddressZ0Z_0));
    Odrv4 I__8321 (
            .O(N__40288),
            .I(sAddressZ0Z_0));
    LocalMux I__8320 (
            .O(N__40283),
            .I(sAddressZ0Z_0));
    LocalMux I__8319 (
            .O(N__40278),
            .I(sAddressZ0Z_0));
    LocalMux I__8318 (
            .O(N__40269),
            .I(sAddressZ0Z_0));
    Odrv4 I__8317 (
            .O(N__40264),
            .I(sAddressZ0Z_0));
    Odrv4 I__8316 (
            .O(N__40261),
            .I(sAddressZ0Z_0));
    LocalMux I__8315 (
            .O(N__40254),
            .I(sAddressZ0Z_0));
    Odrv12 I__8314 (
            .O(N__40251),
            .I(sAddressZ0Z_0));
    InMux I__8313 (
            .O(N__40230),
            .I(N__40227));
    LocalMux I__8312 (
            .O(N__40227),
            .I(N__40224));
    Odrv12 I__8311 (
            .O(N__40224),
            .I(sDAC_mem_35Z0Z_0));
    InMux I__8310 (
            .O(N__40221),
            .I(N__40218));
    LocalMux I__8309 (
            .O(N__40218),
            .I(N__40215));
    Span4Mux_v I__8308 (
            .O(N__40215),
            .I(N__40212));
    Odrv4 I__8307 (
            .O(N__40212),
            .I(sDAC_mem_35Z0Z_2));
    InMux I__8306 (
            .O(N__40209),
            .I(N__40206));
    LocalMux I__8305 (
            .O(N__40206),
            .I(N__40203));
    Span4Mux_v I__8304 (
            .O(N__40203),
            .I(N__40200));
    Span4Mux_h I__8303 (
            .O(N__40200),
            .I(N__40197));
    Odrv4 I__8302 (
            .O(N__40197),
            .I(sDAC_mem_35Z0Z_4));
    InMux I__8301 (
            .O(N__40194),
            .I(N__40191));
    LocalMux I__8300 (
            .O(N__40191),
            .I(N__40188));
    Span4Mux_v I__8299 (
            .O(N__40188),
            .I(N__40185));
    Odrv4 I__8298 (
            .O(N__40185),
            .I(sDAC_mem_35Z0Z_5));
    InMux I__8297 (
            .O(N__40182),
            .I(N__40179));
    LocalMux I__8296 (
            .O(N__40179),
            .I(N__40176));
    Odrv4 I__8295 (
            .O(N__40176),
            .I(sDAC_mem_39Z0Z_2));
    InMux I__8294 (
            .O(N__40173),
            .I(N__40170));
    LocalMux I__8293 (
            .O(N__40170),
            .I(N__40167));
    Span4Mux_v I__8292 (
            .O(N__40167),
            .I(N__40164));
    Odrv4 I__8291 (
            .O(N__40164),
            .I(sDAC_mem_39Z0Z_4));
    InMux I__8290 (
            .O(N__40161),
            .I(N__40158));
    LocalMux I__8289 (
            .O(N__40158),
            .I(N__40155));
    Span4Mux_v I__8288 (
            .O(N__40155),
            .I(N__40152));
    Odrv4 I__8287 (
            .O(N__40152),
            .I(sDAC_mem_39Z0Z_7));
    CEMux I__8286 (
            .O(N__40149),
            .I(N__40146));
    LocalMux I__8285 (
            .O(N__40146),
            .I(N__40143));
    Odrv4 I__8284 (
            .O(N__40143),
            .I(sDAC_mem_37_1_sqmuxa));
    CEMux I__8283 (
            .O(N__40140),
            .I(N__40137));
    LocalMux I__8282 (
            .O(N__40137),
            .I(sDAC_mem_39_1_sqmuxa));
    InMux I__8281 (
            .O(N__40134),
            .I(N__40131));
    LocalMux I__8280 (
            .O(N__40131),
            .I(sDAC_mem_25Z0Z_2));
    InMux I__8279 (
            .O(N__40128),
            .I(N__40125));
    LocalMux I__8278 (
            .O(N__40125),
            .I(N__40122));
    Span4Mux_v I__8277 (
            .O(N__40122),
            .I(N__40119));
    Span4Mux_v I__8276 (
            .O(N__40119),
            .I(N__40116));
    Odrv4 I__8275 (
            .O(N__40116),
            .I(sDAC_mem_25Z0Z_5));
    InMux I__8274 (
            .O(N__40113),
            .I(N__40110));
    LocalMux I__8273 (
            .O(N__40110),
            .I(sDAC_mem_25Z0Z_0));
    InMux I__8272 (
            .O(N__40107),
            .I(N__40104));
    LocalMux I__8271 (
            .O(N__40104),
            .I(N__40101));
    Odrv4 I__8270 (
            .O(N__40101),
            .I(sDAC_mem_25Z0Z_6));
    InMux I__8269 (
            .O(N__40098),
            .I(N__40095));
    LocalMux I__8268 (
            .O(N__40095),
            .I(N__40092));
    Odrv4 I__8267 (
            .O(N__40092),
            .I(sDAC_mem_25Z0Z_3));
    CEMux I__8266 (
            .O(N__40089),
            .I(N__40085));
    CEMux I__8265 (
            .O(N__40088),
            .I(N__40082));
    LocalMux I__8264 (
            .O(N__40085),
            .I(N__40079));
    LocalMux I__8263 (
            .O(N__40082),
            .I(N__40076));
    Span4Mux_v I__8262 (
            .O(N__40079),
            .I(N__40073));
    Odrv12 I__8261 (
            .O(N__40076),
            .I(sDAC_mem_34_1_sqmuxa));
    Odrv4 I__8260 (
            .O(N__40073),
            .I(sDAC_mem_34_1_sqmuxa));
    InMux I__8259 (
            .O(N__40068),
            .I(N__40065));
    LocalMux I__8258 (
            .O(N__40065),
            .I(N__40062));
    Odrv12 I__8257 (
            .O(N__40062),
            .I(sDAC_mem_39Z0Z_0));
    InMux I__8256 (
            .O(N__40059),
            .I(N__40056));
    LocalMux I__8255 (
            .O(N__40056),
            .I(N__40053));
    Span4Mux_h I__8254 (
            .O(N__40053),
            .I(N__40050));
    Odrv4 I__8253 (
            .O(N__40050),
            .I(sDAC_mem_39Z0Z_1));
    CascadeMux I__8252 (
            .O(N__40047),
            .I(sDAC_data_2_39_ns_1_10_cascade_));
    CascadeMux I__8251 (
            .O(N__40044),
            .I(N__40041));
    InMux I__8250 (
            .O(N__40041),
            .I(N__40038));
    LocalMux I__8249 (
            .O(N__40038),
            .I(N__40035));
    Odrv12 I__8248 (
            .O(N__40035),
            .I(sDAC_data_RNO_11Z0Z_10));
    InMux I__8247 (
            .O(N__40032),
            .I(N__40029));
    LocalMux I__8246 (
            .O(N__40029),
            .I(N__40026));
    Odrv4 I__8245 (
            .O(N__40026),
            .I(sDAC_mem_26Z0Z_7));
    InMux I__8244 (
            .O(N__40023),
            .I(N__40020));
    LocalMux I__8243 (
            .O(N__40020),
            .I(sDAC_data_RNO_32Z0Z_10));
    InMux I__8242 (
            .O(N__40017),
            .I(N__40014));
    LocalMux I__8241 (
            .O(N__40014),
            .I(sDAC_mem_29Z0Z_7));
    InMux I__8240 (
            .O(N__40011),
            .I(N__40008));
    LocalMux I__8239 (
            .O(N__40008),
            .I(sDAC_data_RNO_23Z0Z_10));
    InMux I__8238 (
            .O(N__40005),
            .I(N__40002));
    LocalMux I__8237 (
            .O(N__40002),
            .I(N__39999));
    Span4Mux_v I__8236 (
            .O(N__39999),
            .I(N__39996));
    Odrv4 I__8235 (
            .O(N__39996),
            .I(sDAC_mem_31Z0Z_7));
    InMux I__8234 (
            .O(N__39993),
            .I(N__39990));
    LocalMux I__8233 (
            .O(N__39990),
            .I(N__39987));
    Odrv4 I__8232 (
            .O(N__39987),
            .I(sDAC_mem_30Z0Z_7));
    InMux I__8231 (
            .O(N__39984),
            .I(N__39981));
    LocalMux I__8230 (
            .O(N__39981),
            .I(sDAC_data_RNO_24Z0Z_10));
    InMux I__8229 (
            .O(N__39978),
            .I(N__39975));
    LocalMux I__8228 (
            .O(N__39975),
            .I(sDAC_mem_24Z0Z_7));
    CEMux I__8227 (
            .O(N__39972),
            .I(N__39968));
    CEMux I__8226 (
            .O(N__39971),
            .I(N__39964));
    LocalMux I__8225 (
            .O(N__39968),
            .I(N__39961));
    CEMux I__8224 (
            .O(N__39967),
            .I(N__39958));
    LocalMux I__8223 (
            .O(N__39964),
            .I(N__39955));
    Span4Mux_h I__8222 (
            .O(N__39961),
            .I(N__39951));
    LocalMux I__8221 (
            .O(N__39958),
            .I(N__39948));
    Span4Mux_h I__8220 (
            .O(N__39955),
            .I(N__39945));
    CEMux I__8219 (
            .O(N__39954),
            .I(N__39942));
    Span4Mux_h I__8218 (
            .O(N__39951),
            .I(N__39939));
    Span4Mux_h I__8217 (
            .O(N__39948),
            .I(N__39932));
    Span4Mux_h I__8216 (
            .O(N__39945),
            .I(N__39932));
    LocalMux I__8215 (
            .O(N__39942),
            .I(N__39932));
    Span4Mux_v I__8214 (
            .O(N__39939),
            .I(N__39929));
    Span4Mux_v I__8213 (
            .O(N__39932),
            .I(N__39926));
    Odrv4 I__8212 (
            .O(N__39929),
            .I(sDAC_mem_24_1_sqmuxa));
    Odrv4 I__8211 (
            .O(N__39926),
            .I(sDAC_mem_24_1_sqmuxa));
    CascadeMux I__8210 (
            .O(N__39921),
            .I(N__39918));
    InMux I__8209 (
            .O(N__39918),
            .I(N__39915));
    LocalMux I__8208 (
            .O(N__39915),
            .I(N__39912));
    Span4Mux_h I__8207 (
            .O(N__39912),
            .I(N__39909));
    Odrv4 I__8206 (
            .O(N__39909),
            .I(sDAC_data_RNO_32Z0Z_3));
    InMux I__8205 (
            .O(N__39906),
            .I(N__39903));
    LocalMux I__8204 (
            .O(N__39903),
            .I(N__39900));
    Odrv4 I__8203 (
            .O(N__39900),
            .I(sDAC_data_RNO_31Z0Z_3));
    InMux I__8202 (
            .O(N__39897),
            .I(N__39894));
    LocalMux I__8201 (
            .O(N__39894),
            .I(sDAC_mem_25Z0Z_4));
    InMux I__8200 (
            .O(N__39891),
            .I(N__39888));
    LocalMux I__8199 (
            .O(N__39888),
            .I(sDAC_mem_25Z0Z_7));
    InMux I__8198 (
            .O(N__39885),
            .I(N__39882));
    LocalMux I__8197 (
            .O(N__39882),
            .I(N__39879));
    Span4Mux_v I__8196 (
            .O(N__39879),
            .I(N__39876));
    Span4Mux_h I__8195 (
            .O(N__39876),
            .I(N__39873));
    Span4Mux_v I__8194 (
            .O(N__39873),
            .I(N__39870));
    Odrv4 I__8193 (
            .O(N__39870),
            .I(sDAC_mem_23Z0Z_5));
    InMux I__8192 (
            .O(N__39867),
            .I(N__39864));
    LocalMux I__8191 (
            .O(N__39864),
            .I(sDAC_mem_22Z0Z_5));
    InMux I__8190 (
            .O(N__39861),
            .I(N__39858));
    LocalMux I__8189 (
            .O(N__39858),
            .I(N__39855));
    Span4Mux_v I__8188 (
            .O(N__39855),
            .I(N__39852));
    Span4Mux_h I__8187 (
            .O(N__39852),
            .I(N__39849));
    Span4Mux_v I__8186 (
            .O(N__39849),
            .I(N__39846));
    Odrv4 I__8185 (
            .O(N__39846),
            .I(sDAC_mem_23Z0Z_6));
    InMux I__8184 (
            .O(N__39843),
            .I(N__39840));
    LocalMux I__8183 (
            .O(N__39840),
            .I(N__39837));
    Span4Mux_v I__8182 (
            .O(N__39837),
            .I(N__39834));
    Odrv4 I__8181 (
            .O(N__39834),
            .I(sDAC_data_RNO_21Z0Z_9));
    InMux I__8180 (
            .O(N__39831),
            .I(N__39828));
    LocalMux I__8179 (
            .O(N__39828),
            .I(sDAC_mem_22Z0Z_6));
    CEMux I__8178 (
            .O(N__39825),
            .I(N__39821));
    CEMux I__8177 (
            .O(N__39824),
            .I(N__39818));
    LocalMux I__8176 (
            .O(N__39821),
            .I(N__39814));
    LocalMux I__8175 (
            .O(N__39818),
            .I(N__39811));
    CEMux I__8174 (
            .O(N__39817),
            .I(N__39808));
    Span4Mux_v I__8173 (
            .O(N__39814),
            .I(N__39805));
    Span4Mux_v I__8172 (
            .O(N__39811),
            .I(N__39802));
    LocalMux I__8171 (
            .O(N__39808),
            .I(N__39799));
    Span4Mux_h I__8170 (
            .O(N__39805),
            .I(N__39794));
    Span4Mux_h I__8169 (
            .O(N__39802),
            .I(N__39794));
    Span4Mux_h I__8168 (
            .O(N__39799),
            .I(N__39791));
    Odrv4 I__8167 (
            .O(N__39794),
            .I(sDAC_mem_22_1_sqmuxa));
    Odrv4 I__8166 (
            .O(N__39791),
            .I(sDAC_mem_22_1_sqmuxa));
    InMux I__8165 (
            .O(N__39786),
            .I(N__39783));
    LocalMux I__8164 (
            .O(N__39783),
            .I(sDAC_mem_29Z0Z_1));
    InMux I__8163 (
            .O(N__39780),
            .I(N__39777));
    LocalMux I__8162 (
            .O(N__39777),
            .I(sDAC_mem_30Z0Z_1));
    InMux I__8161 (
            .O(N__39774),
            .I(N__39771));
    LocalMux I__8160 (
            .O(N__39771),
            .I(N__39768));
    Span4Mux_h I__8159 (
            .O(N__39768),
            .I(N__39765));
    Odrv4 I__8158 (
            .O(N__39765),
            .I(sDAC_mem_31Z0Z_1));
    InMux I__8157 (
            .O(N__39762),
            .I(N__39759));
    LocalMux I__8156 (
            .O(N__39759),
            .I(N__39756));
    Span4Mux_h I__8155 (
            .O(N__39756),
            .I(N__39753));
    Odrv4 I__8154 (
            .O(N__39753),
            .I(sDAC_mem_31Z0Z_4));
    InMux I__8153 (
            .O(N__39750),
            .I(N__39747));
    LocalMux I__8152 (
            .O(N__39747),
            .I(sDAC_mem_30Z0Z_4));
    InMux I__8151 (
            .O(N__39744),
            .I(N__39741));
    LocalMux I__8150 (
            .O(N__39741),
            .I(N__39738));
    Odrv4 I__8149 (
            .O(N__39738),
            .I(sDAC_data_RNO_24Z0Z_7));
    CascadeMux I__8148 (
            .O(N__39735),
            .I(sDAC_data_RNO_31Z0Z_10_cascade_));
    CascadeMux I__8147 (
            .O(N__39732),
            .I(N_142_cascade_));
    InMux I__8146 (
            .O(N__39729),
            .I(N__39726));
    LocalMux I__8145 (
            .O(N__39726),
            .I(N__39723));
    Odrv4 I__8144 (
            .O(N__39723),
            .I(sDAC_mem_30Z0Z_2));
    InMux I__8143 (
            .O(N__39720),
            .I(N__39717));
    LocalMux I__8142 (
            .O(N__39717),
            .I(N__39714));
    Span4Mux_v I__8141 (
            .O(N__39714),
            .I(N__39711));
    Odrv4 I__8140 (
            .O(N__39711),
            .I(sDAC_mem_30Z0Z_3));
    InMux I__8139 (
            .O(N__39708),
            .I(N__39705));
    LocalMux I__8138 (
            .O(N__39705),
            .I(N__39702));
    Odrv4 I__8137 (
            .O(N__39702),
            .I(sDAC_mem_30Z0Z_5));
    InMux I__8136 (
            .O(N__39699),
            .I(N__39696));
    LocalMux I__8135 (
            .O(N__39696),
            .I(sDAC_mem_30Z0Z_6));
    CEMux I__8134 (
            .O(N__39693),
            .I(N__39690));
    LocalMux I__8133 (
            .O(N__39690),
            .I(sDAC_mem_30_1_sqmuxa));
    InMux I__8132 (
            .O(N__39687),
            .I(N__39684));
    LocalMux I__8131 (
            .O(N__39684),
            .I(N__39681));
    Span12Mux_v I__8130 (
            .O(N__39681),
            .I(N__39678));
    Odrv12 I__8129 (
            .O(N__39678),
            .I(sDAC_mem_36Z0Z_0));
    InMux I__8128 (
            .O(N__39675),
            .I(N__39672));
    LocalMux I__8127 (
            .O(N__39672),
            .I(N__39669));
    Span4Mux_v I__8126 (
            .O(N__39669),
            .I(N__39666));
    Span4Mux_v I__8125 (
            .O(N__39666),
            .I(N__39663));
    Odrv4 I__8124 (
            .O(N__39663),
            .I(sDAC_mem_37Z0Z_0));
    CascadeMux I__8123 (
            .O(N__39660),
            .I(sDAC_data_2_13_am_1_3_cascade_));
    InMux I__8122 (
            .O(N__39657),
            .I(N__39654));
    LocalMux I__8121 (
            .O(N__39654),
            .I(N__39651));
    Span12Mux_h I__8120 (
            .O(N__39651),
            .I(N__39648));
    Odrv12 I__8119 (
            .O(N__39648),
            .I(sDAC_mem_5Z0Z_0));
    InMux I__8118 (
            .O(N__39645),
            .I(N__39642));
    LocalMux I__8117 (
            .O(N__39642),
            .I(sDAC_mem_4Z0Z_0));
    CEMux I__8116 (
            .O(N__39639),
            .I(N__39636));
    LocalMux I__8115 (
            .O(N__39636),
            .I(N__39632));
    CEMux I__8114 (
            .O(N__39635),
            .I(N__39628));
    Span4Mux_v I__8113 (
            .O(N__39632),
            .I(N__39624));
    CEMux I__8112 (
            .O(N__39631),
            .I(N__39621));
    LocalMux I__8111 (
            .O(N__39628),
            .I(N__39618));
    CEMux I__8110 (
            .O(N__39627),
            .I(N__39615));
    Span4Mux_h I__8109 (
            .O(N__39624),
            .I(N__39610));
    LocalMux I__8108 (
            .O(N__39621),
            .I(N__39610));
    Span4Mux_h I__8107 (
            .O(N__39618),
            .I(N__39607));
    LocalMux I__8106 (
            .O(N__39615),
            .I(N__39604));
    Odrv4 I__8105 (
            .O(N__39610),
            .I(sDAC_mem_4_1_sqmuxa));
    Odrv4 I__8104 (
            .O(N__39607),
            .I(sDAC_mem_4_1_sqmuxa));
    Odrv4 I__8103 (
            .O(N__39604),
            .I(sDAC_mem_4_1_sqmuxa));
    InMux I__8102 (
            .O(N__39597),
            .I(N__39594));
    LocalMux I__8101 (
            .O(N__39594),
            .I(N__39591));
    Odrv12 I__8100 (
            .O(N__39591),
            .I(sDAC_mem_36Z0Z_1));
    InMux I__8099 (
            .O(N__39588),
            .I(N__39585));
    LocalMux I__8098 (
            .O(N__39585),
            .I(N__39582));
    Span4Mux_v I__8097 (
            .O(N__39582),
            .I(N__39579));
    Span4Mux_h I__8096 (
            .O(N__39579),
            .I(N__39576));
    Span4Mux_v I__8095 (
            .O(N__39576),
            .I(N__39573));
    Odrv4 I__8094 (
            .O(N__39573),
            .I(sDAC_mem_4Z0Z_1));
    InMux I__8093 (
            .O(N__39570),
            .I(N__39567));
    LocalMux I__8092 (
            .O(N__39567),
            .I(N__39564));
    Span4Mux_v I__8091 (
            .O(N__39564),
            .I(N__39561));
    Span4Mux_v I__8090 (
            .O(N__39561),
            .I(N__39558));
    Odrv4 I__8089 (
            .O(N__39558),
            .I(sDAC_mem_37Z0Z_1));
    CascadeMux I__8088 (
            .O(N__39555),
            .I(sDAC_data_2_13_am_1_4_cascade_));
    InMux I__8087 (
            .O(N__39552),
            .I(N__39549));
    LocalMux I__8086 (
            .O(N__39549),
            .I(N__39546));
    Span4Mux_v I__8085 (
            .O(N__39546),
            .I(N__39543));
    Span4Mux_v I__8084 (
            .O(N__39543),
            .I(N__39540));
    Odrv4 I__8083 (
            .O(N__39540),
            .I(sDAC_mem_5Z0Z_1));
    InMux I__8082 (
            .O(N__39537),
            .I(N__39534));
    LocalMux I__8081 (
            .O(N__39534),
            .I(N__39531));
    Odrv4 I__8080 (
            .O(N__39531),
            .I(sDAC_data_RNO_20Z0Z_10));
    CEMux I__8079 (
            .O(N__39528),
            .I(N__39525));
    LocalMux I__8078 (
            .O(N__39525),
            .I(N__39522));
    Span4Mux_h I__8077 (
            .O(N__39522),
            .I(N__39519));
    Span4Mux_h I__8076 (
            .O(N__39519),
            .I(N__39516));
    Odrv4 I__8075 (
            .O(N__39516),
            .I(sDAC_mem_26_1_sqmuxa));
    InMux I__8074 (
            .O(N__39513),
            .I(N__39510));
    LocalMux I__8073 (
            .O(N__39510),
            .I(N__39507));
    Odrv4 I__8072 (
            .O(N__39507),
            .I(sDAC_data_RNO_14Z0Z_10));
    InMux I__8071 (
            .O(N__39504),
            .I(N__39501));
    LocalMux I__8070 (
            .O(N__39501),
            .I(N__39498));
    Odrv4 I__8069 (
            .O(N__39498),
            .I(sDAC_data_RNO_5Z0Z_10));
    CascadeMux I__8068 (
            .O(N__39495),
            .I(sDAC_data_2_14_ns_1_10_cascade_));
    InMux I__8067 (
            .O(N__39492),
            .I(N__39489));
    LocalMux I__8066 (
            .O(N__39489),
            .I(sDAC_data_RNO_10Z0Z_10));
    InMux I__8065 (
            .O(N__39486),
            .I(N__39483));
    LocalMux I__8064 (
            .O(N__39483),
            .I(sDAC_data_RNO_2Z0Z_10));
    CascadeMux I__8063 (
            .O(N__39480),
            .I(sDAC_data_2_41_ns_1_10_cascade_));
    InMux I__8062 (
            .O(N__39477),
            .I(N__39474));
    LocalMux I__8061 (
            .O(N__39474),
            .I(sDAC_data_RNO_1Z0Z_10));
    CascadeMux I__8060 (
            .O(N__39471),
            .I(sDAC_data_2_10_cascade_));
    InMux I__8059 (
            .O(N__39468),
            .I(N__39465));
    LocalMux I__8058 (
            .O(N__39465),
            .I(N__39462));
    Span4Mux_v I__8057 (
            .O(N__39462),
            .I(N__39459));
    Span4Mux_h I__8056 (
            .O(N__39459),
            .I(N__39456));
    Sp12to4 I__8055 (
            .O(N__39456),
            .I(N__39453));
    Odrv12 I__8054 (
            .O(N__39453),
            .I(sDAC_dataZ0Z_10));
    InMux I__8053 (
            .O(N__39450),
            .I(N__39447));
    LocalMux I__8052 (
            .O(N__39447),
            .I(N__39444));
    Span12Mux_v I__8051 (
            .O(N__39444),
            .I(N__39441));
    Odrv12 I__8050 (
            .O(N__39441),
            .I(sDAC_mem_36Z0Z_7));
    InMux I__8049 (
            .O(N__39438),
            .I(N__39435));
    LocalMux I__8048 (
            .O(N__39435),
            .I(N__39432));
    Sp12to4 I__8047 (
            .O(N__39432),
            .I(N__39429));
    Odrv12 I__8046 (
            .O(N__39429),
            .I(sDAC_mem_37Z0Z_7));
    CascadeMux I__8045 (
            .O(N__39426),
            .I(sDAC_data_2_13_am_1_10_cascade_));
    InMux I__8044 (
            .O(N__39423),
            .I(N__39420));
    LocalMux I__8043 (
            .O(N__39420),
            .I(N__39417));
    Span12Mux_v I__8042 (
            .O(N__39417),
            .I(N__39414));
    Odrv12 I__8041 (
            .O(N__39414),
            .I(sDAC_mem_5Z0Z_7));
    InMux I__8040 (
            .O(N__39411),
            .I(N__39408));
    LocalMux I__8039 (
            .O(N__39408),
            .I(sDAC_data_RNO_4Z0Z_10));
    InMux I__8038 (
            .O(N__39405),
            .I(N__39402));
    LocalMux I__8037 (
            .O(N__39402),
            .I(sDAC_mem_4Z0Z_7));
    CascadeMux I__8036 (
            .O(N__39399),
            .I(N__39396));
    InMux I__8035 (
            .O(N__39396),
            .I(N__39393));
    LocalMux I__8034 (
            .O(N__39393),
            .I(N__39390));
    Span12Mux_h I__8033 (
            .O(N__39390),
            .I(N__39387));
    Odrv12 I__8032 (
            .O(N__39387),
            .I(sDAC_mem_2Z0Z_5));
    InMux I__8031 (
            .O(N__39384),
            .I(N__39381));
    LocalMux I__8030 (
            .O(N__39381),
            .I(N__39378));
    Span4Mux_v I__8029 (
            .O(N__39378),
            .I(N__39375));
    Span4Mux_v I__8028 (
            .O(N__39375),
            .I(N__39372));
    Odrv4 I__8027 (
            .O(N__39372),
            .I(sDAC_mem_34Z0Z_5));
    CascadeMux I__8026 (
            .O(N__39369),
            .I(sDAC_data_2_6_bm_1_8_cascade_));
    InMux I__8025 (
            .O(N__39366),
            .I(N__39363));
    LocalMux I__8024 (
            .O(N__39363),
            .I(sDAC_mem_3Z0Z_5));
    InMux I__8023 (
            .O(N__39360),
            .I(N__39357));
    LocalMux I__8022 (
            .O(N__39357),
            .I(N__39354));
    Span4Mux_h I__8021 (
            .O(N__39354),
            .I(N__39351));
    Span4Mux_h I__8020 (
            .O(N__39351),
            .I(N__39348));
    Odrv4 I__8019 (
            .O(N__39348),
            .I(sDAC_mem_33Z0Z_7));
    CascadeMux I__8018 (
            .O(N__39345),
            .I(sDAC_data_RNO_26Z0Z_10_cascade_));
    CascadeMux I__8017 (
            .O(N__39342),
            .I(N__39338));
    CascadeMux I__8016 (
            .O(N__39341),
            .I(N__39335));
    InMux I__8015 (
            .O(N__39338),
            .I(N__39330));
    InMux I__8014 (
            .O(N__39335),
            .I(N__39330));
    LocalMux I__8013 (
            .O(N__39330),
            .I(N__39327));
    Span4Mux_v I__8012 (
            .O(N__39327),
            .I(N__39324));
    Odrv4 I__8011 (
            .O(N__39324),
            .I(sDAC_mem_1Z0Z_7));
    InMux I__8010 (
            .O(N__39321),
            .I(N__39315));
    InMux I__8009 (
            .O(N__39320),
            .I(N__39315));
    LocalMux I__8008 (
            .O(N__39315),
            .I(N__39312));
    Span4Mux_h I__8007 (
            .O(N__39312),
            .I(N__39309));
    Odrv4 I__8006 (
            .O(N__39309),
            .I(sDAC_mem_32Z0Z_7));
    InMux I__8005 (
            .O(N__39306),
            .I(N__39303));
    LocalMux I__8004 (
            .O(N__39303),
            .I(sDAC_data_RNO_27Z0Z_10));
    CascadeMux I__8003 (
            .O(N__39300),
            .I(N__39297));
    InMux I__8002 (
            .O(N__39297),
            .I(N__39293));
    CascadeMux I__8001 (
            .O(N__39296),
            .I(N__39290));
    LocalMux I__8000 (
            .O(N__39293),
            .I(N__39287));
    InMux I__7999 (
            .O(N__39290),
            .I(N__39284));
    Span4Mux_h I__7998 (
            .O(N__39287),
            .I(N__39279));
    LocalMux I__7997 (
            .O(N__39284),
            .I(N__39279));
    Span4Mux_h I__7996 (
            .O(N__39279),
            .I(N__39276));
    Span4Mux_h I__7995 (
            .O(N__39276),
            .I(N__39273));
    Odrv4 I__7994 (
            .O(N__39273),
            .I(sDAC_mem_1Z0Z_0));
    InMux I__7993 (
            .O(N__39270),
            .I(N__39267));
    LocalMux I__7992 (
            .O(N__39267),
            .I(N__39264));
    Span4Mux_h I__7991 (
            .O(N__39264),
            .I(N__39260));
    InMux I__7990 (
            .O(N__39263),
            .I(N__39257));
    Odrv4 I__7989 (
            .O(N__39260),
            .I(sDAC_mem_32Z0Z_0));
    LocalMux I__7988 (
            .O(N__39257),
            .I(sDAC_mem_32Z0Z_0));
    InMux I__7987 (
            .O(N__39252),
            .I(N__39249));
    LocalMux I__7986 (
            .O(N__39249),
            .I(N__39246));
    Span4Mux_v I__7985 (
            .O(N__39246),
            .I(N__39243));
    Span4Mux_h I__7984 (
            .O(N__39243),
            .I(N__39240));
    Odrv4 I__7983 (
            .O(N__39240),
            .I(sDAC_mem_33Z0Z_0));
    CascadeMux I__7982 (
            .O(N__39237),
            .I(sDAC_data_RNO_26Z0Z_3_cascade_));
    InMux I__7981 (
            .O(N__39234),
            .I(N__39231));
    LocalMux I__7980 (
            .O(N__39231),
            .I(N__39228));
    Odrv4 I__7979 (
            .O(N__39228),
            .I(sDAC_data_RNO_27Z0Z_3));
    InMux I__7978 (
            .O(N__39225),
            .I(N__39222));
    LocalMux I__7977 (
            .O(N__39222),
            .I(N__39219));
    Span4Mux_v I__7976 (
            .O(N__39219),
            .I(N__39216));
    Odrv4 I__7975 (
            .O(N__39216),
            .I(sDAC_data_RNO_21Z0Z_10));
    CascadeMux I__7974 (
            .O(N__39213),
            .I(N__39210));
    InMux I__7973 (
            .O(N__39210),
            .I(N__39207));
    LocalMux I__7972 (
            .O(N__39207),
            .I(N__39204));
    Odrv12 I__7971 (
            .O(N__39204),
            .I(sDAC_data_RNO_30Z0Z_10));
    InMux I__7970 (
            .O(N__39201),
            .I(N__39198));
    LocalMux I__7969 (
            .O(N__39198),
            .I(sDAC_data_2_32_ns_1_10));
    InMux I__7968 (
            .O(N__39195),
            .I(N__39192));
    LocalMux I__7967 (
            .O(N__39192),
            .I(sDAC_data_RNO_4Z0Z_9));
    InMux I__7966 (
            .O(N__39189),
            .I(N__39186));
    LocalMux I__7965 (
            .O(N__39186),
            .I(N__39183));
    Span4Mux_v I__7964 (
            .O(N__39183),
            .I(N__39180));
    Odrv4 I__7963 (
            .O(N__39180),
            .I(sDAC_data_RNO_2Z0Z_9));
    CascadeMux I__7962 (
            .O(N__39177),
            .I(sDAC_data_RNO_1Z0Z_9_cascade_));
    CascadeMux I__7961 (
            .O(N__39174),
            .I(sDAC_data_2_9_cascade_));
    InMux I__7960 (
            .O(N__39171),
            .I(N__39168));
    LocalMux I__7959 (
            .O(N__39168),
            .I(N__39165));
    Span4Mux_v I__7958 (
            .O(N__39165),
            .I(N__39162));
    Span4Mux_h I__7957 (
            .O(N__39162),
            .I(N__39159));
    Odrv4 I__7956 (
            .O(N__39159),
            .I(sDAC_dataZ0Z_9));
    CascadeMux I__7955 (
            .O(N__39156),
            .I(N__39153));
    InMux I__7954 (
            .O(N__39153),
            .I(N__39150));
    LocalMux I__7953 (
            .O(N__39150),
            .I(N__39147));
    Odrv4 I__7952 (
            .O(N__39147),
            .I(sDAC_data_RNO_15Z0Z_9));
    InMux I__7951 (
            .O(N__39144),
            .I(N__39141));
    LocalMux I__7950 (
            .O(N__39141),
            .I(N__39138));
    Span4Mux_v I__7949 (
            .O(N__39138),
            .I(N__39135));
    Odrv4 I__7948 (
            .O(N__39135),
            .I(sDAC_data_RNO_14Z0Z_9));
    InMux I__7947 (
            .O(N__39132),
            .I(N__39129));
    LocalMux I__7946 (
            .O(N__39129),
            .I(sDAC_data_2_14_ns_1_9));
    InMux I__7945 (
            .O(N__39126),
            .I(N__39123));
    LocalMux I__7944 (
            .O(N__39123),
            .I(sDAC_data_RNO_29Z0Z_9));
    InMux I__7943 (
            .O(N__39120),
            .I(N__39117));
    LocalMux I__7942 (
            .O(N__39117),
            .I(N__39114));
    Span4Mux_h I__7941 (
            .O(N__39114),
            .I(N__39111));
    Odrv4 I__7940 (
            .O(N__39111),
            .I(sDAC_data_RNO_30Z0Z_9));
    CascadeMux I__7939 (
            .O(N__39108),
            .I(sDAC_data_2_32_ns_1_9_cascade_));
    InMux I__7938 (
            .O(N__39105),
            .I(N__39102));
    LocalMux I__7937 (
            .O(N__39102),
            .I(N__39099));
    Odrv4 I__7936 (
            .O(N__39099),
            .I(sDAC_data_RNO_20Z0Z_9));
    CascadeMux I__7935 (
            .O(N__39096),
            .I(sDAC_data_RNO_10Z0Z_9_cascade_));
    InMux I__7934 (
            .O(N__39093),
            .I(N__39090));
    LocalMux I__7933 (
            .O(N__39090),
            .I(sDAC_data_RNO_11Z0Z_9));
    InMux I__7932 (
            .O(N__39087),
            .I(N__39084));
    LocalMux I__7931 (
            .O(N__39084),
            .I(sDAC_data_2_41_ns_1_9));
    InMux I__7930 (
            .O(N__39081),
            .I(N__39078));
    LocalMux I__7929 (
            .O(N__39078),
            .I(sDAC_mem_3Z0Z_4));
    CascadeMux I__7928 (
            .O(N__39075),
            .I(sDAC_data_2_6_bm_1_7_cascade_));
    InMux I__7927 (
            .O(N__39072),
            .I(N__39069));
    LocalMux I__7926 (
            .O(N__39069),
            .I(sDAC_data_RNO_15Z0Z_7));
    InMux I__7925 (
            .O(N__39066),
            .I(N__39063));
    LocalMux I__7924 (
            .O(N__39063),
            .I(N__39060));
    Odrv12 I__7923 (
            .O(N__39060),
            .I(sDAC_mem_36Z0Z_5));
    InMux I__7922 (
            .O(N__39057),
            .I(N__39054));
    LocalMux I__7921 (
            .O(N__39054),
            .I(N__39051));
    Odrv12 I__7920 (
            .O(N__39051),
            .I(sDAC_mem_37Z0Z_5));
    CascadeMux I__7919 (
            .O(N__39048),
            .I(sDAC_data_2_13_am_1_8_cascade_));
    InMux I__7918 (
            .O(N__39045),
            .I(N__39042));
    LocalMux I__7917 (
            .O(N__39042),
            .I(N__39039));
    Span4Mux_v I__7916 (
            .O(N__39039),
            .I(N__39036));
    Odrv4 I__7915 (
            .O(N__39036),
            .I(sDAC_mem_5Z0Z_5));
    InMux I__7914 (
            .O(N__39033),
            .I(N__39030));
    LocalMux I__7913 (
            .O(N__39030),
            .I(sDAC_mem_4Z0Z_5));
    InMux I__7912 (
            .O(N__39027),
            .I(N__39024));
    LocalMux I__7911 (
            .O(N__39024),
            .I(N__39021));
    Odrv12 I__7910 (
            .O(N__39021),
            .I(sDAC_mem_36Z0Z_6));
    InMux I__7909 (
            .O(N__39018),
            .I(N__39015));
    LocalMux I__7908 (
            .O(N__39015),
            .I(N__39012));
    Odrv12 I__7907 (
            .O(N__39012),
            .I(sDAC_mem_37Z0Z_6));
    CascadeMux I__7906 (
            .O(N__39009),
            .I(sDAC_data_2_13_am_1_9_cascade_));
    InMux I__7905 (
            .O(N__39006),
            .I(N__39003));
    LocalMux I__7904 (
            .O(N__39003),
            .I(N__39000));
    Span4Mux_v I__7903 (
            .O(N__39000),
            .I(N__38997));
    Odrv4 I__7902 (
            .O(N__38997),
            .I(sDAC_mem_5Z0Z_6));
    InMux I__7901 (
            .O(N__38994),
            .I(N__38991));
    LocalMux I__7900 (
            .O(N__38991),
            .I(sDAC_mem_4Z0Z_6));
    InMux I__7899 (
            .O(N__38988),
            .I(N__38985));
    LocalMux I__7898 (
            .O(N__38985),
            .I(N__38982));
    Span4Mux_v I__7897 (
            .O(N__38982),
            .I(N__38979));
    Odrv4 I__7896 (
            .O(N__38979),
            .I(sDAC_mem_6Z0Z_7));
    CascadeMux I__7895 (
            .O(N__38976),
            .I(sDAC_data_2_13_bm_1_10_cascade_));
    InMux I__7894 (
            .O(N__38973),
            .I(N__38970));
    LocalMux I__7893 (
            .O(N__38970),
            .I(N__38967));
    Span4Mux_v I__7892 (
            .O(N__38967),
            .I(N__38964));
    Odrv4 I__7891 (
            .O(N__38964),
            .I(sDAC_mem_7Z0Z_7));
    InMux I__7890 (
            .O(N__38961),
            .I(N__38958));
    LocalMux I__7889 (
            .O(N__38958),
            .I(sDAC_mem_20Z0Z_6));
    InMux I__7888 (
            .O(N__38955),
            .I(N__38952));
    LocalMux I__7887 (
            .O(N__38952),
            .I(N__38949));
    Odrv12 I__7886 (
            .O(N__38949),
            .I(sDAC_mem_23Z0Z_7));
    InMux I__7885 (
            .O(N__38946),
            .I(N__38943));
    LocalMux I__7884 (
            .O(N__38943),
            .I(N__38940));
    Span4Mux_h I__7883 (
            .O(N__38940),
            .I(N__38937));
    Span4Mux_h I__7882 (
            .O(N__38937),
            .I(N__38934));
    Odrv4 I__7881 (
            .O(N__38934),
            .I(sDAC_mem_22Z0Z_7));
    InMux I__7880 (
            .O(N__38931),
            .I(N__38928));
    LocalMux I__7879 (
            .O(N__38928),
            .I(N__38925));
    Odrv12 I__7878 (
            .O(N__38925),
            .I(sDAC_mem_23Z0Z_0));
    InMux I__7877 (
            .O(N__38922),
            .I(N__38919));
    LocalMux I__7876 (
            .O(N__38919),
            .I(N__38916));
    Span4Mux_h I__7875 (
            .O(N__38916),
            .I(N__38913));
    Span4Mux_h I__7874 (
            .O(N__38913),
            .I(N__38910));
    Odrv4 I__7873 (
            .O(N__38910),
            .I(sDAC_mem_22Z0Z_0));
    CascadeMux I__7872 (
            .O(N__38907),
            .I(sDAC_data_2_13_bm_1_7_cascade_));
    InMux I__7871 (
            .O(N__38904),
            .I(N__38901));
    LocalMux I__7870 (
            .O(N__38901),
            .I(N__38898));
    Span4Mux_v I__7869 (
            .O(N__38898),
            .I(N__38895));
    Odrv4 I__7868 (
            .O(N__38895),
            .I(sDAC_mem_7Z0Z_4));
    InMux I__7867 (
            .O(N__38892),
            .I(N__38889));
    LocalMux I__7866 (
            .O(N__38889),
            .I(sDAC_data_RNO_5Z0Z_7));
    CascadeMux I__7865 (
            .O(N__38886),
            .I(N__38883));
    InMux I__7864 (
            .O(N__38883),
            .I(N__38880));
    LocalMux I__7863 (
            .O(N__38880),
            .I(N__38877));
    Span4Mux_h I__7862 (
            .O(N__38877),
            .I(N__38874));
    Span4Mux_v I__7861 (
            .O(N__38874),
            .I(N__38871));
    Odrv4 I__7860 (
            .O(N__38871),
            .I(sDAC_data_RNO_30Z0Z_7));
    InMux I__7859 (
            .O(N__38868),
            .I(N__38865));
    LocalMux I__7858 (
            .O(N__38865),
            .I(sDAC_data_RNO_29Z0Z_7));
    InMux I__7857 (
            .O(N__38862),
            .I(N__38859));
    LocalMux I__7856 (
            .O(N__38859),
            .I(sDAC_data_2_32_ns_1_7));
    CascadeMux I__7855 (
            .O(N__38856),
            .I(N__38853));
    InMux I__7854 (
            .O(N__38853),
            .I(N__38850));
    LocalMux I__7853 (
            .O(N__38850),
            .I(N__38847));
    Span4Mux_v I__7852 (
            .O(N__38847),
            .I(N__38844));
    Odrv4 I__7851 (
            .O(N__38844),
            .I(sDAC_mem_34Z0Z_4));
    InMux I__7850 (
            .O(N__38841),
            .I(N__38838));
    LocalMux I__7849 (
            .O(N__38838),
            .I(N__38835));
    Span4Mux_h I__7848 (
            .O(N__38835),
            .I(N__38832));
    Odrv4 I__7847 (
            .O(N__38832),
            .I(sDAC_mem_2Z0Z_4));
    InMux I__7846 (
            .O(N__38829),
            .I(N__38826));
    LocalMux I__7845 (
            .O(N__38826),
            .I(N__38823));
    Span4Mux_h I__7844 (
            .O(N__38823),
            .I(N__38820));
    Odrv4 I__7843 (
            .O(N__38820),
            .I(sDAC_mem_8Z0Z_4));
    InMux I__7842 (
            .O(N__38817),
            .I(N__38814));
    LocalMux I__7841 (
            .O(N__38814),
            .I(N__38811));
    Odrv4 I__7840 (
            .O(N__38811),
            .I(sDAC_mem_8Z0Z_6));
    InMux I__7839 (
            .O(N__38808),
            .I(N__38805));
    LocalMux I__7838 (
            .O(N__38805),
            .I(N__38802));
    Span4Mux_v I__7837 (
            .O(N__38802),
            .I(N__38799));
    Odrv4 I__7836 (
            .O(N__38799),
            .I(sDAC_mem_8Z0Z_7));
    CEMux I__7835 (
            .O(N__38796),
            .I(N__38793));
    LocalMux I__7834 (
            .O(N__38793),
            .I(sDAC_mem_8_1_sqmuxa));
    InMux I__7833 (
            .O(N__38790),
            .I(N__38787));
    LocalMux I__7832 (
            .O(N__38787),
            .I(N__38784));
    Odrv4 I__7831 (
            .O(N__38784),
            .I(sDAC_data_RNO_20Z0Z_7));
    InMux I__7830 (
            .O(N__38781),
            .I(N__38778));
    LocalMux I__7829 (
            .O(N__38778),
            .I(sDAC_mem_20Z0Z_4));
    InMux I__7828 (
            .O(N__38775),
            .I(N__38772));
    LocalMux I__7827 (
            .O(N__38772),
            .I(sDAC_mem_20Z0Z_5));
    InMux I__7826 (
            .O(N__38769),
            .I(N__38766));
    LocalMux I__7825 (
            .O(N__38766),
            .I(N__38763));
    Odrv4 I__7824 (
            .O(N__38763),
            .I(sDAC_mem_37Z0Z_2));
    InMux I__7823 (
            .O(N__38760),
            .I(N__38757));
    LocalMux I__7822 (
            .O(N__38757),
            .I(N__38754));
    Odrv4 I__7821 (
            .O(N__38754),
            .I(sDAC_mem_37Z0Z_3));
    InMux I__7820 (
            .O(N__38751),
            .I(N__38748));
    LocalMux I__7819 (
            .O(N__38748),
            .I(N__38745));
    Odrv4 I__7818 (
            .O(N__38745),
            .I(sDAC_mem_37Z0Z_4));
    InMux I__7817 (
            .O(N__38742),
            .I(N__38739));
    LocalMux I__7816 (
            .O(N__38739),
            .I(N__38736));
    Odrv4 I__7815 (
            .O(N__38736),
            .I(sDAC_mem_8Z0Z_2));
    InMux I__7814 (
            .O(N__38733),
            .I(N__38730));
    LocalMux I__7813 (
            .O(N__38730),
            .I(N__38727));
    Span4Mux_h I__7812 (
            .O(N__38727),
            .I(N__38724));
    Odrv4 I__7811 (
            .O(N__38724),
            .I(sDAC_mem_36Z0Z_2));
    InMux I__7810 (
            .O(N__38721),
            .I(N__38718));
    LocalMux I__7809 (
            .O(N__38718),
            .I(N__38715));
    Span4Mux_h I__7808 (
            .O(N__38715),
            .I(N__38712));
    Odrv4 I__7807 (
            .O(N__38712),
            .I(sDAC_mem_36Z0Z_3));
    InMux I__7806 (
            .O(N__38709),
            .I(N__38706));
    LocalMux I__7805 (
            .O(N__38706),
            .I(N__38703));
    Span4Mux_v I__7804 (
            .O(N__38703),
            .I(N__38700));
    Odrv4 I__7803 (
            .O(N__38700),
            .I(sDAC_mem_36Z0Z_4));
    InMux I__7802 (
            .O(N__38697),
            .I(N__38694));
    LocalMux I__7801 (
            .O(N__38694),
            .I(N__38691));
    Span4Mux_v I__7800 (
            .O(N__38691),
            .I(N__38688));
    Odrv4 I__7799 (
            .O(N__38688),
            .I(sDAC_mem_31Z0Z_2));
    InMux I__7798 (
            .O(N__38685),
            .I(N__38682));
    LocalMux I__7797 (
            .O(N__38682),
            .I(sDAC_data_RNO_24Z0Z_5));
    InMux I__7796 (
            .O(N__38679),
            .I(N__38676));
    LocalMux I__7795 (
            .O(N__38676),
            .I(sDAC_mem_24Z0Z_2));
    CascadeMux I__7794 (
            .O(N__38673),
            .I(N__38670));
    InMux I__7793 (
            .O(N__38670),
            .I(N__38667));
    LocalMux I__7792 (
            .O(N__38667),
            .I(sDAC_data_RNO_31Z0Z_6));
    InMux I__7791 (
            .O(N__38664),
            .I(N__38661));
    LocalMux I__7790 (
            .O(N__38661),
            .I(sDAC_data_2_39_ns_1_6));
    InMux I__7789 (
            .O(N__38658),
            .I(N__38655));
    LocalMux I__7788 (
            .O(N__38655),
            .I(N__38652));
    Odrv4 I__7787 (
            .O(N__38652),
            .I(sDAC_mem_29Z0Z_4));
    InMux I__7786 (
            .O(N__38649),
            .I(N__38646));
    LocalMux I__7785 (
            .O(N__38646),
            .I(N__38643));
    Odrv4 I__7784 (
            .O(N__38643),
            .I(sDAC_data_RNO_23Z0Z_7));
    InMux I__7783 (
            .O(N__38640),
            .I(N__38637));
    LocalMux I__7782 (
            .O(N__38637),
            .I(N__38634));
    Odrv12 I__7781 (
            .O(N__38634),
            .I(sDAC_mem_26Z0Z_3));
    InMux I__7780 (
            .O(N__38631),
            .I(N__38628));
    LocalMux I__7779 (
            .O(N__38628),
            .I(sDAC_data_RNO_32Z0Z_6));
    InMux I__7778 (
            .O(N__38625),
            .I(N__38622));
    LocalMux I__7777 (
            .O(N__38622),
            .I(N__38619));
    Span4Mux_h I__7776 (
            .O(N__38619),
            .I(N__38616));
    Span4Mux_v I__7775 (
            .O(N__38616),
            .I(N__38613));
    Odrv4 I__7774 (
            .O(N__38613),
            .I(sDAC_mem_24Z0Z_0));
    InMux I__7773 (
            .O(N__38610),
            .I(N__38607));
    LocalMux I__7772 (
            .O(N__38607),
            .I(N__38604));
    Span4Mux_h I__7771 (
            .O(N__38604),
            .I(N__38601));
    Sp12to4 I__7770 (
            .O(N__38601),
            .I(N__38598));
    Odrv12 I__7769 (
            .O(N__38598),
            .I(sDAC_mem_17Z0Z_3));
    InMux I__7768 (
            .O(N__38595),
            .I(N__38591));
    InMux I__7767 (
            .O(N__38594),
            .I(N__38588));
    LocalMux I__7766 (
            .O(N__38591),
            .I(N__38585));
    LocalMux I__7765 (
            .O(N__38588),
            .I(N__38582));
    Span4Mux_v I__7764 (
            .O(N__38585),
            .I(N__38579));
    Span4Mux_v I__7763 (
            .O(N__38582),
            .I(N__38576));
    Span4Mux_h I__7762 (
            .O(N__38579),
            .I(N__38573));
    Span4Mux_h I__7761 (
            .O(N__38576),
            .I(N__38570));
    Odrv4 I__7760 (
            .O(N__38573),
            .I(\spi_slave_inst.spi_miso ));
    Odrv4 I__7759 (
            .O(N__38570),
            .I(\spi_slave_inst.spi_miso ));
    InMux I__7758 (
            .O(N__38565),
            .I(N__38558));
    InMux I__7757 (
            .O(N__38564),
            .I(N__38558));
    InMux I__7756 (
            .O(N__38563),
            .I(N__38555));
    LocalMux I__7755 (
            .O(N__38558),
            .I(N__38549));
    LocalMux I__7754 (
            .O(N__38555),
            .I(N__38546));
    InMux I__7753 (
            .O(N__38554),
            .I(N__38541));
    InMux I__7752 (
            .O(N__38553),
            .I(N__38541));
    InMux I__7751 (
            .O(N__38552),
            .I(N__38538));
    Span4Mux_v I__7750 (
            .O(N__38549),
            .I(N__38535));
    Span4Mux_h I__7749 (
            .O(N__38546),
            .I(N__38528));
    LocalMux I__7748 (
            .O(N__38541),
            .I(N__38528));
    LocalMux I__7747 (
            .O(N__38538),
            .I(N__38528));
    Span4Mux_v I__7746 (
            .O(N__38535),
            .I(N__38522));
    Span4Mux_h I__7745 (
            .O(N__38528),
            .I(N__38519));
    InMux I__7744 (
            .O(N__38527),
            .I(N__38512));
    InMux I__7743 (
            .O(N__38526),
            .I(N__38512));
    InMux I__7742 (
            .O(N__38525),
            .I(N__38512));
    Sp12to4 I__7741 (
            .O(N__38522),
            .I(N__38509));
    Span4Mux_v I__7740 (
            .O(N__38519),
            .I(N__38506));
    LocalMux I__7739 (
            .O(N__38512),
            .I(N__38503));
    Span12Mux_h I__7738 (
            .O(N__38509),
            .I(N__38496));
    Sp12to4 I__7737 (
            .O(N__38506),
            .I(N__38496));
    Span12Mux_s11_v I__7736 (
            .O(N__38503),
            .I(N__38496));
    Span12Mux_h I__7735 (
            .O(N__38496),
            .I(N__38493));
    Odrv12 I__7734 (
            .O(N__38493),
            .I(spi_select_c));
    IoInMux I__7733 (
            .O(N__38490),
            .I(N__38487));
    LocalMux I__7732 (
            .O(N__38487),
            .I(N__38484));
    Span4Mux_s3_v I__7731 (
            .O(N__38484),
            .I(N__38481));
    Span4Mux_h I__7730 (
            .O(N__38481),
            .I(N__38478));
    Span4Mux_h I__7729 (
            .O(N__38478),
            .I(N__38475));
    Odrv4 I__7728 (
            .O(N__38475),
            .I(spi_miso_ft_c));
    CascadeMux I__7727 (
            .O(N__38472),
            .I(sDAC_data_2_39_ns_1_7_cascade_));
    InMux I__7726 (
            .O(N__38469),
            .I(N__38466));
    LocalMux I__7725 (
            .O(N__38466),
            .I(N__38463));
    Span12Mux_v I__7724 (
            .O(N__38463),
            .I(N__38460));
    Odrv12 I__7723 (
            .O(N__38460),
            .I(sDAC_data_RNO_11Z0Z_7));
    InMux I__7722 (
            .O(N__38457),
            .I(N__38454));
    LocalMux I__7721 (
            .O(N__38454),
            .I(sDAC_mem_28Z0Z_3));
    InMux I__7720 (
            .O(N__38451),
            .I(N__38448));
    LocalMux I__7719 (
            .O(N__38448),
            .I(N__38445));
    Odrv4 I__7718 (
            .O(N__38445),
            .I(sDAC_mem_26Z0Z_4));
    InMux I__7717 (
            .O(N__38442),
            .I(N__38439));
    LocalMux I__7716 (
            .O(N__38439),
            .I(sDAC_data_RNO_32Z0Z_7));
    InMux I__7715 (
            .O(N__38436),
            .I(N__38433));
    LocalMux I__7714 (
            .O(N__38433),
            .I(N__38430));
    Span4Mux_v I__7713 (
            .O(N__38430),
            .I(N__38427));
    Odrv4 I__7712 (
            .O(N__38427),
            .I(sDAC_mem_31Z0Z_3));
    InMux I__7711 (
            .O(N__38424),
            .I(N__38421));
    LocalMux I__7710 (
            .O(N__38421),
            .I(sDAC_data_RNO_24Z0Z_6));
    CascadeMux I__7709 (
            .O(N__38418),
            .I(sDAC_data_RNO_31Z0Z_5_cascade_));
    CascadeMux I__7708 (
            .O(N__38415),
            .I(sDAC_data_2_39_ns_1_5_cascade_));
    InMux I__7707 (
            .O(N__38412),
            .I(N__38409));
    LocalMux I__7706 (
            .O(N__38409),
            .I(N__38406));
    Span4Mux_v I__7705 (
            .O(N__38406),
            .I(N__38403));
    Span4Mux_v I__7704 (
            .O(N__38403),
            .I(N__38400));
    Odrv4 I__7703 (
            .O(N__38400),
            .I(sDAC_data_RNO_11Z0Z_5));
    InMux I__7702 (
            .O(N__38397),
            .I(N__38394));
    LocalMux I__7701 (
            .O(N__38394),
            .I(N__38391));
    Odrv12 I__7700 (
            .O(N__38391),
            .I(sDAC_mem_26Z0Z_2));
    InMux I__7699 (
            .O(N__38388),
            .I(N__38385));
    LocalMux I__7698 (
            .O(N__38385),
            .I(N__38382));
    Odrv4 I__7697 (
            .O(N__38382),
            .I(sDAC_data_RNO_32Z0Z_5));
    InMux I__7696 (
            .O(N__38379),
            .I(N__38376));
    LocalMux I__7695 (
            .O(N__38376),
            .I(N__38373));
    Odrv4 I__7694 (
            .O(N__38373),
            .I(sDAC_mem_29Z0Z_2));
    InMux I__7693 (
            .O(N__38370),
            .I(N__38367));
    LocalMux I__7692 (
            .O(N__38367),
            .I(sDAC_data_RNO_23Z0Z_5));
    InMux I__7691 (
            .O(N__38364),
            .I(N__38361));
    LocalMux I__7690 (
            .O(N__38361),
            .I(N__38358));
    Odrv12 I__7689 (
            .O(N__38358),
            .I(sDAC_mem_29Z0Z_5));
    InMux I__7688 (
            .O(N__38355),
            .I(N__38352));
    LocalMux I__7687 (
            .O(N__38352),
            .I(N__38349));
    Odrv12 I__7686 (
            .O(N__38349),
            .I(sDAC_mem_29Z0Z_6));
    CEMux I__7685 (
            .O(N__38346),
            .I(N__38343));
    LocalMux I__7684 (
            .O(N__38343),
            .I(N__38340));
    Span4Mux_h I__7683 (
            .O(N__38340),
            .I(N__38337));
    Span4Mux_v I__7682 (
            .O(N__38337),
            .I(N__38334));
    Odrv4 I__7681 (
            .O(N__38334),
            .I(sDAC_mem_29_1_sqmuxa));
    InMux I__7680 (
            .O(N__38331),
            .I(N__38328));
    LocalMux I__7679 (
            .O(N__38328),
            .I(sDAC_mem_29Z0Z_3));
    InMux I__7678 (
            .O(N__38325),
            .I(N__38322));
    LocalMux I__7677 (
            .O(N__38322),
            .I(sDAC_data_RNO_23Z0Z_6));
    InMux I__7676 (
            .O(N__38319),
            .I(N__38316));
    LocalMux I__7675 (
            .O(N__38316),
            .I(N__38313));
    Span4Mux_h I__7674 (
            .O(N__38313),
            .I(N__38310));
    Odrv4 I__7673 (
            .O(N__38310),
            .I(sDAC_mem_24Z0Z_4));
    CascadeMux I__7672 (
            .O(N__38307),
            .I(sDAC_data_RNO_31Z0Z_7_cascade_));
    CascadeMux I__7671 (
            .O(N__38304),
            .I(sDAC_data_RNO_18Z0Z_9_cascade_));
    InMux I__7670 (
            .O(N__38301),
            .I(N__38298));
    LocalMux I__7669 (
            .O(N__38298),
            .I(sDAC_data_RNO_19Z0Z_9));
    InMux I__7668 (
            .O(N__38295),
            .I(N__38292));
    LocalMux I__7667 (
            .O(N__38292),
            .I(N__38289));
    Span4Mux_v I__7666 (
            .O(N__38289),
            .I(N__38286));
    Odrv4 I__7665 (
            .O(N__38286),
            .I(sDAC_data_2_24_ns_1_9));
    InMux I__7664 (
            .O(N__38283),
            .I(N__38279));
    InMux I__7663 (
            .O(N__38282),
            .I(N__38276));
    LocalMux I__7662 (
            .O(N__38279),
            .I(N__38273));
    LocalMux I__7661 (
            .O(N__38276),
            .I(sCounterADCZ0Z_1));
    Odrv12 I__7660 (
            .O(N__38273),
            .I(sCounterADCZ0Z_1));
    InMux I__7659 (
            .O(N__38268),
            .I(N__38264));
    InMux I__7658 (
            .O(N__38267),
            .I(N__38261));
    LocalMux I__7657 (
            .O(N__38264),
            .I(N__38258));
    LocalMux I__7656 (
            .O(N__38261),
            .I(sCounterADCZ0Z_0));
    Odrv4 I__7655 (
            .O(N__38258),
            .I(sCounterADCZ0Z_0));
    InMux I__7654 (
            .O(N__38253),
            .I(N__38250));
    LocalMux I__7653 (
            .O(N__38250),
            .I(un11_sacqtime_NE_3));
    InMux I__7652 (
            .O(N__38247),
            .I(N__38244));
    LocalMux I__7651 (
            .O(N__38244),
            .I(un11_sacqtime_NE_2));
    CascadeMux I__7650 (
            .O(N__38241),
            .I(un11_sacqtime_NE_0_0_cascade_));
    InMux I__7649 (
            .O(N__38238),
            .I(N__38235));
    LocalMux I__7648 (
            .O(N__38235),
            .I(N__38232));
    Odrv4 I__7647 (
            .O(N__38232),
            .I(un11_sacqtime_NE_1));
    CascadeMux I__7646 (
            .O(N__38229),
            .I(N__38222));
    InMux I__7645 (
            .O(N__38228),
            .I(N__38213));
    InMux I__7644 (
            .O(N__38227),
            .I(N__38213));
    InMux I__7643 (
            .O(N__38226),
            .I(N__38213));
    InMux I__7642 (
            .O(N__38225),
            .I(N__38213));
    InMux I__7641 (
            .O(N__38222),
            .I(N__38210));
    LocalMux I__7640 (
            .O(N__38213),
            .I(N__38207));
    LocalMux I__7639 (
            .O(N__38210),
            .I(N__38200));
    Span4Mux_h I__7638 (
            .O(N__38207),
            .I(N__38197));
    InMux I__7637 (
            .O(N__38206),
            .I(N__38188));
    InMux I__7636 (
            .O(N__38205),
            .I(N__38188));
    InMux I__7635 (
            .O(N__38204),
            .I(N__38188));
    InMux I__7634 (
            .O(N__38203),
            .I(N__38188));
    Span4Mux_v I__7633 (
            .O(N__38200),
            .I(N__38185));
    Span4Mux_h I__7632 (
            .O(N__38197),
            .I(N__38178));
    LocalMux I__7631 (
            .O(N__38188),
            .I(N__38178));
    Span4Mux_h I__7630 (
            .O(N__38185),
            .I(N__38178));
    Odrv4 I__7629 (
            .O(N__38178),
            .I(un11_sacqtime_NE_0));
    InMux I__7628 (
            .O(N__38175),
            .I(N__38172));
    LocalMux I__7627 (
            .O(N__38172),
            .I(sDAC_mem_31Z0Z_6));
    InMux I__7626 (
            .O(N__38169),
            .I(N__38166));
    LocalMux I__7625 (
            .O(N__38166),
            .I(N__38163));
    Span4Mux_v I__7624 (
            .O(N__38163),
            .I(N__38160));
    Odrv4 I__7623 (
            .O(N__38160),
            .I(sDAC_data_RNO_24Z0Z_9));
    InMux I__7622 (
            .O(N__38157),
            .I(N__38154));
    LocalMux I__7621 (
            .O(N__38154),
            .I(sDAC_mem_24Z0Z_5));
    CascadeMux I__7620 (
            .O(N__38151),
            .I(N__38148));
    InMux I__7619 (
            .O(N__38148),
            .I(N__38145));
    LocalMux I__7618 (
            .O(N__38145),
            .I(N__38142));
    Span4Mux_h I__7617 (
            .O(N__38142),
            .I(N__38139));
    Span4Mux_v I__7616 (
            .O(N__38139),
            .I(N__38136));
    Odrv4 I__7615 (
            .O(N__38136),
            .I(sDAC_data_RNO_31Z0Z_9));
    InMux I__7614 (
            .O(N__38133),
            .I(N__38130));
    LocalMux I__7613 (
            .O(N__38130),
            .I(N__38127));
    Span4Mux_v I__7612 (
            .O(N__38127),
            .I(N__38124));
    Odrv4 I__7611 (
            .O(N__38124),
            .I(sDAC_data_RNO_32Z0Z_9));
    InMux I__7610 (
            .O(N__38121),
            .I(N__38118));
    LocalMux I__7609 (
            .O(N__38118),
            .I(N__38115));
    Odrv4 I__7608 (
            .O(N__38115),
            .I(sDAC_data_2_39_ns_1_9));
    InMux I__7607 (
            .O(N__38112),
            .I(N__38109));
    LocalMux I__7606 (
            .O(N__38109),
            .I(N__38106));
    Span4Mux_v I__7605 (
            .O(N__38106),
            .I(N__38103));
    Odrv4 I__7604 (
            .O(N__38103),
            .I(sDAC_mem_26Z0Z_0));
    InMux I__7603 (
            .O(N__38100),
            .I(N__38097));
    LocalMux I__7602 (
            .O(N__38097),
            .I(sDAC_mem_26Z0Z_5));
    InMux I__7601 (
            .O(N__38094),
            .I(N__38091));
    LocalMux I__7600 (
            .O(N__38091),
            .I(N__38088));
    Span4Mux_v I__7599 (
            .O(N__38088),
            .I(N__38085));
    Odrv4 I__7598 (
            .O(N__38085),
            .I(sDAC_mem_26Z0Z_6));
    CascadeMux I__7597 (
            .O(N__38082),
            .I(N__38065));
    CascadeMux I__7596 (
            .O(N__38081),
            .I(N__38062));
    CascadeMux I__7595 (
            .O(N__38080),
            .I(N__38059));
    CascadeMux I__7594 (
            .O(N__38079),
            .I(N__38056));
    CascadeMux I__7593 (
            .O(N__38078),
            .I(N__38053));
    CascadeMux I__7592 (
            .O(N__38077),
            .I(N__38050));
    CascadeMux I__7591 (
            .O(N__38076),
            .I(N__38047));
    CascadeMux I__7590 (
            .O(N__38075),
            .I(N__38044));
    CascadeMux I__7589 (
            .O(N__38074),
            .I(N__38040));
    CascadeMux I__7588 (
            .O(N__38073),
            .I(N__38037));
    CascadeMux I__7587 (
            .O(N__38072),
            .I(N__38034));
    CascadeMux I__7586 (
            .O(N__38071),
            .I(N__38030));
    CascadeMux I__7585 (
            .O(N__38070),
            .I(N__38027));
    CascadeMux I__7584 (
            .O(N__38069),
            .I(N__38024));
    CascadeMux I__7583 (
            .O(N__38068),
            .I(N__38021));
    InMux I__7582 (
            .O(N__38065),
            .I(N__38009));
    InMux I__7581 (
            .O(N__38062),
            .I(N__38009));
    InMux I__7580 (
            .O(N__38059),
            .I(N__38009));
    InMux I__7579 (
            .O(N__38056),
            .I(N__38009));
    InMux I__7578 (
            .O(N__38053),
            .I(N__38000));
    InMux I__7577 (
            .O(N__38050),
            .I(N__38000));
    InMux I__7576 (
            .O(N__38047),
            .I(N__38000));
    InMux I__7575 (
            .O(N__38044),
            .I(N__38000));
    InMux I__7574 (
            .O(N__38043),
            .I(N__37991));
    InMux I__7573 (
            .O(N__38040),
            .I(N__37991));
    InMux I__7572 (
            .O(N__38037),
            .I(N__37991));
    InMux I__7571 (
            .O(N__38034),
            .I(N__37991));
    InMux I__7570 (
            .O(N__38033),
            .I(N__37982));
    InMux I__7569 (
            .O(N__38030),
            .I(N__37982));
    InMux I__7568 (
            .O(N__38027),
            .I(N__37982));
    InMux I__7567 (
            .O(N__38024),
            .I(N__37982));
    InMux I__7566 (
            .O(N__38021),
            .I(N__37977));
    InMux I__7565 (
            .O(N__38020),
            .I(N__37977));
    InMux I__7564 (
            .O(N__38019),
            .I(N__37972));
    InMux I__7563 (
            .O(N__38018),
            .I(N__37972));
    LocalMux I__7562 (
            .O(N__38009),
            .I(N__37959));
    LocalMux I__7561 (
            .O(N__38000),
            .I(N__37959));
    LocalMux I__7560 (
            .O(N__37991),
            .I(N__37954));
    LocalMux I__7559 (
            .O(N__37982),
            .I(N__37954));
    LocalMux I__7558 (
            .O(N__37977),
            .I(N__37951));
    LocalMux I__7557 (
            .O(N__37972),
            .I(N__37948));
    CascadeMux I__7556 (
            .O(N__37971),
            .I(N__37945));
    CascadeMux I__7555 (
            .O(N__37970),
            .I(N__37941));
    CascadeMux I__7554 (
            .O(N__37969),
            .I(N__37937));
    CascadeMux I__7553 (
            .O(N__37968),
            .I(N__37933));
    CascadeMux I__7552 (
            .O(N__37967),
            .I(N__37925));
    CascadeMux I__7551 (
            .O(N__37966),
            .I(N__37921));
    CascadeMux I__7550 (
            .O(N__37965),
            .I(N__37917));
    CascadeMux I__7549 (
            .O(N__37964),
            .I(N__37913));
    Span4Mux_v I__7548 (
            .O(N__37959),
            .I(N__37904));
    Span4Mux_v I__7547 (
            .O(N__37954),
            .I(N__37898));
    Span4Mux_v I__7546 (
            .O(N__37951),
            .I(N__37898));
    Span4Mux_h I__7545 (
            .O(N__37948),
            .I(N__37895));
    InMux I__7544 (
            .O(N__37945),
            .I(N__37878));
    InMux I__7543 (
            .O(N__37944),
            .I(N__37878));
    InMux I__7542 (
            .O(N__37941),
            .I(N__37878));
    InMux I__7541 (
            .O(N__37940),
            .I(N__37878));
    InMux I__7540 (
            .O(N__37937),
            .I(N__37878));
    InMux I__7539 (
            .O(N__37936),
            .I(N__37878));
    InMux I__7538 (
            .O(N__37933),
            .I(N__37878));
    InMux I__7537 (
            .O(N__37932),
            .I(N__37878));
    CascadeMux I__7536 (
            .O(N__37931),
            .I(N__37875));
    CascadeMux I__7535 (
            .O(N__37930),
            .I(N__37870));
    CascadeMux I__7534 (
            .O(N__37929),
            .I(N__37866));
    CascadeMux I__7533 (
            .O(N__37928),
            .I(N__37862));
    InMux I__7532 (
            .O(N__37925),
            .I(N__37845));
    InMux I__7531 (
            .O(N__37924),
            .I(N__37845));
    InMux I__7530 (
            .O(N__37921),
            .I(N__37845));
    InMux I__7529 (
            .O(N__37920),
            .I(N__37845));
    InMux I__7528 (
            .O(N__37917),
            .I(N__37845));
    InMux I__7527 (
            .O(N__37916),
            .I(N__37845));
    InMux I__7526 (
            .O(N__37913),
            .I(N__37845));
    InMux I__7525 (
            .O(N__37912),
            .I(N__37845));
    CascadeMux I__7524 (
            .O(N__37911),
            .I(N__37842));
    CascadeMux I__7523 (
            .O(N__37910),
            .I(N__37838));
    CascadeMux I__7522 (
            .O(N__37909),
            .I(N__37834));
    CascadeMux I__7521 (
            .O(N__37908),
            .I(N__37830));
    CascadeMux I__7520 (
            .O(N__37907),
            .I(N__37825));
    Sp12to4 I__7519 (
            .O(N__37904),
            .I(N__37821));
    InMux I__7518 (
            .O(N__37903),
            .I(N__37818));
    Span4Mux_v I__7517 (
            .O(N__37898),
            .I(N__37811));
    Span4Mux_h I__7516 (
            .O(N__37895),
            .I(N__37811));
    LocalMux I__7515 (
            .O(N__37878),
            .I(N__37811));
    InMux I__7514 (
            .O(N__37875),
            .I(N__37794));
    InMux I__7513 (
            .O(N__37874),
            .I(N__37794));
    InMux I__7512 (
            .O(N__37873),
            .I(N__37794));
    InMux I__7511 (
            .O(N__37870),
            .I(N__37794));
    InMux I__7510 (
            .O(N__37869),
            .I(N__37794));
    InMux I__7509 (
            .O(N__37866),
            .I(N__37794));
    InMux I__7508 (
            .O(N__37865),
            .I(N__37794));
    InMux I__7507 (
            .O(N__37862),
            .I(N__37794));
    LocalMux I__7506 (
            .O(N__37845),
            .I(N__37791));
    InMux I__7505 (
            .O(N__37842),
            .I(N__37774));
    InMux I__7504 (
            .O(N__37841),
            .I(N__37774));
    InMux I__7503 (
            .O(N__37838),
            .I(N__37774));
    InMux I__7502 (
            .O(N__37837),
            .I(N__37774));
    InMux I__7501 (
            .O(N__37834),
            .I(N__37774));
    InMux I__7500 (
            .O(N__37833),
            .I(N__37774));
    InMux I__7499 (
            .O(N__37830),
            .I(N__37774));
    InMux I__7498 (
            .O(N__37829),
            .I(N__37774));
    InMux I__7497 (
            .O(N__37828),
            .I(N__37767));
    InMux I__7496 (
            .O(N__37825),
            .I(N__37767));
    InMux I__7495 (
            .O(N__37824),
            .I(N__37767));
    Span12Mux_h I__7494 (
            .O(N__37821),
            .I(N__37762));
    LocalMux I__7493 (
            .O(N__37818),
            .I(N__37762));
    Span4Mux_h I__7492 (
            .O(N__37811),
            .I(N__37757));
    LocalMux I__7491 (
            .O(N__37794),
            .I(N__37757));
    Span4Mux_v I__7490 (
            .O(N__37791),
            .I(N__37752));
    LocalMux I__7489 (
            .O(N__37774),
            .I(N__37752));
    LocalMux I__7488 (
            .O(N__37767),
            .I(N__37749));
    Span12Mux_v I__7487 (
            .O(N__37762),
            .I(N__37746));
    Span4Mux_v I__7486 (
            .O(N__37757),
            .I(N__37743));
    Span4Mux_h I__7485 (
            .O(N__37752),
            .I(N__37738));
    Span4Mux_v I__7484 (
            .O(N__37749),
            .I(N__37738));
    Odrv12 I__7483 (
            .O(N__37746),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__7482 (
            .O(N__37743),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__7481 (
            .O(N__37738),
            .I(CONSTANT_ONE_NET));
    InMux I__7480 (
            .O(N__37731),
            .I(N__37728));
    LocalMux I__7479 (
            .O(N__37728),
            .I(N__37725));
    Span12Mux_h I__7478 (
            .O(N__37725),
            .I(N__37722));
    Odrv12 I__7477 (
            .O(N__37722),
            .I(sDAC_dataZ0Z_13));
    InMux I__7476 (
            .O(N__37719),
            .I(N__37716));
    LocalMux I__7475 (
            .O(N__37716),
            .I(N__37713));
    Span4Mux_h I__7474 (
            .O(N__37713),
            .I(N__37710));
    Span4Mux_v I__7473 (
            .O(N__37710),
            .I(N__37707));
    Span4Mux_h I__7472 (
            .O(N__37707),
            .I(N__37704));
    Odrv4 I__7471 (
            .O(N__37704),
            .I(sDAC_dataZ0Z_14));
    InMux I__7470 (
            .O(N__37701),
            .I(N__37698));
    LocalMux I__7469 (
            .O(N__37698),
            .I(N__37695));
    Span4Mux_h I__7468 (
            .O(N__37695),
            .I(N__37692));
    Span4Mux_v I__7467 (
            .O(N__37692),
            .I(N__37689));
    Span4Mux_h I__7466 (
            .O(N__37689),
            .I(N__37686));
    Odrv4 I__7465 (
            .O(N__37686),
            .I(sDAC_dataZ0Z_15));
    CascadeMux I__7464 (
            .O(N__37683),
            .I(sDAC_data_RNO_31Z0Z_8_cascade_));
    CascadeMux I__7463 (
            .O(N__37680),
            .I(sDAC_data_2_39_ns_1_8_cascade_));
    InMux I__7462 (
            .O(N__37677),
            .I(N__37674));
    LocalMux I__7461 (
            .O(N__37674),
            .I(sDAC_data_RNO_32Z0Z_8));
    InMux I__7460 (
            .O(N__37671),
            .I(N__37668));
    LocalMux I__7459 (
            .O(N__37668),
            .I(sDAC_data_RNO_23Z0Z_8));
    InMux I__7458 (
            .O(N__37665),
            .I(N__37662));
    LocalMux I__7457 (
            .O(N__37662),
            .I(sDAC_mem_31Z0Z_5));
    InMux I__7456 (
            .O(N__37659),
            .I(N__37656));
    LocalMux I__7455 (
            .O(N__37656),
            .I(sDAC_data_RNO_24Z0Z_8));
    InMux I__7454 (
            .O(N__37653),
            .I(N__37650));
    LocalMux I__7453 (
            .O(N__37650),
            .I(sDAC_data_RNO_17Z0Z_10));
    InMux I__7452 (
            .O(N__37647),
            .I(N__37644));
    LocalMux I__7451 (
            .O(N__37644),
            .I(sDAC_data_2_24_ns_1_10));
    CascadeMux I__7450 (
            .O(N__37641),
            .I(sDAC_data_RNO_8Z0Z_10_cascade_));
    CascadeMux I__7449 (
            .O(N__37638),
            .I(sDAC_data_2_20_am_1_10_cascade_));
    InMux I__7448 (
            .O(N__37635),
            .I(N__37632));
    LocalMux I__7447 (
            .O(N__37632),
            .I(sDAC_data_RNO_7Z0Z_10));
    InMux I__7446 (
            .O(N__37629),
            .I(N__37626));
    LocalMux I__7445 (
            .O(N__37626),
            .I(sDAC_mem_28Z0Z_6));
    InMux I__7444 (
            .O(N__37623),
            .I(N__37620));
    LocalMux I__7443 (
            .O(N__37620),
            .I(N__37617));
    Span4Mux_h I__7442 (
            .O(N__37617),
            .I(N__37614));
    Span4Mux_h I__7441 (
            .O(N__37614),
            .I(N__37611));
    Span4Mux_v I__7440 (
            .O(N__37611),
            .I(N__37608));
    Odrv4 I__7439 (
            .O(N__37608),
            .I(sDAC_dataZ0Z_1));
    InMux I__7438 (
            .O(N__37605),
            .I(N__37602));
    LocalMux I__7437 (
            .O(N__37602),
            .I(N__37599));
    Span4Mux_v I__7436 (
            .O(N__37599),
            .I(N__37596));
    Span4Mux_v I__7435 (
            .O(N__37596),
            .I(N__37593));
    Span4Mux_h I__7434 (
            .O(N__37593),
            .I(N__37590));
    Odrv4 I__7433 (
            .O(N__37590),
            .I(sDAC_dataZ0Z_11));
    InMux I__7432 (
            .O(N__37587),
            .I(N__37584));
    LocalMux I__7431 (
            .O(N__37584),
            .I(N__37581));
    Span4Mux_v I__7430 (
            .O(N__37581),
            .I(N__37578));
    Span4Mux_v I__7429 (
            .O(N__37578),
            .I(N__37575));
    Span4Mux_h I__7428 (
            .O(N__37575),
            .I(N__37572));
    Odrv4 I__7427 (
            .O(N__37572),
            .I(sDAC_dataZ0Z_12));
    InMux I__7426 (
            .O(N__37569),
            .I(N__37566));
    LocalMux I__7425 (
            .O(N__37566),
            .I(N__37563));
    Odrv4 I__7424 (
            .O(N__37563),
            .I(sDAC_mem_17Z0Z_6));
    InMux I__7423 (
            .O(N__37560),
            .I(N__37557));
    LocalMux I__7422 (
            .O(N__37557),
            .I(sDAC_mem_16Z0Z_6));
    InMux I__7421 (
            .O(N__37554),
            .I(sDAC_mem_pointer_0_cry_1));
    InMux I__7420 (
            .O(N__37551),
            .I(sDAC_mem_pointer_0_cry_2));
    InMux I__7419 (
            .O(N__37548),
            .I(sDAC_mem_pointer_0_cry_3));
    InMux I__7418 (
            .O(N__37545),
            .I(sDAC_mem_pointer_0_cry_4));
    CascadeMux I__7417 (
            .O(N__37542),
            .I(sDAC_data_RNO_23Z0Z_9_cascade_));
    CascadeMux I__7416 (
            .O(N__37539),
            .I(sDAC_data_RNO_17Z0Z_9_cascade_));
    CascadeMux I__7415 (
            .O(N__37536),
            .I(sDAC_data_RNO_8Z0Z_9_cascade_));
    CascadeMux I__7414 (
            .O(N__37533),
            .I(sDAC_data_2_20_am_1_9_cascade_));
    InMux I__7413 (
            .O(N__37530),
            .I(N__37527));
    LocalMux I__7412 (
            .O(N__37527),
            .I(sDAC_data_RNO_7Z0Z_9));
    InMux I__7411 (
            .O(N__37524),
            .I(N__37521));
    LocalMux I__7410 (
            .O(N__37521),
            .I(N__37518));
    Odrv4 I__7409 (
            .O(N__37518),
            .I(sDAC_mem_17Z0Z_4));
    InMux I__7408 (
            .O(N__37515),
            .I(N__37512));
    LocalMux I__7407 (
            .O(N__37512),
            .I(sDAC_mem_16Z0Z_4));
    InMux I__7406 (
            .O(N__37509),
            .I(N__37506));
    LocalMux I__7405 (
            .O(N__37506),
            .I(N__37503));
    Odrv12 I__7404 (
            .O(N__37503),
            .I(sDAC_mem_17Z0Z_5));
    InMux I__7403 (
            .O(N__37500),
            .I(N__37497));
    LocalMux I__7402 (
            .O(N__37497),
            .I(sDAC_mem_16Z0Z_5));
    InMux I__7401 (
            .O(N__37494),
            .I(N__37476));
    InMux I__7400 (
            .O(N__37493),
            .I(N__37476));
    InMux I__7399 (
            .O(N__37492),
            .I(N__37476));
    InMux I__7398 (
            .O(N__37491),
            .I(N__37476));
    InMux I__7397 (
            .O(N__37490),
            .I(N__37476));
    InMux I__7396 (
            .O(N__37489),
            .I(N__37476));
    LocalMux I__7395 (
            .O(N__37476),
            .I(N_279));
    CascadeMux I__7394 (
            .O(N__37473),
            .I(N_279_cascade_));
    InMux I__7393 (
            .O(N__37470),
            .I(N__37467));
    LocalMux I__7392 (
            .O(N__37467),
            .I(N__37464));
    Odrv4 I__7391 (
            .O(N__37464),
            .I(sDAC_data_RNO_21Z0Z_7));
    CascadeMux I__7390 (
            .O(N__37461),
            .I(sDAC_data_2_14_ns_1_7_cascade_));
    InMux I__7389 (
            .O(N__37458),
            .I(N__37455));
    LocalMux I__7388 (
            .O(N__37455),
            .I(N__37452));
    Odrv4 I__7387 (
            .O(N__37452),
            .I(sDAC_data_RNO_4Z0Z_7));
    InMux I__7386 (
            .O(N__37449),
            .I(N__37446));
    LocalMux I__7385 (
            .O(N__37446),
            .I(sDAC_data_RNO_10Z0Z_7));
    InMux I__7384 (
            .O(N__37443),
            .I(N__37440));
    LocalMux I__7383 (
            .O(N__37440),
            .I(sDAC_data_RNO_2Z0Z_7));
    CascadeMux I__7382 (
            .O(N__37437),
            .I(sDAC_data_2_41_ns_1_7_cascade_));
    InMux I__7381 (
            .O(N__37434),
            .I(N__37431));
    LocalMux I__7380 (
            .O(N__37431),
            .I(sDAC_data_RNO_1Z0Z_7));
    CascadeMux I__7379 (
            .O(N__37428),
            .I(sDAC_data_2_7_cascade_));
    InMux I__7378 (
            .O(N__37425),
            .I(N__37422));
    LocalMux I__7377 (
            .O(N__37422),
            .I(N__37419));
    Span4Mux_h I__7376 (
            .O(N__37419),
            .I(N__37416));
    Odrv4 I__7375 (
            .O(N__37416),
            .I(sDAC_dataZ0Z_7));
    InMux I__7374 (
            .O(N__37413),
            .I(N__37410));
    LocalMux I__7373 (
            .O(N__37410),
            .I(sDAC_mem_5Z0Z_4));
    CEMux I__7372 (
            .O(N__37407),
            .I(N__37404));
    LocalMux I__7371 (
            .O(N__37404),
            .I(N__37401));
    Span4Mux_h I__7370 (
            .O(N__37401),
            .I(N__37398));
    Odrv4 I__7369 (
            .O(N__37398),
            .I(sDAC_mem_2_1_sqmuxa));
    CEMux I__7368 (
            .O(N__37395),
            .I(N__37392));
    LocalMux I__7367 (
            .O(N__37392),
            .I(N__37389));
    Span4Mux_v I__7366 (
            .O(N__37389),
            .I(N__37386));
    Odrv4 I__7365 (
            .O(N__37386),
            .I(sDAC_mem_5_1_sqmuxa));
    CEMux I__7364 (
            .O(N__37383),
            .I(N__37380));
    LocalMux I__7363 (
            .O(N__37380),
            .I(N__37377));
    Span4Mux_v I__7362 (
            .O(N__37377),
            .I(N__37374));
    Span4Mux_h I__7361 (
            .O(N__37374),
            .I(N__37371));
    Odrv4 I__7360 (
            .O(N__37371),
            .I(sDAC_mem_7_1_sqmuxa));
    InMux I__7359 (
            .O(N__37368),
            .I(N__37365));
    LocalMux I__7358 (
            .O(N__37365),
            .I(N__37362));
    Odrv4 I__7357 (
            .O(N__37362),
            .I(sDAC_mem_7Z0Z_2));
    InMux I__7356 (
            .O(N__37359),
            .I(N__37356));
    LocalMux I__7355 (
            .O(N__37356),
            .I(sDAC_mem_5Z0Z_2));
    InMux I__7354 (
            .O(N__37353),
            .I(N__37350));
    LocalMux I__7353 (
            .O(N__37350),
            .I(sDAC_mem_5Z0Z_3));
    InMux I__7352 (
            .O(N__37347),
            .I(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4 ));
    InMux I__7351 (
            .O(N__37344),
            .I(N__37340));
    InMux I__7350 (
            .O(N__37343),
            .I(N__37337));
    LocalMux I__7349 (
            .O(N__37340),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5 ));
    LocalMux I__7348 (
            .O(N__37337),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5 ));
    InMux I__7347 (
            .O(N__37332),
            .I(N__37329));
    LocalMux I__7346 (
            .O(N__37329),
            .I(N__37326));
    Span4Mux_v I__7345 (
            .O(N__37326),
            .I(N__37323));
    Odrv4 I__7344 (
            .O(N__37323),
            .I(sDAC_mem_34Z0Z_0));
    InMux I__7343 (
            .O(N__37320),
            .I(N__37317));
    LocalMux I__7342 (
            .O(N__37317),
            .I(N__37314));
    Span4Mux_v I__7341 (
            .O(N__37314),
            .I(N__37311));
    Odrv4 I__7340 (
            .O(N__37311),
            .I(sDAC_mem_34Z0Z_2));
    InMux I__7339 (
            .O(N__37308),
            .I(N__37305));
    LocalMux I__7338 (
            .O(N__37305),
            .I(N__37302));
    Span4Mux_v I__7337 (
            .O(N__37302),
            .I(N__37299));
    Odrv4 I__7336 (
            .O(N__37299),
            .I(sDAC_mem_34Z0Z_6));
    InMux I__7335 (
            .O(N__37296),
            .I(N__37293));
    LocalMux I__7334 (
            .O(N__37293),
            .I(sDAC_mem_7Z0Z_0));
    InMux I__7333 (
            .O(N__37290),
            .I(N__37287));
    LocalMux I__7332 (
            .O(N__37287),
            .I(sDAC_mem_7Z0Z_1));
    InMux I__7331 (
            .O(N__37284),
            .I(N__37281));
    LocalMux I__7330 (
            .O(N__37281),
            .I(sDAC_mem_16Z0Z_2));
    InMux I__7329 (
            .O(N__37278),
            .I(N__37275));
    LocalMux I__7328 (
            .O(N__37275),
            .I(sDAC_mem_pointerZ0Z_6));
    InMux I__7327 (
            .O(N__37272),
            .I(N__37269));
    LocalMux I__7326 (
            .O(N__37269),
            .I(sDAC_mem_pointerZ0Z_7));
    CascadeMux I__7325 (
            .O(N__37266),
            .I(N__37262));
    InMux I__7324 (
            .O(N__37265),
            .I(N__37259));
    InMux I__7323 (
            .O(N__37262),
            .I(N__37256));
    LocalMux I__7322 (
            .O(N__37259),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1 ));
    LocalMux I__7321 (
            .O(N__37256),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1 ));
    InMux I__7320 (
            .O(N__37251),
            .I(N__37248));
    LocalMux I__7319 (
            .O(N__37248),
            .I(N__37245));
    Span4Mux_h I__7318 (
            .O(N__37245),
            .I(N__37241));
    CascadeMux I__7317 (
            .O(N__37244),
            .I(N__37237));
    Span4Mux_v I__7316 (
            .O(N__37241),
            .I(N__37234));
    InMux I__7315 (
            .O(N__37240),
            .I(N__37231));
    InMux I__7314 (
            .O(N__37237),
            .I(N__37228));
    Odrv4 I__7313 (
            .O(N__37234),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0 ));
    LocalMux I__7312 (
            .O(N__37231),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0 ));
    LocalMux I__7311 (
            .O(N__37228),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0 ));
    InMux I__7310 (
            .O(N__37221),
            .I(N__37215));
    InMux I__7309 (
            .O(N__37220),
            .I(N__37215));
    LocalMux I__7308 (
            .O(N__37215),
            .I(N__37212));
    Span4Mux_h I__7307 (
            .O(N__37212),
            .I(N__37209));
    Span4Mux_v I__7306 (
            .O(N__37209),
            .I(N__37204));
    InMux I__7305 (
            .O(N__37208),
            .I(N__37201));
    InMux I__7304 (
            .O(N__37207),
            .I(N__37198));
    Odrv4 I__7303 (
            .O(N__37204),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1 ));
    LocalMux I__7302 (
            .O(N__37201),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1 ));
    LocalMux I__7301 (
            .O(N__37198),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1 ));
    InMux I__7300 (
            .O(N__37191),
            .I(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0 ));
    CascadeMux I__7299 (
            .O(N__37188),
            .I(N__37182));
    InMux I__7298 (
            .O(N__37187),
            .I(N__37177));
    InMux I__7297 (
            .O(N__37186),
            .I(N__37177));
    InMux I__7296 (
            .O(N__37185),
            .I(N__37174));
    InMux I__7295 (
            .O(N__37182),
            .I(N__37171));
    LocalMux I__7294 (
            .O(N__37177),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_i6 ));
    LocalMux I__7293 (
            .O(N__37174),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_i6 ));
    LocalMux I__7292 (
            .O(N__37171),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_i6 ));
    InMux I__7291 (
            .O(N__37164),
            .I(N__37157));
    InMux I__7290 (
            .O(N__37163),
            .I(N__37157));
    InMux I__7289 (
            .O(N__37162),
            .I(N__37154));
    LocalMux I__7288 (
            .O(N__37157),
            .I(N__37148));
    LocalMux I__7287 (
            .O(N__37154),
            .I(N__37148));
    InMux I__7286 (
            .O(N__37153),
            .I(N__37145));
    Span4Mux_v I__7285 (
            .O(N__37148),
            .I(N__37140));
    LocalMux I__7284 (
            .O(N__37145),
            .I(N__37140));
    Span4Mux_h I__7283 (
            .O(N__37140),
            .I(N__37135));
    InMux I__7282 (
            .O(N__37139),
            .I(N__37132));
    InMux I__7281 (
            .O(N__37138),
            .I(N__37129));
    Odrv4 I__7280 (
            .O(N__37135),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2 ));
    LocalMux I__7279 (
            .O(N__37132),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2 ));
    LocalMux I__7278 (
            .O(N__37129),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2 ));
    InMux I__7277 (
            .O(N__37122),
            .I(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1 ));
    InMux I__7276 (
            .O(N__37119),
            .I(N__37115));
    InMux I__7275 (
            .O(N__37118),
            .I(N__37112));
    LocalMux I__7274 (
            .O(N__37115),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3 ));
    LocalMux I__7273 (
            .O(N__37112),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3 ));
    InMux I__7272 (
            .O(N__37107),
            .I(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2 ));
    InMux I__7271 (
            .O(N__37104),
            .I(N__37100));
    InMux I__7270 (
            .O(N__37103),
            .I(N__37097));
    LocalMux I__7269 (
            .O(N__37100),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4 ));
    LocalMux I__7268 (
            .O(N__37097),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4 ));
    InMux I__7267 (
            .O(N__37092),
            .I(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3 ));
    CascadeMux I__7266 (
            .O(N__37089),
            .I(N__37084));
    InMux I__7265 (
            .O(N__37088),
            .I(N__37080));
    InMux I__7264 (
            .O(N__37087),
            .I(N__37076));
    InMux I__7263 (
            .O(N__37084),
            .I(N__37071));
    CascadeMux I__7262 (
            .O(N__37083),
            .I(N__37068));
    LocalMux I__7261 (
            .O(N__37080),
            .I(N__37065));
    InMux I__7260 (
            .O(N__37079),
            .I(N__37062));
    LocalMux I__7259 (
            .O(N__37076),
            .I(N__37059));
    InMux I__7258 (
            .O(N__37075),
            .I(N__37055));
    InMux I__7257 (
            .O(N__37074),
            .I(N__37050));
    LocalMux I__7256 (
            .O(N__37071),
            .I(N__37047));
    InMux I__7255 (
            .O(N__37068),
            .I(N__37044));
    Span4Mux_h I__7254 (
            .O(N__37065),
            .I(N__37039));
    LocalMux I__7253 (
            .O(N__37062),
            .I(N__37039));
    Span4Mux_v I__7252 (
            .O(N__37059),
            .I(N__37036));
    InMux I__7251 (
            .O(N__37058),
            .I(N__37033));
    LocalMux I__7250 (
            .O(N__37055),
            .I(N__37030));
    InMux I__7249 (
            .O(N__37054),
            .I(N__37027));
    InMux I__7248 (
            .O(N__37053),
            .I(N__37024));
    LocalMux I__7247 (
            .O(N__37050),
            .I(N__37021));
    Span4Mux_v I__7246 (
            .O(N__37047),
            .I(N__37016));
    LocalMux I__7245 (
            .O(N__37044),
            .I(N__37016));
    Span4Mux_v I__7244 (
            .O(N__37039),
            .I(N__37009));
    Span4Mux_h I__7243 (
            .O(N__37036),
            .I(N__37009));
    LocalMux I__7242 (
            .O(N__37033),
            .I(N__37009));
    Span4Mux_h I__7241 (
            .O(N__37030),
            .I(N__37006));
    LocalMux I__7240 (
            .O(N__37027),
            .I(un7_spon_23));
    LocalMux I__7239 (
            .O(N__37024),
            .I(un7_spon_23));
    Odrv12 I__7238 (
            .O(N__37021),
            .I(un7_spon_23));
    Odrv4 I__7237 (
            .O(N__37016),
            .I(un7_spon_23));
    Odrv4 I__7236 (
            .O(N__37009),
            .I(un7_spon_23));
    Odrv4 I__7235 (
            .O(N__37006),
            .I(un7_spon_23));
    InMux I__7234 (
            .O(N__36993),
            .I(N__36990));
    LocalMux I__7233 (
            .O(N__36990),
            .I(N__36987));
    Span4Mux_v I__7232 (
            .O(N__36987),
            .I(N__36984));
    Span4Mux_v I__7231 (
            .O(N__36984),
            .I(N__36981));
    Odrv4 I__7230 (
            .O(N__36981),
            .I(un17_sdacdyn_1));
    InMux I__7229 (
            .O(N__36978),
            .I(N__36975));
    LocalMux I__7228 (
            .O(N__36975),
            .I(N__36969));
    InMux I__7227 (
            .O(N__36974),
            .I(N__36964));
    InMux I__7226 (
            .O(N__36973),
            .I(N__36964));
    InMux I__7225 (
            .O(N__36972),
            .I(N__36961));
    Span4Mux_h I__7224 (
            .O(N__36969),
            .I(N__36952));
    LocalMux I__7223 (
            .O(N__36964),
            .I(N__36949));
    LocalMux I__7222 (
            .O(N__36961),
            .I(N__36946));
    InMux I__7221 (
            .O(N__36960),
            .I(N__36941));
    InMux I__7220 (
            .O(N__36959),
            .I(N__36941));
    InMux I__7219 (
            .O(N__36958),
            .I(N__36938));
    InMux I__7218 (
            .O(N__36957),
            .I(N__36935));
    InMux I__7217 (
            .O(N__36956),
            .I(N__36931));
    InMux I__7216 (
            .O(N__36955),
            .I(N__36928));
    Span4Mux_h I__7215 (
            .O(N__36952),
            .I(N__36925));
    Span4Mux_h I__7214 (
            .O(N__36949),
            .I(N__36922));
    Span4Mux_v I__7213 (
            .O(N__36946),
            .I(N__36917));
    LocalMux I__7212 (
            .O(N__36941),
            .I(N__36917));
    LocalMux I__7211 (
            .O(N__36938),
            .I(N__36914));
    LocalMux I__7210 (
            .O(N__36935),
            .I(N__36911));
    InMux I__7209 (
            .O(N__36934),
            .I(N__36908));
    LocalMux I__7208 (
            .O(N__36931),
            .I(N__36901));
    LocalMux I__7207 (
            .O(N__36928),
            .I(N__36901));
    Span4Mux_v I__7206 (
            .O(N__36925),
            .I(N__36901));
    Odrv4 I__7205 (
            .O(N__36922),
            .I(N_1479));
    Odrv4 I__7204 (
            .O(N__36917),
            .I(N_1479));
    Odrv4 I__7203 (
            .O(N__36914),
            .I(N_1479));
    Odrv4 I__7202 (
            .O(N__36911),
            .I(N_1479));
    LocalMux I__7201 (
            .O(N__36908),
            .I(N_1479));
    Odrv4 I__7200 (
            .O(N__36901),
            .I(N_1479));
    CascadeMux I__7199 (
            .O(N__36888),
            .I(N__36885));
    InMux I__7198 (
            .O(N__36885),
            .I(N__36879));
    CascadeMux I__7197 (
            .O(N__36884),
            .I(N__36874));
    CascadeMux I__7196 (
            .O(N__36883),
            .I(N__36870));
    CascadeMux I__7195 (
            .O(N__36882),
            .I(N__36867));
    LocalMux I__7194 (
            .O(N__36879),
            .I(N__36864));
    CascadeMux I__7193 (
            .O(N__36878),
            .I(N__36861));
    InMux I__7192 (
            .O(N__36877),
            .I(N__36856));
    InMux I__7191 (
            .O(N__36874),
            .I(N__36852));
    CascadeMux I__7190 (
            .O(N__36873),
            .I(N__36849));
    InMux I__7189 (
            .O(N__36870),
            .I(N__36845));
    InMux I__7188 (
            .O(N__36867),
            .I(N__36841));
    Span4Mux_v I__7187 (
            .O(N__36864),
            .I(N__36837));
    InMux I__7186 (
            .O(N__36861),
            .I(N__36832));
    InMux I__7185 (
            .O(N__36860),
            .I(N__36832));
    InMux I__7184 (
            .O(N__36859),
            .I(N__36829));
    LocalMux I__7183 (
            .O(N__36856),
            .I(N__36826));
    InMux I__7182 (
            .O(N__36855),
            .I(N__36823));
    LocalMux I__7181 (
            .O(N__36852),
            .I(N__36820));
    InMux I__7180 (
            .O(N__36849),
            .I(N__36814));
    InMux I__7179 (
            .O(N__36848),
            .I(N__36814));
    LocalMux I__7178 (
            .O(N__36845),
            .I(N__36810));
    InMux I__7177 (
            .O(N__36844),
            .I(N__36807));
    LocalMux I__7176 (
            .O(N__36841),
            .I(N__36801));
    InMux I__7175 (
            .O(N__36840),
            .I(N__36798));
    Span4Mux_h I__7174 (
            .O(N__36837),
            .I(N__36795));
    LocalMux I__7173 (
            .O(N__36832),
            .I(N__36786));
    LocalMux I__7172 (
            .O(N__36829),
            .I(N__36786));
    Span4Mux_v I__7171 (
            .O(N__36826),
            .I(N__36786));
    LocalMux I__7170 (
            .O(N__36823),
            .I(N__36786));
    Span4Mux_h I__7169 (
            .O(N__36820),
            .I(N__36783));
    InMux I__7168 (
            .O(N__36819),
            .I(N__36779));
    LocalMux I__7167 (
            .O(N__36814),
            .I(N__36776));
    InMux I__7166 (
            .O(N__36813),
            .I(N__36773));
    Span4Mux_h I__7165 (
            .O(N__36810),
            .I(N__36768));
    LocalMux I__7164 (
            .O(N__36807),
            .I(N__36768));
    InMux I__7163 (
            .O(N__36806),
            .I(N__36763));
    InMux I__7162 (
            .O(N__36805),
            .I(N__36763));
    InMux I__7161 (
            .O(N__36804),
            .I(N__36760));
    Span4Mux_v I__7160 (
            .O(N__36801),
            .I(N__36753));
    LocalMux I__7159 (
            .O(N__36798),
            .I(N__36753));
    Span4Mux_v I__7158 (
            .O(N__36795),
            .I(N__36753));
    Span4Mux_v I__7157 (
            .O(N__36786),
            .I(N__36748));
    Span4Mux_h I__7156 (
            .O(N__36783),
            .I(N__36748));
    InMux I__7155 (
            .O(N__36782),
            .I(N__36745));
    LocalMux I__7154 (
            .O(N__36779),
            .I(N__36742));
    Odrv12 I__7153 (
            .O(N__36776),
            .I(un7_spon_4));
    LocalMux I__7152 (
            .O(N__36773),
            .I(un7_spon_4));
    Odrv4 I__7151 (
            .O(N__36768),
            .I(un7_spon_4));
    LocalMux I__7150 (
            .O(N__36763),
            .I(un7_spon_4));
    LocalMux I__7149 (
            .O(N__36760),
            .I(un7_spon_4));
    Odrv4 I__7148 (
            .O(N__36753),
            .I(un7_spon_4));
    Odrv4 I__7147 (
            .O(N__36748),
            .I(un7_spon_4));
    LocalMux I__7146 (
            .O(N__36745),
            .I(un7_spon_4));
    Odrv4 I__7145 (
            .O(N__36742),
            .I(un7_spon_4));
    InMux I__7144 (
            .O(N__36723),
            .I(bfn_14_19_0_));
    InMux I__7143 (
            .O(N__36720),
            .I(N__36717));
    LocalMux I__7142 (
            .O(N__36717),
            .I(N__36714));
    Span4Mux_v I__7141 (
            .O(N__36714),
            .I(N__36711));
    Odrv4 I__7140 (
            .O(N__36711),
            .I(sDAC_mem_24Z0Z_3));
    InMux I__7139 (
            .O(N__36708),
            .I(N__36705));
    LocalMux I__7138 (
            .O(N__36705),
            .I(N__36702));
    Span4Mux_v I__7137 (
            .O(N__36702),
            .I(N__36699));
    Odrv4 I__7136 (
            .O(N__36699),
            .I(sDAC_mem_24Z0Z_6));
    InMux I__7135 (
            .O(N__36696),
            .I(N__36693));
    LocalMux I__7134 (
            .O(N__36693),
            .I(N__36690));
    Span4Mux_v I__7133 (
            .O(N__36690),
            .I(N__36687));
    Span4Mux_v I__7132 (
            .O(N__36687),
            .I(N__36684));
    Odrv4 I__7131 (
            .O(N__36684),
            .I(sDAC_mem_17Z0Z_2));
    CascadeMux I__7130 (
            .O(N__36681),
            .I(N__36678));
    InMux I__7129 (
            .O(N__36678),
            .I(N__36675));
    LocalMux I__7128 (
            .O(N__36675),
            .I(N__36672));
    Span4Mux_v I__7127 (
            .O(N__36672),
            .I(N__36669));
    Span4Mux_v I__7126 (
            .O(N__36669),
            .I(N__36666));
    Span4Mux_v I__7125 (
            .O(N__36666),
            .I(N__36663));
    Odrv4 I__7124 (
            .O(N__36663),
            .I(sDAC_data_RNO_29Z0Z_5));
    InMux I__7123 (
            .O(N__36660),
            .I(N__36656));
    InMux I__7122 (
            .O(N__36659),
            .I(N__36650));
    LocalMux I__7121 (
            .O(N__36656),
            .I(N__36647));
    InMux I__7120 (
            .O(N__36655),
            .I(N__36644));
    InMux I__7119 (
            .O(N__36654),
            .I(N__36641));
    CascadeMux I__7118 (
            .O(N__36653),
            .I(N__36638));
    LocalMux I__7117 (
            .O(N__36650),
            .I(N__36634));
    Span4Mux_h I__7116 (
            .O(N__36647),
            .I(N__36630));
    LocalMux I__7115 (
            .O(N__36644),
            .I(N__36626));
    LocalMux I__7114 (
            .O(N__36641),
            .I(N__36623));
    InMux I__7113 (
            .O(N__36638),
            .I(N__36620));
    InMux I__7112 (
            .O(N__36637),
            .I(N__36617));
    Span12Mux_v I__7111 (
            .O(N__36634),
            .I(N__36613));
    InMux I__7110 (
            .O(N__36633),
            .I(N__36610));
    Span4Mux_h I__7109 (
            .O(N__36630),
            .I(N__36607));
    InMux I__7108 (
            .O(N__36629),
            .I(N__36604));
    Span4Mux_h I__7107 (
            .O(N__36626),
            .I(N__36599));
    Span4Mux_h I__7106 (
            .O(N__36623),
            .I(N__36599));
    LocalMux I__7105 (
            .O(N__36620),
            .I(N__36596));
    LocalMux I__7104 (
            .O(N__36617),
            .I(N__36593));
    InMux I__7103 (
            .O(N__36616),
            .I(N__36590));
    Odrv12 I__7102 (
            .O(N__36613),
            .I(un7_spon_15));
    LocalMux I__7101 (
            .O(N__36610),
            .I(un7_spon_15));
    Odrv4 I__7100 (
            .O(N__36607),
            .I(un7_spon_15));
    LocalMux I__7099 (
            .O(N__36604),
            .I(un7_spon_15));
    Odrv4 I__7098 (
            .O(N__36599),
            .I(un7_spon_15));
    Odrv4 I__7097 (
            .O(N__36596),
            .I(un7_spon_15));
    Odrv12 I__7096 (
            .O(N__36593),
            .I(un7_spon_15));
    LocalMux I__7095 (
            .O(N__36590),
            .I(un7_spon_15));
    InMux I__7094 (
            .O(N__36573),
            .I(N__36570));
    LocalMux I__7093 (
            .O(N__36570),
            .I(N__36566));
    InMux I__7092 (
            .O(N__36569),
            .I(N__36563));
    Span4Mux_v I__7091 (
            .O(N__36566),
            .I(N__36558));
    LocalMux I__7090 (
            .O(N__36563),
            .I(N__36558));
    Odrv4 I__7089 (
            .O(N__36558),
            .I(sEEACQZ0Z_15));
    CascadeMux I__7088 (
            .O(N__36555),
            .I(N__36552));
    InMux I__7087 (
            .O(N__36552),
            .I(N__36549));
    LocalMux I__7086 (
            .O(N__36549),
            .I(sEEACQ_i_15));
    CascadeMux I__7085 (
            .O(N__36546),
            .I(N__36542));
    CascadeMux I__7084 (
            .O(N__36545),
            .I(N__36538));
    InMux I__7083 (
            .O(N__36542),
            .I(N__36535));
    InMux I__7082 (
            .O(N__36541),
            .I(N__36532));
    InMux I__7081 (
            .O(N__36538),
            .I(N__36526));
    LocalMux I__7080 (
            .O(N__36535),
            .I(N__36522));
    LocalMux I__7079 (
            .O(N__36532),
            .I(N__36518));
    InMux I__7078 (
            .O(N__36531),
            .I(N__36514));
    InMux I__7077 (
            .O(N__36530),
            .I(N__36511));
    InMux I__7076 (
            .O(N__36529),
            .I(N__36508));
    LocalMux I__7075 (
            .O(N__36526),
            .I(N__36504));
    InMux I__7074 (
            .O(N__36525),
            .I(N__36501));
    Span4Mux_h I__7073 (
            .O(N__36522),
            .I(N__36498));
    InMux I__7072 (
            .O(N__36521),
            .I(N__36495));
    Span4Mux_v I__7071 (
            .O(N__36518),
            .I(N__36492));
    InMux I__7070 (
            .O(N__36517),
            .I(N__36489));
    LocalMux I__7069 (
            .O(N__36514),
            .I(N__36486));
    LocalMux I__7068 (
            .O(N__36511),
            .I(N__36483));
    LocalMux I__7067 (
            .O(N__36508),
            .I(N__36480));
    InMux I__7066 (
            .O(N__36507),
            .I(N__36477));
    Span4Mux_h I__7065 (
            .O(N__36504),
            .I(N__36472));
    LocalMux I__7064 (
            .O(N__36501),
            .I(N__36472));
    Span4Mux_v I__7063 (
            .O(N__36498),
            .I(N__36463));
    LocalMux I__7062 (
            .O(N__36495),
            .I(N__36463));
    Span4Mux_h I__7061 (
            .O(N__36492),
            .I(N__36463));
    LocalMux I__7060 (
            .O(N__36489),
            .I(N__36463));
    Span4Mux_v I__7059 (
            .O(N__36486),
            .I(N__36458));
    Span4Mux_v I__7058 (
            .O(N__36483),
            .I(N__36458));
    Span4Mux_v I__7057 (
            .O(N__36480),
            .I(N__36455));
    LocalMux I__7056 (
            .O(N__36477),
            .I(un7_spon_16));
    Odrv4 I__7055 (
            .O(N__36472),
            .I(un7_spon_16));
    Odrv4 I__7054 (
            .O(N__36463),
            .I(un7_spon_16));
    Odrv4 I__7053 (
            .O(N__36458),
            .I(un7_spon_16));
    Odrv4 I__7052 (
            .O(N__36455),
            .I(un7_spon_16));
    InMux I__7051 (
            .O(N__36444),
            .I(N__36438));
    CascadeMux I__7050 (
            .O(N__36443),
            .I(N__36435));
    InMux I__7049 (
            .O(N__36442),
            .I(N__36432));
    InMux I__7048 (
            .O(N__36441),
            .I(N__36427));
    LocalMux I__7047 (
            .O(N__36438),
            .I(N__36423));
    InMux I__7046 (
            .O(N__36435),
            .I(N__36420));
    LocalMux I__7045 (
            .O(N__36432),
            .I(N__36417));
    InMux I__7044 (
            .O(N__36431),
            .I(N__36413));
    InMux I__7043 (
            .O(N__36430),
            .I(N__36410));
    LocalMux I__7042 (
            .O(N__36427),
            .I(N__36407));
    InMux I__7041 (
            .O(N__36426),
            .I(N__36402));
    Span4Mux_h I__7040 (
            .O(N__36423),
            .I(N__36397));
    LocalMux I__7039 (
            .O(N__36420),
            .I(N__36397));
    Span4Mux_v I__7038 (
            .O(N__36417),
            .I(N__36394));
    InMux I__7037 (
            .O(N__36416),
            .I(N__36391));
    LocalMux I__7036 (
            .O(N__36413),
            .I(N__36388));
    LocalMux I__7035 (
            .O(N__36410),
            .I(N__36385));
    Span4Mux_v I__7034 (
            .O(N__36407),
            .I(N__36382));
    InMux I__7033 (
            .O(N__36406),
            .I(N__36379));
    InMux I__7032 (
            .O(N__36405),
            .I(N__36376));
    LocalMux I__7031 (
            .O(N__36402),
            .I(N__36373));
    Span4Mux_v I__7030 (
            .O(N__36397),
            .I(N__36366));
    Span4Mux_h I__7029 (
            .O(N__36394),
            .I(N__36366));
    LocalMux I__7028 (
            .O(N__36391),
            .I(N__36366));
    Span4Mux_v I__7027 (
            .O(N__36388),
            .I(N__36361));
    Span4Mux_h I__7026 (
            .O(N__36385),
            .I(N__36361));
    Odrv4 I__7025 (
            .O(N__36382),
            .I(un7_spon_17));
    LocalMux I__7024 (
            .O(N__36379),
            .I(un7_spon_17));
    LocalMux I__7023 (
            .O(N__36376),
            .I(un7_spon_17));
    Odrv12 I__7022 (
            .O(N__36373),
            .I(un7_spon_17));
    Odrv4 I__7021 (
            .O(N__36366),
            .I(un7_spon_17));
    Odrv4 I__7020 (
            .O(N__36361),
            .I(un7_spon_17));
    CascadeMux I__7019 (
            .O(N__36348),
            .I(N__36342));
    InMux I__7018 (
            .O(N__36347),
            .I(N__36339));
    CascadeMux I__7017 (
            .O(N__36346),
            .I(N__36336));
    InMux I__7016 (
            .O(N__36345),
            .I(N__36333));
    InMux I__7015 (
            .O(N__36342),
            .I(N__36329));
    LocalMux I__7014 (
            .O(N__36339),
            .I(N__36324));
    InMux I__7013 (
            .O(N__36336),
            .I(N__36320));
    LocalMux I__7012 (
            .O(N__36333),
            .I(N__36317));
    InMux I__7011 (
            .O(N__36332),
            .I(N__36314));
    LocalMux I__7010 (
            .O(N__36329),
            .I(N__36311));
    InMux I__7009 (
            .O(N__36328),
            .I(N__36306));
    InMux I__7008 (
            .O(N__36327),
            .I(N__36303));
    Span4Mux_v I__7007 (
            .O(N__36324),
            .I(N__36300));
    InMux I__7006 (
            .O(N__36323),
            .I(N__36297));
    LocalMux I__7005 (
            .O(N__36320),
            .I(N__36290));
    Span4Mux_v I__7004 (
            .O(N__36317),
            .I(N__36290));
    LocalMux I__7003 (
            .O(N__36314),
            .I(N__36290));
    Span4Mux_h I__7002 (
            .O(N__36311),
            .I(N__36287));
    InMux I__7001 (
            .O(N__36310),
            .I(N__36284));
    InMux I__7000 (
            .O(N__36309),
            .I(N__36281));
    LocalMux I__6999 (
            .O(N__36306),
            .I(N__36278));
    LocalMux I__6998 (
            .O(N__36303),
            .I(N__36271));
    Span4Mux_h I__6997 (
            .O(N__36300),
            .I(N__36271));
    LocalMux I__6996 (
            .O(N__36297),
            .I(N__36271));
    Span4Mux_h I__6995 (
            .O(N__36290),
            .I(N__36268));
    Odrv4 I__6994 (
            .O(N__36287),
            .I(un7_spon_18));
    LocalMux I__6993 (
            .O(N__36284),
            .I(un7_spon_18));
    LocalMux I__6992 (
            .O(N__36281),
            .I(un7_spon_18));
    Odrv4 I__6991 (
            .O(N__36278),
            .I(un7_spon_18));
    Odrv4 I__6990 (
            .O(N__36271),
            .I(un7_spon_18));
    Odrv4 I__6989 (
            .O(N__36268),
            .I(un7_spon_18));
    InMux I__6988 (
            .O(N__36255),
            .I(N__36248));
    InMux I__6987 (
            .O(N__36254),
            .I(N__36244));
    InMux I__6986 (
            .O(N__36253),
            .I(N__36241));
    InMux I__6985 (
            .O(N__36252),
            .I(N__36238));
    InMux I__6984 (
            .O(N__36251),
            .I(N__36235));
    LocalMux I__6983 (
            .O(N__36248),
            .I(N__36232));
    InMux I__6982 (
            .O(N__36247),
            .I(N__36225));
    LocalMux I__6981 (
            .O(N__36244),
            .I(N__36220));
    LocalMux I__6980 (
            .O(N__36241),
            .I(N__36220));
    LocalMux I__6979 (
            .O(N__36238),
            .I(N__36217));
    LocalMux I__6978 (
            .O(N__36235),
            .I(N__36214));
    Span4Mux_v I__6977 (
            .O(N__36232),
            .I(N__36211));
    InMux I__6976 (
            .O(N__36231),
            .I(N__36208));
    InMux I__6975 (
            .O(N__36230),
            .I(N__36205));
    InMux I__6974 (
            .O(N__36229),
            .I(N__36202));
    InMux I__6973 (
            .O(N__36228),
            .I(N__36199));
    LocalMux I__6972 (
            .O(N__36225),
            .I(N__36196));
    Span4Mux_h I__6971 (
            .O(N__36220),
            .I(N__36191));
    Span4Mux_h I__6970 (
            .O(N__36217),
            .I(N__36191));
    Span4Mux_v I__6969 (
            .O(N__36214),
            .I(N__36184));
    Span4Mux_h I__6968 (
            .O(N__36211),
            .I(N__36184));
    LocalMux I__6967 (
            .O(N__36208),
            .I(N__36184));
    LocalMux I__6966 (
            .O(N__36205),
            .I(un7_spon_19));
    LocalMux I__6965 (
            .O(N__36202),
            .I(un7_spon_19));
    LocalMux I__6964 (
            .O(N__36199),
            .I(un7_spon_19));
    Odrv4 I__6963 (
            .O(N__36196),
            .I(un7_spon_19));
    Odrv4 I__6962 (
            .O(N__36191),
            .I(un7_spon_19));
    Odrv4 I__6961 (
            .O(N__36184),
            .I(un7_spon_19));
    CascadeMux I__6960 (
            .O(N__36171),
            .I(N__36166));
    InMux I__6959 (
            .O(N__36170),
            .I(N__36163));
    CascadeMux I__6958 (
            .O(N__36169),
            .I(N__36159));
    InMux I__6957 (
            .O(N__36166),
            .I(N__36155));
    LocalMux I__6956 (
            .O(N__36163),
            .I(N__36152));
    InMux I__6955 (
            .O(N__36162),
            .I(N__36149));
    InMux I__6954 (
            .O(N__36159),
            .I(N__36141));
    InMux I__6953 (
            .O(N__36158),
            .I(N__36141));
    LocalMux I__6952 (
            .O(N__36155),
            .I(N__36138));
    Span4Mux_h I__6951 (
            .O(N__36152),
            .I(N__36133));
    LocalMux I__6950 (
            .O(N__36149),
            .I(N__36130));
    InMux I__6949 (
            .O(N__36148),
            .I(N__36125));
    InMux I__6948 (
            .O(N__36147),
            .I(N__36125));
    InMux I__6947 (
            .O(N__36146),
            .I(N__36122));
    LocalMux I__6946 (
            .O(N__36141),
            .I(N__36119));
    Span4Mux_v I__6945 (
            .O(N__36138),
            .I(N__36116));
    InMux I__6944 (
            .O(N__36137),
            .I(N__36113));
    InMux I__6943 (
            .O(N__36136),
            .I(N__36110));
    Span4Mux_h I__6942 (
            .O(N__36133),
            .I(N__36107));
    Span4Mux_v I__6941 (
            .O(N__36130),
            .I(N__36102));
    LocalMux I__6940 (
            .O(N__36125),
            .I(N__36102));
    LocalMux I__6939 (
            .O(N__36122),
            .I(N__36099));
    Span4Mux_h I__6938 (
            .O(N__36119),
            .I(N__36096));
    Odrv4 I__6937 (
            .O(N__36116),
            .I(un7_spon_20));
    LocalMux I__6936 (
            .O(N__36113),
            .I(un7_spon_20));
    LocalMux I__6935 (
            .O(N__36110),
            .I(un7_spon_20));
    Odrv4 I__6934 (
            .O(N__36107),
            .I(un7_spon_20));
    Odrv4 I__6933 (
            .O(N__36102),
            .I(un7_spon_20));
    Odrv12 I__6932 (
            .O(N__36099),
            .I(un7_spon_20));
    Odrv4 I__6931 (
            .O(N__36096),
            .I(un7_spon_20));
    InMux I__6930 (
            .O(N__36081),
            .I(N__36076));
    CascadeMux I__6929 (
            .O(N__36080),
            .I(N__36073));
    InMux I__6928 (
            .O(N__36079),
            .I(N__36069));
    LocalMux I__6927 (
            .O(N__36076),
            .I(N__36066));
    InMux I__6926 (
            .O(N__36073),
            .I(N__36060));
    InMux I__6925 (
            .O(N__36072),
            .I(N__36057));
    LocalMux I__6924 (
            .O(N__36069),
            .I(N__36054));
    Span4Mux_h I__6923 (
            .O(N__36066),
            .I(N__36050));
    InMux I__6922 (
            .O(N__36065),
            .I(N__36047));
    InMux I__6921 (
            .O(N__36064),
            .I(N__36044));
    InMux I__6920 (
            .O(N__36063),
            .I(N__36041));
    LocalMux I__6919 (
            .O(N__36060),
            .I(N__36038));
    LocalMux I__6918 (
            .O(N__36057),
            .I(N__36035));
    Span4Mux_v I__6917 (
            .O(N__36054),
            .I(N__36032));
    InMux I__6916 (
            .O(N__36053),
            .I(N__36029));
    Span4Mux_h I__6915 (
            .O(N__36050),
            .I(N__36026));
    LocalMux I__6914 (
            .O(N__36047),
            .I(N__36023));
    LocalMux I__6913 (
            .O(N__36044),
            .I(N__36018));
    LocalMux I__6912 (
            .O(N__36041),
            .I(N__36018));
    Span4Mux_h I__6911 (
            .O(N__36038),
            .I(N__36013));
    Span4Mux_h I__6910 (
            .O(N__36035),
            .I(N__36013));
    Odrv4 I__6909 (
            .O(N__36032),
            .I(un7_spon_21));
    LocalMux I__6908 (
            .O(N__36029),
            .I(un7_spon_21));
    Odrv4 I__6907 (
            .O(N__36026),
            .I(un7_spon_21));
    Odrv4 I__6906 (
            .O(N__36023),
            .I(un7_spon_21));
    Odrv12 I__6905 (
            .O(N__36018),
            .I(un7_spon_21));
    Odrv4 I__6904 (
            .O(N__36013),
            .I(un7_spon_21));
    CascadeMux I__6903 (
            .O(N__36000),
            .I(N__35997));
    InMux I__6902 (
            .O(N__35997),
            .I(N__35991));
    CascadeMux I__6901 (
            .O(N__35996),
            .I(N__35988));
    CascadeMux I__6900 (
            .O(N__35995),
            .I(N__35985));
    InMux I__6899 (
            .O(N__35994),
            .I(N__35982));
    LocalMux I__6898 (
            .O(N__35991),
            .I(N__35976));
    InMux I__6897 (
            .O(N__35988),
            .I(N__35973));
    InMux I__6896 (
            .O(N__35985),
            .I(N__35970));
    LocalMux I__6895 (
            .O(N__35982),
            .I(N__35967));
    InMux I__6894 (
            .O(N__35981),
            .I(N__35964));
    CascadeMux I__6893 (
            .O(N__35980),
            .I(N__35961));
    CascadeMux I__6892 (
            .O(N__35979),
            .I(N__35957));
    Span4Mux_h I__6891 (
            .O(N__35976),
            .I(N__35952));
    LocalMux I__6890 (
            .O(N__35973),
            .I(N__35952));
    LocalMux I__6889 (
            .O(N__35970),
            .I(N__35947));
    Span4Mux_h I__6888 (
            .O(N__35967),
            .I(N__35944));
    LocalMux I__6887 (
            .O(N__35964),
            .I(N__35941));
    InMux I__6886 (
            .O(N__35961),
            .I(N__35938));
    InMux I__6885 (
            .O(N__35960),
            .I(N__35935));
    InMux I__6884 (
            .O(N__35957),
            .I(N__35932));
    Span4Mux_v I__6883 (
            .O(N__35952),
            .I(N__35929));
    InMux I__6882 (
            .O(N__35951),
            .I(N__35926));
    InMux I__6881 (
            .O(N__35950),
            .I(N__35923));
    Span4Mux_v I__6880 (
            .O(N__35947),
            .I(N__35920));
    Span4Mux_h I__6879 (
            .O(N__35944),
            .I(N__35917));
    Span4Mux_v I__6878 (
            .O(N__35941),
            .I(N__35912));
    LocalMux I__6877 (
            .O(N__35938),
            .I(N__35912));
    LocalMux I__6876 (
            .O(N__35935),
            .I(N__35909));
    LocalMux I__6875 (
            .O(N__35932),
            .I(N__35906));
    Odrv4 I__6874 (
            .O(N__35929),
            .I(un7_spon_22));
    LocalMux I__6873 (
            .O(N__35926),
            .I(un7_spon_22));
    LocalMux I__6872 (
            .O(N__35923),
            .I(un7_spon_22));
    Odrv4 I__6871 (
            .O(N__35920),
            .I(un7_spon_22));
    Odrv4 I__6870 (
            .O(N__35917),
            .I(un7_spon_22));
    Odrv4 I__6869 (
            .O(N__35912),
            .I(un7_spon_22));
    Odrv12 I__6868 (
            .O(N__35909),
            .I(un7_spon_22));
    Odrv12 I__6867 (
            .O(N__35906),
            .I(un7_spon_22));
    CascadeMux I__6866 (
            .O(N__35889),
            .I(N__35885));
    CascadeMux I__6865 (
            .O(N__35888),
            .I(N__35882));
    InMux I__6864 (
            .O(N__35885),
            .I(N__35878));
    InMux I__6863 (
            .O(N__35882),
            .I(N__35874));
    CascadeMux I__6862 (
            .O(N__35881),
            .I(N__35871));
    LocalMux I__6861 (
            .O(N__35878),
            .I(N__35867));
    InMux I__6860 (
            .O(N__35877),
            .I(N__35864));
    LocalMux I__6859 (
            .O(N__35874),
            .I(N__35861));
    InMux I__6858 (
            .O(N__35871),
            .I(N__35858));
    InMux I__6857 (
            .O(N__35870),
            .I(N__35854));
    Span4Mux_h I__6856 (
            .O(N__35867),
            .I(N__35851));
    LocalMux I__6855 (
            .O(N__35864),
            .I(N__35846));
    Span4Mux_h I__6854 (
            .O(N__35861),
            .I(N__35843));
    LocalMux I__6853 (
            .O(N__35858),
            .I(N__35839));
    InMux I__6852 (
            .O(N__35857),
            .I(N__35836));
    LocalMux I__6851 (
            .O(N__35854),
            .I(N__35833));
    Span4Mux_v I__6850 (
            .O(N__35851),
            .I(N__35830));
    InMux I__6849 (
            .O(N__35850),
            .I(N__35827));
    InMux I__6848 (
            .O(N__35849),
            .I(N__35824));
    Span4Mux_v I__6847 (
            .O(N__35846),
            .I(N__35819));
    Span4Mux_h I__6846 (
            .O(N__35843),
            .I(N__35819));
    InMux I__6845 (
            .O(N__35842),
            .I(N__35816));
    Span4Mux_h I__6844 (
            .O(N__35839),
            .I(N__35811));
    LocalMux I__6843 (
            .O(N__35836),
            .I(N__35811));
    Span4Mux_v I__6842 (
            .O(N__35833),
            .I(N__35808));
    Odrv4 I__6841 (
            .O(N__35830),
            .I(un7_spon_8));
    LocalMux I__6840 (
            .O(N__35827),
            .I(un7_spon_8));
    LocalMux I__6839 (
            .O(N__35824),
            .I(un7_spon_8));
    Odrv4 I__6838 (
            .O(N__35819),
            .I(un7_spon_8));
    LocalMux I__6837 (
            .O(N__35816),
            .I(un7_spon_8));
    Odrv4 I__6836 (
            .O(N__35811),
            .I(un7_spon_8));
    Odrv4 I__6835 (
            .O(N__35808),
            .I(un7_spon_8));
    InMux I__6834 (
            .O(N__35793),
            .I(N__35789));
    InMux I__6833 (
            .O(N__35792),
            .I(N__35786));
    LocalMux I__6832 (
            .O(N__35789),
            .I(N__35783));
    LocalMux I__6831 (
            .O(N__35786),
            .I(N__35780));
    Odrv4 I__6830 (
            .O(N__35783),
            .I(sEEACQZ0Z_8));
    Odrv4 I__6829 (
            .O(N__35780),
            .I(sEEACQZ0Z_8));
    InMux I__6828 (
            .O(N__35775),
            .I(N__35772));
    LocalMux I__6827 (
            .O(N__35772),
            .I(sEEACQ_i_8));
    InMux I__6826 (
            .O(N__35769),
            .I(N__35764));
    InMux I__6825 (
            .O(N__35768),
            .I(N__35758));
    InMux I__6824 (
            .O(N__35767),
            .I(N__35755));
    LocalMux I__6823 (
            .O(N__35764),
            .I(N__35752));
    InMux I__6822 (
            .O(N__35763),
            .I(N__35749));
    InMux I__6821 (
            .O(N__35762),
            .I(N__35746));
    CascadeMux I__6820 (
            .O(N__35761),
            .I(N__35743));
    LocalMux I__6819 (
            .O(N__35758),
            .I(N__35740));
    LocalMux I__6818 (
            .O(N__35755),
            .I(N__35735));
    Span4Mux_v I__6817 (
            .O(N__35752),
            .I(N__35732));
    LocalMux I__6816 (
            .O(N__35749),
            .I(N__35728));
    LocalMux I__6815 (
            .O(N__35746),
            .I(N__35725));
    InMux I__6814 (
            .O(N__35743),
            .I(N__35722));
    Span4Mux_v I__6813 (
            .O(N__35740),
            .I(N__35719));
    InMux I__6812 (
            .O(N__35739),
            .I(N__35716));
    InMux I__6811 (
            .O(N__35738),
            .I(N__35713));
    Span4Mux_v I__6810 (
            .O(N__35735),
            .I(N__35708));
    Span4Mux_h I__6809 (
            .O(N__35732),
            .I(N__35708));
    InMux I__6808 (
            .O(N__35731),
            .I(N__35705));
    Span4Mux_h I__6807 (
            .O(N__35728),
            .I(N__35698));
    Span4Mux_h I__6806 (
            .O(N__35725),
            .I(N__35698));
    LocalMux I__6805 (
            .O(N__35722),
            .I(N__35698));
    Span4Mux_h I__6804 (
            .O(N__35719),
            .I(N__35695));
    LocalMux I__6803 (
            .O(N__35716),
            .I(un7_spon_9));
    LocalMux I__6802 (
            .O(N__35713),
            .I(un7_spon_9));
    Odrv4 I__6801 (
            .O(N__35708),
            .I(un7_spon_9));
    LocalMux I__6800 (
            .O(N__35705),
            .I(un7_spon_9));
    Odrv4 I__6799 (
            .O(N__35698),
            .I(un7_spon_9));
    Odrv4 I__6798 (
            .O(N__35695),
            .I(un7_spon_9));
    InMux I__6797 (
            .O(N__35682),
            .I(N__35678));
    InMux I__6796 (
            .O(N__35681),
            .I(N__35675));
    LocalMux I__6795 (
            .O(N__35678),
            .I(N__35672));
    LocalMux I__6794 (
            .O(N__35675),
            .I(N__35669));
    Odrv4 I__6793 (
            .O(N__35672),
            .I(sEEACQZ0Z_9));
    Odrv4 I__6792 (
            .O(N__35669),
            .I(sEEACQZ0Z_9));
    CascadeMux I__6791 (
            .O(N__35664),
            .I(N__35661));
    InMux I__6790 (
            .O(N__35661),
            .I(N__35658));
    LocalMux I__6789 (
            .O(N__35658),
            .I(sEEACQ_i_9));
    CascadeMux I__6788 (
            .O(N__35655),
            .I(N__35651));
    CascadeMux I__6787 (
            .O(N__35654),
            .I(N__35648));
    InMux I__6786 (
            .O(N__35651),
            .I(N__35643));
    InMux I__6785 (
            .O(N__35648),
            .I(N__35640));
    InMux I__6784 (
            .O(N__35647),
            .I(N__35637));
    InMux I__6783 (
            .O(N__35646),
            .I(N__35634));
    LocalMux I__6782 (
            .O(N__35643),
            .I(N__35628));
    LocalMux I__6781 (
            .O(N__35640),
            .I(N__35624));
    LocalMux I__6780 (
            .O(N__35637),
            .I(N__35621));
    LocalMux I__6779 (
            .O(N__35634),
            .I(N__35618));
    InMux I__6778 (
            .O(N__35633),
            .I(N__35614));
    InMux I__6777 (
            .O(N__35632),
            .I(N__35609));
    InMux I__6776 (
            .O(N__35631),
            .I(N__35609));
    Span4Mux_h I__6775 (
            .O(N__35628),
            .I(N__35606));
    InMux I__6774 (
            .O(N__35627),
            .I(N__35603));
    Span4Mux_h I__6773 (
            .O(N__35624),
            .I(N__35598));
    Span4Mux_h I__6772 (
            .O(N__35621),
            .I(N__35598));
    Span12Mux_s11_v I__6771 (
            .O(N__35618),
            .I(N__35595));
    InMux I__6770 (
            .O(N__35617),
            .I(N__35592));
    LocalMux I__6769 (
            .O(N__35614),
            .I(N__35589));
    LocalMux I__6768 (
            .O(N__35609),
            .I(N__35586));
    Odrv4 I__6767 (
            .O(N__35606),
            .I(un7_spon_10));
    LocalMux I__6766 (
            .O(N__35603),
            .I(un7_spon_10));
    Odrv4 I__6765 (
            .O(N__35598),
            .I(un7_spon_10));
    Odrv12 I__6764 (
            .O(N__35595),
            .I(un7_spon_10));
    LocalMux I__6763 (
            .O(N__35592),
            .I(un7_spon_10));
    Odrv4 I__6762 (
            .O(N__35589),
            .I(un7_spon_10));
    Odrv4 I__6761 (
            .O(N__35586),
            .I(un7_spon_10));
    InMux I__6760 (
            .O(N__35571),
            .I(N__35568));
    LocalMux I__6759 (
            .O(N__35568),
            .I(N__35564));
    InMux I__6758 (
            .O(N__35567),
            .I(N__35561));
    Span4Mux_h I__6757 (
            .O(N__35564),
            .I(N__35558));
    LocalMux I__6756 (
            .O(N__35561),
            .I(N__35555));
    Odrv4 I__6755 (
            .O(N__35558),
            .I(sEEACQZ0Z_10));
    Odrv12 I__6754 (
            .O(N__35555),
            .I(sEEACQZ0Z_10));
    CascadeMux I__6753 (
            .O(N__35550),
            .I(N__35547));
    InMux I__6752 (
            .O(N__35547),
            .I(N__35544));
    LocalMux I__6751 (
            .O(N__35544),
            .I(sEEACQ_i_10));
    InMux I__6750 (
            .O(N__35541),
            .I(N__35537));
    InMux I__6749 (
            .O(N__35540),
            .I(N__35533));
    LocalMux I__6748 (
            .O(N__35537),
            .I(N__35529));
    InMux I__6747 (
            .O(N__35536),
            .I(N__35526));
    LocalMux I__6746 (
            .O(N__35533),
            .I(N__35523));
    InMux I__6745 (
            .O(N__35532),
            .I(N__35517));
    Span4Mux_h I__6744 (
            .O(N__35529),
            .I(N__35511));
    LocalMux I__6743 (
            .O(N__35526),
            .I(N__35511));
    Span4Mux_v I__6742 (
            .O(N__35523),
            .I(N__35508));
    InMux I__6741 (
            .O(N__35522),
            .I(N__35503));
    InMux I__6740 (
            .O(N__35521),
            .I(N__35503));
    InMux I__6739 (
            .O(N__35520),
            .I(N__35500));
    LocalMux I__6738 (
            .O(N__35517),
            .I(N__35497));
    InMux I__6737 (
            .O(N__35516),
            .I(N__35493));
    Span4Mux_v I__6736 (
            .O(N__35511),
            .I(N__35488));
    Span4Mux_h I__6735 (
            .O(N__35508),
            .I(N__35488));
    LocalMux I__6734 (
            .O(N__35503),
            .I(N__35485));
    LocalMux I__6733 (
            .O(N__35500),
            .I(N__35482));
    Span4Mux_h I__6732 (
            .O(N__35497),
            .I(N__35479));
    InMux I__6731 (
            .O(N__35496),
            .I(N__35476));
    LocalMux I__6730 (
            .O(N__35493),
            .I(un7_spon_11));
    Odrv4 I__6729 (
            .O(N__35488),
            .I(un7_spon_11));
    Odrv4 I__6728 (
            .O(N__35485),
            .I(un7_spon_11));
    Odrv4 I__6727 (
            .O(N__35482),
            .I(un7_spon_11));
    Odrv4 I__6726 (
            .O(N__35479),
            .I(un7_spon_11));
    LocalMux I__6725 (
            .O(N__35476),
            .I(un7_spon_11));
    InMux I__6724 (
            .O(N__35463),
            .I(N__35459));
    InMux I__6723 (
            .O(N__35462),
            .I(N__35456));
    LocalMux I__6722 (
            .O(N__35459),
            .I(N__35453));
    LocalMux I__6721 (
            .O(N__35456),
            .I(N__35450));
    Odrv4 I__6720 (
            .O(N__35453),
            .I(sEEACQZ0Z_11));
    Odrv12 I__6719 (
            .O(N__35450),
            .I(sEEACQZ0Z_11));
    CascadeMux I__6718 (
            .O(N__35445),
            .I(N__35442));
    InMux I__6717 (
            .O(N__35442),
            .I(N__35439));
    LocalMux I__6716 (
            .O(N__35439),
            .I(sEEACQ_i_11));
    InMux I__6715 (
            .O(N__35436),
            .I(N__35432));
    InMux I__6714 (
            .O(N__35435),
            .I(N__35429));
    LocalMux I__6713 (
            .O(N__35432),
            .I(N__35426));
    LocalMux I__6712 (
            .O(N__35429),
            .I(N__35423));
    Odrv4 I__6711 (
            .O(N__35426),
            .I(sEEACQZ0Z_12));
    Odrv12 I__6710 (
            .O(N__35423),
            .I(sEEACQZ0Z_12));
    CascadeMux I__6709 (
            .O(N__35418),
            .I(N__35415));
    InMux I__6708 (
            .O(N__35415),
            .I(N__35411));
    CascadeMux I__6707 (
            .O(N__35414),
            .I(N__35406));
    LocalMux I__6706 (
            .O(N__35411),
            .I(N__35403));
    InMux I__6705 (
            .O(N__35410),
            .I(N__35400));
    InMux I__6704 (
            .O(N__35409),
            .I(N__35397));
    InMux I__6703 (
            .O(N__35406),
            .I(N__35393));
    Span4Mux_h I__6702 (
            .O(N__35403),
            .I(N__35388));
    LocalMux I__6701 (
            .O(N__35400),
            .I(N__35388));
    LocalMux I__6700 (
            .O(N__35397),
            .I(N__35385));
    CascadeMux I__6699 (
            .O(N__35396),
            .I(N__35381));
    LocalMux I__6698 (
            .O(N__35393),
            .I(N__35376));
    Span4Mux_h I__6697 (
            .O(N__35388),
            .I(N__35373));
    Span4Mux_h I__6696 (
            .O(N__35385),
            .I(N__35370));
    InMux I__6695 (
            .O(N__35384),
            .I(N__35366));
    InMux I__6694 (
            .O(N__35381),
            .I(N__35361));
    InMux I__6693 (
            .O(N__35380),
            .I(N__35361));
    InMux I__6692 (
            .O(N__35379),
            .I(N__35358));
    Span4Mux_v I__6691 (
            .O(N__35376),
            .I(N__35353));
    Span4Mux_v I__6690 (
            .O(N__35373),
            .I(N__35353));
    Span4Mux_h I__6689 (
            .O(N__35370),
            .I(N__35350));
    InMux I__6688 (
            .O(N__35369),
            .I(N__35347));
    LocalMux I__6687 (
            .O(N__35366),
            .I(N__35344));
    LocalMux I__6686 (
            .O(N__35361),
            .I(N__35341));
    LocalMux I__6685 (
            .O(N__35358),
            .I(un7_spon_12));
    Odrv4 I__6684 (
            .O(N__35353),
            .I(un7_spon_12));
    Odrv4 I__6683 (
            .O(N__35350),
            .I(un7_spon_12));
    LocalMux I__6682 (
            .O(N__35347),
            .I(un7_spon_12));
    Odrv4 I__6681 (
            .O(N__35344),
            .I(un7_spon_12));
    Odrv4 I__6680 (
            .O(N__35341),
            .I(un7_spon_12));
    CascadeMux I__6679 (
            .O(N__35328),
            .I(N__35325));
    InMux I__6678 (
            .O(N__35325),
            .I(N__35322));
    LocalMux I__6677 (
            .O(N__35322),
            .I(sEEACQ_i_12));
    CascadeMux I__6676 (
            .O(N__35319),
            .I(N__35316));
    InMux I__6675 (
            .O(N__35316),
            .I(N__35312));
    InMux I__6674 (
            .O(N__35315),
            .I(N__35307));
    LocalMux I__6673 (
            .O(N__35312),
            .I(N__35303));
    InMux I__6672 (
            .O(N__35311),
            .I(N__35299));
    CascadeMux I__6671 (
            .O(N__35310),
            .I(N__35295));
    LocalMux I__6670 (
            .O(N__35307),
            .I(N__35292));
    InMux I__6669 (
            .O(N__35306),
            .I(N__35288));
    Span4Mux_h I__6668 (
            .O(N__35303),
            .I(N__35285));
    InMux I__6667 (
            .O(N__35302),
            .I(N__35281));
    LocalMux I__6666 (
            .O(N__35299),
            .I(N__35278));
    InMux I__6665 (
            .O(N__35298),
            .I(N__35273));
    InMux I__6664 (
            .O(N__35295),
            .I(N__35273));
    Span4Mux_v I__6663 (
            .O(N__35292),
            .I(N__35270));
    InMux I__6662 (
            .O(N__35291),
            .I(N__35267));
    LocalMux I__6661 (
            .O(N__35288),
            .I(N__35264));
    Span4Mux_h I__6660 (
            .O(N__35285),
            .I(N__35261));
    InMux I__6659 (
            .O(N__35284),
            .I(N__35258));
    LocalMux I__6658 (
            .O(N__35281),
            .I(N__35255));
    Span4Mux_h I__6657 (
            .O(N__35278),
            .I(N__35250));
    LocalMux I__6656 (
            .O(N__35273),
            .I(N__35250));
    Odrv4 I__6655 (
            .O(N__35270),
            .I(un7_spon_13));
    LocalMux I__6654 (
            .O(N__35267),
            .I(un7_spon_13));
    Odrv12 I__6653 (
            .O(N__35264),
            .I(un7_spon_13));
    Odrv4 I__6652 (
            .O(N__35261),
            .I(un7_spon_13));
    LocalMux I__6651 (
            .O(N__35258),
            .I(un7_spon_13));
    Odrv4 I__6650 (
            .O(N__35255),
            .I(un7_spon_13));
    Odrv4 I__6649 (
            .O(N__35250),
            .I(un7_spon_13));
    InMux I__6648 (
            .O(N__35235),
            .I(N__35232));
    LocalMux I__6647 (
            .O(N__35232),
            .I(N__35228));
    InMux I__6646 (
            .O(N__35231),
            .I(N__35225));
    Span4Mux_v I__6645 (
            .O(N__35228),
            .I(N__35222));
    LocalMux I__6644 (
            .O(N__35225),
            .I(N__35219));
    Odrv4 I__6643 (
            .O(N__35222),
            .I(sEEACQZ0Z_13));
    Odrv12 I__6642 (
            .O(N__35219),
            .I(sEEACQZ0Z_13));
    InMux I__6641 (
            .O(N__35214),
            .I(N__35211));
    LocalMux I__6640 (
            .O(N__35211),
            .I(sEEACQ_i_13));
    CascadeMux I__6639 (
            .O(N__35208),
            .I(N__35205));
    InMux I__6638 (
            .O(N__35205),
            .I(N__35199));
    CascadeMux I__6637 (
            .O(N__35204),
            .I(N__35196));
    InMux I__6636 (
            .O(N__35203),
            .I(N__35192));
    CascadeMux I__6635 (
            .O(N__35202),
            .I(N__35189));
    LocalMux I__6634 (
            .O(N__35199),
            .I(N__35185));
    InMux I__6633 (
            .O(N__35196),
            .I(N__35182));
    InMux I__6632 (
            .O(N__35195),
            .I(N__35179));
    LocalMux I__6631 (
            .O(N__35192),
            .I(N__35176));
    InMux I__6630 (
            .O(N__35189),
            .I(N__35173));
    InMux I__6629 (
            .O(N__35188),
            .I(N__35170));
    Span4Mux_h I__6628 (
            .O(N__35185),
            .I(N__35165));
    LocalMux I__6627 (
            .O(N__35182),
            .I(N__35165));
    LocalMux I__6626 (
            .O(N__35179),
            .I(N__35160));
    Span4Mux_h I__6625 (
            .O(N__35176),
            .I(N__35157));
    LocalMux I__6624 (
            .O(N__35173),
            .I(N__35153));
    LocalMux I__6623 (
            .O(N__35170),
            .I(N__35150));
    Span4Mux_v I__6622 (
            .O(N__35165),
            .I(N__35147));
    InMux I__6621 (
            .O(N__35164),
            .I(N__35144));
    InMux I__6620 (
            .O(N__35163),
            .I(N__35141));
    Span4Mux_v I__6619 (
            .O(N__35160),
            .I(N__35136));
    Span4Mux_h I__6618 (
            .O(N__35157),
            .I(N__35136));
    InMux I__6617 (
            .O(N__35156),
            .I(N__35133));
    Span4Mux_v I__6616 (
            .O(N__35153),
            .I(N__35128));
    Span4Mux_h I__6615 (
            .O(N__35150),
            .I(N__35128));
    Odrv4 I__6614 (
            .O(N__35147),
            .I(un7_spon_14));
    LocalMux I__6613 (
            .O(N__35144),
            .I(un7_spon_14));
    LocalMux I__6612 (
            .O(N__35141),
            .I(un7_spon_14));
    Odrv4 I__6611 (
            .O(N__35136),
            .I(un7_spon_14));
    LocalMux I__6610 (
            .O(N__35133),
            .I(un7_spon_14));
    Odrv4 I__6609 (
            .O(N__35128),
            .I(un7_spon_14));
    InMux I__6608 (
            .O(N__35115),
            .I(N__35112));
    LocalMux I__6607 (
            .O(N__35112),
            .I(N__35108));
    InMux I__6606 (
            .O(N__35111),
            .I(N__35105));
    Span4Mux_v I__6605 (
            .O(N__35108),
            .I(N__35100));
    LocalMux I__6604 (
            .O(N__35105),
            .I(N__35100));
    Odrv4 I__6603 (
            .O(N__35100),
            .I(sEEACQZ0Z_14));
    CascadeMux I__6602 (
            .O(N__35097),
            .I(N__35094));
    InMux I__6601 (
            .O(N__35094),
            .I(N__35091));
    LocalMux I__6600 (
            .O(N__35091),
            .I(sEEACQ_i_14));
    InMux I__6599 (
            .O(N__35088),
            .I(N__35085));
    LocalMux I__6598 (
            .O(N__35085),
            .I(sEEACQ_i_0));
    InMux I__6597 (
            .O(N__35082),
            .I(N__35079));
    LocalMux I__6596 (
            .O(N__35079),
            .I(N__35076));
    Span4Mux_v I__6595 (
            .O(N__35076),
            .I(N__35072));
    InMux I__6594 (
            .O(N__35075),
            .I(N__35069));
    Odrv4 I__6593 (
            .O(N__35072),
            .I(sEEACQZ0Z_1));
    LocalMux I__6592 (
            .O(N__35069),
            .I(sEEACQZ0Z_1));
    CascadeMux I__6591 (
            .O(N__35064),
            .I(N__35059));
    CascadeMux I__6590 (
            .O(N__35063),
            .I(N__35055));
    InMux I__6589 (
            .O(N__35062),
            .I(N__35052));
    InMux I__6588 (
            .O(N__35059),
            .I(N__35047));
    InMux I__6587 (
            .O(N__35058),
            .I(N__35044));
    InMux I__6586 (
            .O(N__35055),
            .I(N__35041));
    LocalMux I__6585 (
            .O(N__35052),
            .I(N__35038));
    InMux I__6584 (
            .O(N__35051),
            .I(N__35035));
    InMux I__6583 (
            .O(N__35050),
            .I(N__35031));
    LocalMux I__6582 (
            .O(N__35047),
            .I(N__35028));
    LocalMux I__6581 (
            .O(N__35044),
            .I(N__35025));
    LocalMux I__6580 (
            .O(N__35041),
            .I(N__35020));
    Span4Mux_v I__6579 (
            .O(N__35038),
            .I(N__35017));
    LocalMux I__6578 (
            .O(N__35035),
            .I(N__35014));
    InMux I__6577 (
            .O(N__35034),
            .I(N__35011));
    LocalMux I__6576 (
            .O(N__35031),
            .I(N__35008));
    Span4Mux_h I__6575 (
            .O(N__35028),
            .I(N__35003));
    Span4Mux_h I__6574 (
            .O(N__35025),
            .I(N__35003));
    InMux I__6573 (
            .O(N__35024),
            .I(N__35000));
    InMux I__6572 (
            .O(N__35023),
            .I(N__34997));
    Span4Mux_v I__6571 (
            .O(N__35020),
            .I(N__34990));
    Span4Mux_h I__6570 (
            .O(N__35017),
            .I(N__34990));
    Span4Mux_v I__6569 (
            .O(N__35014),
            .I(N__34990));
    LocalMux I__6568 (
            .O(N__35011),
            .I(un7_spon_1));
    Odrv4 I__6567 (
            .O(N__35008),
            .I(un7_spon_1));
    Odrv4 I__6566 (
            .O(N__35003),
            .I(un7_spon_1));
    LocalMux I__6565 (
            .O(N__35000),
            .I(un7_spon_1));
    LocalMux I__6564 (
            .O(N__34997),
            .I(un7_spon_1));
    Odrv4 I__6563 (
            .O(N__34990),
            .I(un7_spon_1));
    CascadeMux I__6562 (
            .O(N__34977),
            .I(N__34974));
    InMux I__6561 (
            .O(N__34974),
            .I(N__34971));
    LocalMux I__6560 (
            .O(N__34971),
            .I(sEEACQ_i_1));
    CascadeMux I__6559 (
            .O(N__34968),
            .I(N__34965));
    InMux I__6558 (
            .O(N__34965),
            .I(N__34961));
    CascadeMux I__6557 (
            .O(N__34964),
            .I(N__34958));
    LocalMux I__6556 (
            .O(N__34961),
            .I(N__34953));
    InMux I__6555 (
            .O(N__34958),
            .I(N__34950));
    InMux I__6554 (
            .O(N__34957),
            .I(N__34946));
    InMux I__6553 (
            .O(N__34956),
            .I(N__34943));
    Span4Mux_v I__6552 (
            .O(N__34953),
            .I(N__34936));
    LocalMux I__6551 (
            .O(N__34950),
            .I(N__34936));
    InMux I__6550 (
            .O(N__34949),
            .I(N__34933));
    LocalMux I__6549 (
            .O(N__34946),
            .I(N__34930));
    LocalMux I__6548 (
            .O(N__34943),
            .I(N__34926));
    InMux I__6547 (
            .O(N__34942),
            .I(N__34922));
    InMux I__6546 (
            .O(N__34941),
            .I(N__34919));
    Span4Mux_h I__6545 (
            .O(N__34936),
            .I(N__34914));
    LocalMux I__6544 (
            .O(N__34933),
            .I(N__34914));
    Span4Mux_h I__6543 (
            .O(N__34930),
            .I(N__34911));
    InMux I__6542 (
            .O(N__34929),
            .I(N__34908));
    Span12Mux_v I__6541 (
            .O(N__34926),
            .I(N__34905));
    InMux I__6540 (
            .O(N__34925),
            .I(N__34902));
    LocalMux I__6539 (
            .O(N__34922),
            .I(N__34899));
    LocalMux I__6538 (
            .O(N__34919),
            .I(un7_spon_2));
    Odrv4 I__6537 (
            .O(N__34914),
            .I(un7_spon_2));
    Odrv4 I__6536 (
            .O(N__34911),
            .I(un7_spon_2));
    LocalMux I__6535 (
            .O(N__34908),
            .I(un7_spon_2));
    Odrv12 I__6534 (
            .O(N__34905),
            .I(un7_spon_2));
    LocalMux I__6533 (
            .O(N__34902),
            .I(un7_spon_2));
    Odrv4 I__6532 (
            .O(N__34899),
            .I(un7_spon_2));
    InMux I__6531 (
            .O(N__34884),
            .I(N__34881));
    LocalMux I__6530 (
            .O(N__34881),
            .I(N__34878));
    Span4Mux_h I__6529 (
            .O(N__34878),
            .I(N__34874));
    InMux I__6528 (
            .O(N__34877),
            .I(N__34871));
    Odrv4 I__6527 (
            .O(N__34874),
            .I(sEEACQZ0Z_2));
    LocalMux I__6526 (
            .O(N__34871),
            .I(sEEACQZ0Z_2));
    CascadeMux I__6525 (
            .O(N__34866),
            .I(N__34863));
    InMux I__6524 (
            .O(N__34863),
            .I(N__34860));
    LocalMux I__6523 (
            .O(N__34860),
            .I(sEEACQ_i_2));
    InMux I__6522 (
            .O(N__34857),
            .I(N__34853));
    InMux I__6521 (
            .O(N__34856),
            .I(N__34848));
    LocalMux I__6520 (
            .O(N__34853),
            .I(N__34845));
    InMux I__6519 (
            .O(N__34852),
            .I(N__34842));
    InMux I__6518 (
            .O(N__34851),
            .I(N__34839));
    LocalMux I__6517 (
            .O(N__34848),
            .I(N__34836));
    Span4Mux_h I__6516 (
            .O(N__34845),
            .I(N__34828));
    LocalMux I__6515 (
            .O(N__34842),
            .I(N__34828));
    LocalMux I__6514 (
            .O(N__34839),
            .I(N__34824));
    Span4Mux_v I__6513 (
            .O(N__34836),
            .I(N__34821));
    InMux I__6512 (
            .O(N__34835),
            .I(N__34818));
    InMux I__6511 (
            .O(N__34834),
            .I(N__34814));
    InMux I__6510 (
            .O(N__34833),
            .I(N__34811));
    Span4Mux_h I__6509 (
            .O(N__34828),
            .I(N__34808));
    InMux I__6508 (
            .O(N__34827),
            .I(N__34805));
    Span4Mux_v I__6507 (
            .O(N__34824),
            .I(N__34800));
    Span4Mux_h I__6506 (
            .O(N__34821),
            .I(N__34800));
    LocalMux I__6505 (
            .O(N__34818),
            .I(N__34797));
    InMux I__6504 (
            .O(N__34817),
            .I(N__34794));
    LocalMux I__6503 (
            .O(N__34814),
            .I(un7_spon_3));
    LocalMux I__6502 (
            .O(N__34811),
            .I(un7_spon_3));
    Odrv4 I__6501 (
            .O(N__34808),
            .I(un7_spon_3));
    LocalMux I__6500 (
            .O(N__34805),
            .I(un7_spon_3));
    Odrv4 I__6499 (
            .O(N__34800),
            .I(un7_spon_3));
    Odrv4 I__6498 (
            .O(N__34797),
            .I(un7_spon_3));
    LocalMux I__6497 (
            .O(N__34794),
            .I(un7_spon_3));
    InMux I__6496 (
            .O(N__34779),
            .I(N__34776));
    LocalMux I__6495 (
            .O(N__34776),
            .I(N__34773));
    Span4Mux_h I__6494 (
            .O(N__34773),
            .I(N__34769));
    InMux I__6493 (
            .O(N__34772),
            .I(N__34766));
    Odrv4 I__6492 (
            .O(N__34769),
            .I(sEEACQZ0Z_3));
    LocalMux I__6491 (
            .O(N__34766),
            .I(sEEACQZ0Z_3));
    CascadeMux I__6490 (
            .O(N__34761),
            .I(N__34758));
    InMux I__6489 (
            .O(N__34758),
            .I(N__34755));
    LocalMux I__6488 (
            .O(N__34755),
            .I(sEEACQ_i_3));
    InMux I__6487 (
            .O(N__34752),
            .I(N__34749));
    LocalMux I__6486 (
            .O(N__34749),
            .I(N__34746));
    Span4Mux_h I__6485 (
            .O(N__34746),
            .I(N__34742));
    InMux I__6484 (
            .O(N__34745),
            .I(N__34739));
    Odrv4 I__6483 (
            .O(N__34742),
            .I(sEEACQZ0Z_4));
    LocalMux I__6482 (
            .O(N__34739),
            .I(sEEACQZ0Z_4));
    InMux I__6481 (
            .O(N__34734),
            .I(N__34731));
    LocalMux I__6480 (
            .O(N__34731),
            .I(sEEACQ_i_4));
    InMux I__6479 (
            .O(N__34728),
            .I(N__34723));
    CascadeMux I__6478 (
            .O(N__34727),
            .I(N__34720));
    InMux I__6477 (
            .O(N__34726),
            .I(N__34717));
    LocalMux I__6476 (
            .O(N__34723),
            .I(N__34714));
    InMux I__6475 (
            .O(N__34720),
            .I(N__34711));
    LocalMux I__6474 (
            .O(N__34717),
            .I(N__34707));
    Span4Mux_h I__6473 (
            .O(N__34714),
            .I(N__34701));
    LocalMux I__6472 (
            .O(N__34711),
            .I(N__34701));
    InMux I__6471 (
            .O(N__34710),
            .I(N__34696));
    Span4Mux_h I__6470 (
            .O(N__34707),
            .I(N__34692));
    InMux I__6469 (
            .O(N__34706),
            .I(N__34688));
    Span4Mux_v I__6468 (
            .O(N__34701),
            .I(N__34685));
    InMux I__6467 (
            .O(N__34700),
            .I(N__34682));
    InMux I__6466 (
            .O(N__34699),
            .I(N__34679));
    LocalMux I__6465 (
            .O(N__34696),
            .I(N__34676));
    InMux I__6464 (
            .O(N__34695),
            .I(N__34673));
    Span4Mux_h I__6463 (
            .O(N__34692),
            .I(N__34670));
    InMux I__6462 (
            .O(N__34691),
            .I(N__34667));
    LocalMux I__6461 (
            .O(N__34688),
            .I(N__34664));
    Odrv4 I__6460 (
            .O(N__34685),
            .I(un7_spon_5));
    LocalMux I__6459 (
            .O(N__34682),
            .I(un7_spon_5));
    LocalMux I__6458 (
            .O(N__34679),
            .I(un7_spon_5));
    Odrv12 I__6457 (
            .O(N__34676),
            .I(un7_spon_5));
    LocalMux I__6456 (
            .O(N__34673),
            .I(un7_spon_5));
    Odrv4 I__6455 (
            .O(N__34670),
            .I(un7_spon_5));
    LocalMux I__6454 (
            .O(N__34667),
            .I(un7_spon_5));
    Odrv4 I__6453 (
            .O(N__34664),
            .I(un7_spon_5));
    InMux I__6452 (
            .O(N__34647),
            .I(N__34644));
    LocalMux I__6451 (
            .O(N__34644),
            .I(N__34641));
    Span4Mux_v I__6450 (
            .O(N__34641),
            .I(N__34637));
    InMux I__6449 (
            .O(N__34640),
            .I(N__34634));
    Odrv4 I__6448 (
            .O(N__34637),
            .I(sEEACQZ0Z_5));
    LocalMux I__6447 (
            .O(N__34634),
            .I(sEEACQZ0Z_5));
    CascadeMux I__6446 (
            .O(N__34629),
            .I(N__34626));
    InMux I__6445 (
            .O(N__34626),
            .I(N__34623));
    LocalMux I__6444 (
            .O(N__34623),
            .I(sEEACQ_i_5));
    CascadeMux I__6443 (
            .O(N__34620),
            .I(N__34616));
    CascadeMux I__6442 (
            .O(N__34619),
            .I(N__34613));
    InMux I__6441 (
            .O(N__34616),
            .I(N__34609));
    InMux I__6440 (
            .O(N__34613),
            .I(N__34606));
    InMux I__6439 (
            .O(N__34612),
            .I(N__34602));
    LocalMux I__6438 (
            .O(N__34609),
            .I(N__34598));
    LocalMux I__6437 (
            .O(N__34606),
            .I(N__34595));
    InMux I__6436 (
            .O(N__34605),
            .I(N__34591));
    LocalMux I__6435 (
            .O(N__34602),
            .I(N__34588));
    InMux I__6434 (
            .O(N__34601),
            .I(N__34585));
    Span4Mux_v I__6433 (
            .O(N__34598),
            .I(N__34582));
    Span4Mux_v I__6432 (
            .O(N__34595),
            .I(N__34579));
    CascadeMux I__6431 (
            .O(N__34594),
            .I(N__34576));
    LocalMux I__6430 (
            .O(N__34591),
            .I(N__34571));
    Span4Mux_h I__6429 (
            .O(N__34588),
            .I(N__34568));
    LocalMux I__6428 (
            .O(N__34585),
            .I(N__34564));
    Span4Mux_v I__6427 (
            .O(N__34582),
            .I(N__34561));
    Span4Mux_v I__6426 (
            .O(N__34579),
            .I(N__34558));
    InMux I__6425 (
            .O(N__34576),
            .I(N__34555));
    InMux I__6424 (
            .O(N__34575),
            .I(N__34552));
    InMux I__6423 (
            .O(N__34574),
            .I(N__34549));
    Span4Mux_v I__6422 (
            .O(N__34571),
            .I(N__34544));
    Span4Mux_h I__6421 (
            .O(N__34568),
            .I(N__34544));
    InMux I__6420 (
            .O(N__34567),
            .I(N__34541));
    Span4Mux_h I__6419 (
            .O(N__34564),
            .I(N__34538));
    Odrv4 I__6418 (
            .O(N__34561),
            .I(un7_spon_6));
    Odrv4 I__6417 (
            .O(N__34558),
            .I(un7_spon_6));
    LocalMux I__6416 (
            .O(N__34555),
            .I(un7_spon_6));
    LocalMux I__6415 (
            .O(N__34552),
            .I(un7_spon_6));
    LocalMux I__6414 (
            .O(N__34549),
            .I(un7_spon_6));
    Odrv4 I__6413 (
            .O(N__34544),
            .I(un7_spon_6));
    LocalMux I__6412 (
            .O(N__34541),
            .I(un7_spon_6));
    Odrv4 I__6411 (
            .O(N__34538),
            .I(un7_spon_6));
    InMux I__6410 (
            .O(N__34521),
            .I(N__34518));
    LocalMux I__6409 (
            .O(N__34518),
            .I(N__34515));
    Span4Mux_v I__6408 (
            .O(N__34515),
            .I(N__34511));
    InMux I__6407 (
            .O(N__34514),
            .I(N__34508));
    Odrv4 I__6406 (
            .O(N__34511),
            .I(sEEACQZ0Z_6));
    LocalMux I__6405 (
            .O(N__34508),
            .I(sEEACQZ0Z_6));
    CascadeMux I__6404 (
            .O(N__34503),
            .I(N__34500));
    InMux I__6403 (
            .O(N__34500),
            .I(N__34497));
    LocalMux I__6402 (
            .O(N__34497),
            .I(sEEACQ_i_6));
    CascadeMux I__6401 (
            .O(N__34494),
            .I(N__34490));
    CascadeMux I__6400 (
            .O(N__34493),
            .I(N__34486));
    InMux I__6399 (
            .O(N__34490),
            .I(N__34483));
    CascadeMux I__6398 (
            .O(N__34489),
            .I(N__34480));
    InMux I__6397 (
            .O(N__34486),
            .I(N__34476));
    LocalMux I__6396 (
            .O(N__34483),
            .I(N__34472));
    InMux I__6395 (
            .O(N__34480),
            .I(N__34469));
    InMux I__6394 (
            .O(N__34479),
            .I(N__34466));
    LocalMux I__6393 (
            .O(N__34476),
            .I(N__34463));
    CascadeMux I__6392 (
            .O(N__34475),
            .I(N__34460));
    Span4Mux_h I__6391 (
            .O(N__34472),
            .I(N__34455));
    LocalMux I__6390 (
            .O(N__34469),
            .I(N__34455));
    LocalMux I__6389 (
            .O(N__34466),
            .I(N__34449));
    Span4Mux_h I__6388 (
            .O(N__34463),
            .I(N__34446));
    InMux I__6387 (
            .O(N__34460),
            .I(N__34442));
    Span4Mux_v I__6386 (
            .O(N__34455),
            .I(N__34439));
    InMux I__6385 (
            .O(N__34454),
            .I(N__34436));
    InMux I__6384 (
            .O(N__34453),
            .I(N__34433));
    InMux I__6383 (
            .O(N__34452),
            .I(N__34430));
    Span4Mux_v I__6382 (
            .O(N__34449),
            .I(N__34425));
    Span4Mux_h I__6381 (
            .O(N__34446),
            .I(N__34425));
    InMux I__6380 (
            .O(N__34445),
            .I(N__34422));
    LocalMux I__6379 (
            .O(N__34442),
            .I(N__34419));
    Odrv4 I__6378 (
            .O(N__34439),
            .I(un7_spon_7));
    LocalMux I__6377 (
            .O(N__34436),
            .I(un7_spon_7));
    LocalMux I__6376 (
            .O(N__34433),
            .I(un7_spon_7));
    LocalMux I__6375 (
            .O(N__34430),
            .I(un7_spon_7));
    Odrv4 I__6374 (
            .O(N__34425),
            .I(un7_spon_7));
    LocalMux I__6373 (
            .O(N__34422),
            .I(un7_spon_7));
    Odrv4 I__6372 (
            .O(N__34419),
            .I(un7_spon_7));
    InMux I__6371 (
            .O(N__34404),
            .I(N__34401));
    LocalMux I__6370 (
            .O(N__34401),
            .I(N__34398));
    Span4Mux_h I__6369 (
            .O(N__34398),
            .I(N__34394));
    InMux I__6368 (
            .O(N__34397),
            .I(N__34391));
    Odrv4 I__6367 (
            .O(N__34394),
            .I(sEEACQZ0Z_7));
    LocalMux I__6366 (
            .O(N__34391),
            .I(sEEACQZ0Z_7));
    InMux I__6365 (
            .O(N__34386),
            .I(N__34383));
    LocalMux I__6364 (
            .O(N__34383),
            .I(sEEACQ_i_7));
    CEMux I__6363 (
            .O(N__34380),
            .I(N__34377));
    LocalMux I__6362 (
            .O(N__34377),
            .I(N__34374));
    Span4Mux_h I__6361 (
            .O(N__34374),
            .I(N__34371));
    Span4Mux_h I__6360 (
            .O(N__34371),
            .I(N__34368));
    Odrv4 I__6359 (
            .O(N__34368),
            .I(sDAC_mem_31_1_sqmuxa));
    InMux I__6358 (
            .O(N__34365),
            .I(N__34361));
    InMux I__6357 (
            .O(N__34364),
            .I(N__34358));
    LocalMux I__6356 (
            .O(N__34361),
            .I(N__34355));
    LocalMux I__6355 (
            .O(N__34358),
            .I(sCounterADCZ0Z_3));
    Odrv4 I__6354 (
            .O(N__34355),
            .I(sCounterADCZ0Z_3));
    InMux I__6353 (
            .O(N__34350),
            .I(N__34346));
    InMux I__6352 (
            .O(N__34349),
            .I(N__34343));
    LocalMux I__6351 (
            .O(N__34346),
            .I(N__34338));
    LocalMux I__6350 (
            .O(N__34343),
            .I(N__34338));
    Odrv4 I__6349 (
            .O(N__34338),
            .I(sCounterADCZ0Z_2));
    InMux I__6348 (
            .O(N__34335),
            .I(N__34332));
    LocalMux I__6347 (
            .O(N__34332),
            .I(sEEADC_freqZ0Z_2));
    CascadeMux I__6346 (
            .O(N__34329),
            .I(N__34326));
    InMux I__6345 (
            .O(N__34326),
            .I(N__34323));
    LocalMux I__6344 (
            .O(N__34323),
            .I(sEEADC_freqZ0Z_3));
    InMux I__6343 (
            .O(N__34320),
            .I(N__34316));
    InMux I__6342 (
            .O(N__34319),
            .I(N__34313));
    LocalMux I__6341 (
            .O(N__34316),
            .I(N__34308));
    LocalMux I__6340 (
            .O(N__34313),
            .I(N__34308));
    Odrv12 I__6339 (
            .O(N__34308),
            .I(sCounterADCZ0Z_5));
    InMux I__6338 (
            .O(N__34305),
            .I(N__34301));
    InMux I__6337 (
            .O(N__34304),
            .I(N__34298));
    LocalMux I__6336 (
            .O(N__34301),
            .I(N__34295));
    LocalMux I__6335 (
            .O(N__34298),
            .I(sCounterADCZ0Z_4));
    Odrv4 I__6334 (
            .O(N__34295),
            .I(sCounterADCZ0Z_4));
    InMux I__6333 (
            .O(N__34290),
            .I(N__34287));
    LocalMux I__6332 (
            .O(N__34287),
            .I(sEEADC_freqZ0Z_4));
    CascadeMux I__6331 (
            .O(N__34284),
            .I(N__34281));
    InMux I__6330 (
            .O(N__34281),
            .I(N__34278));
    LocalMux I__6329 (
            .O(N__34278),
            .I(sEEADC_freqZ0Z_5));
    InMux I__6328 (
            .O(N__34275),
            .I(N__34271));
    InMux I__6327 (
            .O(N__34274),
            .I(N__34268));
    LocalMux I__6326 (
            .O(N__34271),
            .I(N__34265));
    LocalMux I__6325 (
            .O(N__34268),
            .I(sCounterADCZ0Z_6));
    Odrv4 I__6324 (
            .O(N__34265),
            .I(sCounterADCZ0Z_6));
    InMux I__6323 (
            .O(N__34260),
            .I(N__34256));
    InMux I__6322 (
            .O(N__34259),
            .I(N__34253));
    LocalMux I__6321 (
            .O(N__34256),
            .I(N__34250));
    LocalMux I__6320 (
            .O(N__34253),
            .I(sCounterADCZ0Z_7));
    Odrv12 I__6319 (
            .O(N__34250),
            .I(sCounterADCZ0Z_7));
    CascadeMux I__6318 (
            .O(N__34245),
            .I(N__34240));
    CascadeMux I__6317 (
            .O(N__34244),
            .I(N__34237));
    CascadeMux I__6316 (
            .O(N__34243),
            .I(N__34234));
    InMux I__6315 (
            .O(N__34240),
            .I(N__34231));
    InMux I__6314 (
            .O(N__34237),
            .I(N__34227));
    InMux I__6313 (
            .O(N__34234),
            .I(N__34223));
    LocalMux I__6312 (
            .O(N__34231),
            .I(N__34220));
    InMux I__6311 (
            .O(N__34230),
            .I(N__34217));
    LocalMux I__6310 (
            .O(N__34227),
            .I(N__34214));
    InMux I__6309 (
            .O(N__34226),
            .I(N__34211));
    LocalMux I__6308 (
            .O(N__34223),
            .I(N__34208));
    Span4Mux_h I__6307 (
            .O(N__34220),
            .I(N__34202));
    LocalMux I__6306 (
            .O(N__34217),
            .I(N__34202));
    Span4Mux_h I__6305 (
            .O(N__34214),
            .I(N__34197));
    LocalMux I__6304 (
            .O(N__34211),
            .I(N__34194));
    Span4Mux_v I__6303 (
            .O(N__34208),
            .I(N__34191));
    InMux I__6302 (
            .O(N__34207),
            .I(N__34188));
    Span4Mux_h I__6301 (
            .O(N__34202),
            .I(N__34185));
    InMux I__6300 (
            .O(N__34201),
            .I(N__34182));
    InMux I__6299 (
            .O(N__34200),
            .I(N__34179));
    Span4Mux_h I__6298 (
            .O(N__34197),
            .I(N__34174));
    Span4Mux_v I__6297 (
            .O(N__34194),
            .I(N__34174));
    Odrv4 I__6296 (
            .O(N__34191),
            .I(un7_spon_0));
    LocalMux I__6295 (
            .O(N__34188),
            .I(un7_spon_0));
    Odrv4 I__6294 (
            .O(N__34185),
            .I(un7_spon_0));
    LocalMux I__6293 (
            .O(N__34182),
            .I(un7_spon_0));
    LocalMux I__6292 (
            .O(N__34179),
            .I(un7_spon_0));
    Odrv4 I__6291 (
            .O(N__34174),
            .I(un7_spon_0));
    InMux I__6290 (
            .O(N__34161),
            .I(N__34158));
    LocalMux I__6289 (
            .O(N__34158),
            .I(N__34155));
    Span4Mux_v I__6288 (
            .O(N__34155),
            .I(N__34151));
    InMux I__6287 (
            .O(N__34154),
            .I(N__34148));
    Odrv4 I__6286 (
            .O(N__34151),
            .I(sEEACQZ0Z_0));
    LocalMux I__6285 (
            .O(N__34148),
            .I(sEEACQZ0Z_0));
    InMux I__6284 (
            .O(N__34143),
            .I(N__34140));
    LocalMux I__6283 (
            .O(N__34140),
            .I(sDAC_data_RNO_19Z0Z_6));
    InMux I__6282 (
            .O(N__34137),
            .I(N__34134));
    LocalMux I__6281 (
            .O(N__34134),
            .I(sDAC_mem_12Z0Z_2));
    InMux I__6280 (
            .O(N__34131),
            .I(N__34128));
    LocalMux I__6279 (
            .O(N__34128),
            .I(sDAC_mem_12Z0Z_3));
    CascadeMux I__6278 (
            .O(N__34125),
            .I(N__34122));
    InMux I__6277 (
            .O(N__34122),
            .I(N__34119));
    LocalMux I__6276 (
            .O(N__34119),
            .I(sDAC_mem_19Z0Z_1));
    InMux I__6275 (
            .O(N__34116),
            .I(N__34113));
    LocalMux I__6274 (
            .O(N__34113),
            .I(sDAC_mem_18Z0Z_1));
    InMux I__6273 (
            .O(N__34110),
            .I(N__34107));
    LocalMux I__6272 (
            .O(N__34107),
            .I(sDAC_mem_19Z0Z_2));
    InMux I__6271 (
            .O(N__34104),
            .I(N__34101));
    LocalMux I__6270 (
            .O(N__34101),
            .I(N__34098));
    Odrv12 I__6269 (
            .O(N__34098),
            .I(sDAC_data_RNO_30Z0Z_5));
    InMux I__6268 (
            .O(N__34095),
            .I(N__34092));
    LocalMux I__6267 (
            .O(N__34092),
            .I(sDAC_mem_18Z0Z_2));
    CEMux I__6266 (
            .O(N__34089),
            .I(N__34085));
    CEMux I__6265 (
            .O(N__34088),
            .I(N__34082));
    LocalMux I__6264 (
            .O(N__34085),
            .I(N__34079));
    LocalMux I__6263 (
            .O(N__34082),
            .I(sDAC_mem_18_1_sqmuxa));
    Odrv12 I__6262 (
            .O(N__34079),
            .I(sDAC_mem_18_1_sqmuxa));
    CascadeMux I__6261 (
            .O(N__34074),
            .I(sDAC_data_RNO_18Z0Z_5_cascade_));
    InMux I__6260 (
            .O(N__34071),
            .I(N__34068));
    LocalMux I__6259 (
            .O(N__34068),
            .I(sDAC_data_RNO_19Z0Z_5));
    InMux I__6258 (
            .O(N__34065),
            .I(N__34062));
    LocalMux I__6257 (
            .O(N__34062),
            .I(N__34059));
    Span4Mux_v I__6256 (
            .O(N__34059),
            .I(N__34056));
    Odrv4 I__6255 (
            .O(N__34056),
            .I(sDAC_data_2_24_ns_1_5));
    CascadeMux I__6254 (
            .O(N__34053),
            .I(sDAC_data_RNO_18Z0Z_6_cascade_));
    CascadeMux I__6253 (
            .O(N__34050),
            .I(op_le_op_le_un15_sdacdynlt4_cascade_));
    InMux I__6252 (
            .O(N__34047),
            .I(N__34044));
    LocalMux I__6251 (
            .O(N__34044),
            .I(N__34041));
    Odrv12 I__6250 (
            .O(N__34041),
            .I(un17_sdacdyn_0));
    InMux I__6249 (
            .O(N__34038),
            .I(N__34035));
    LocalMux I__6248 (
            .O(N__34035),
            .I(sDAC_mem_10Z0Z_7));
    InMux I__6247 (
            .O(N__34032),
            .I(N__34029));
    LocalMux I__6246 (
            .O(N__34029),
            .I(sDAC_mem_19Z0Z_7));
    InMux I__6245 (
            .O(N__34026),
            .I(N__34023));
    LocalMux I__6244 (
            .O(N__34023),
            .I(sDAC_mem_18Z0Z_7));
    InMux I__6243 (
            .O(N__34020),
            .I(N__34017));
    LocalMux I__6242 (
            .O(N__34017),
            .I(sDAC_mem_19Z0Z_0));
    InMux I__6241 (
            .O(N__34014),
            .I(N__34011));
    LocalMux I__6240 (
            .O(N__34011),
            .I(sDAC_mem_18Z0Z_0));
    CascadeMux I__6239 (
            .O(N__34008),
            .I(N__34005));
    InMux I__6238 (
            .O(N__34005),
            .I(N__34002));
    LocalMux I__6237 (
            .O(N__34002),
            .I(N__33999));
    Span4Mux_v I__6236 (
            .O(N__33999),
            .I(N__33996));
    Odrv4 I__6235 (
            .O(N__33996),
            .I(sDAC_mem_2Z0Z_6));
    CascadeMux I__6234 (
            .O(N__33993),
            .I(sDAC_data_2_6_bm_1_9_cascade_));
    InMux I__6233 (
            .O(N__33990),
            .I(N__33987));
    LocalMux I__6232 (
            .O(N__33987),
            .I(sDAC_mem_3Z0Z_6));
    InMux I__6231 (
            .O(N__33984),
            .I(N__33981));
    LocalMux I__6230 (
            .O(N__33981),
            .I(N__33978));
    Span4Mux_h I__6229 (
            .O(N__33978),
            .I(N__33975));
    Odrv4 I__6228 (
            .O(N__33975),
            .I(sDAC_mem_33Z0Z_1));
    CascadeMux I__6227 (
            .O(N__33972),
            .I(sDAC_data_RNO_26Z0Z_4_cascade_));
    CascadeMux I__6226 (
            .O(N__33969),
            .I(N__33965));
    CascadeMux I__6225 (
            .O(N__33968),
            .I(N__33962));
    InMux I__6224 (
            .O(N__33965),
            .I(N__33957));
    InMux I__6223 (
            .O(N__33962),
            .I(N__33957));
    LocalMux I__6222 (
            .O(N__33957),
            .I(N__33954));
    Span4Mux_v I__6221 (
            .O(N__33954),
            .I(N__33951));
    Odrv4 I__6220 (
            .O(N__33951),
            .I(sDAC_mem_1Z0Z_1));
    InMux I__6219 (
            .O(N__33948),
            .I(N__33942));
    InMux I__6218 (
            .O(N__33947),
            .I(N__33942));
    LocalMux I__6217 (
            .O(N__33942),
            .I(sDAC_mem_32Z0Z_1));
    InMux I__6216 (
            .O(N__33939),
            .I(N__33936));
    LocalMux I__6215 (
            .O(N__33936),
            .I(sDAC_data_RNO_27Z0Z_4));
    InMux I__6214 (
            .O(N__33933),
            .I(N__33930));
    LocalMux I__6213 (
            .O(N__33930),
            .I(N__33927));
    Span4Mux_v I__6212 (
            .O(N__33927),
            .I(N__33924));
    Odrv4 I__6211 (
            .O(N__33924),
            .I(sDAC_mem_33Z0Z_2));
    CascadeMux I__6210 (
            .O(N__33921),
            .I(sDAC_data_RNO_26Z0Z_5_cascade_));
    CascadeMux I__6209 (
            .O(N__33918),
            .I(N__33915));
    InMux I__6208 (
            .O(N__33915),
            .I(N__33912));
    LocalMux I__6207 (
            .O(N__33912),
            .I(N__33909));
    Odrv12 I__6206 (
            .O(N__33909),
            .I(sDAC_data_RNO_14Z0Z_5));
    CascadeMux I__6205 (
            .O(N__33906),
            .I(N__33903));
    InMux I__6204 (
            .O(N__33903),
            .I(N__33899));
    InMux I__6203 (
            .O(N__33902),
            .I(N__33896));
    LocalMux I__6202 (
            .O(N__33899),
            .I(sDAC_mem_32Z0Z_2));
    LocalMux I__6201 (
            .O(N__33896),
            .I(sDAC_mem_32Z0Z_2));
    InMux I__6200 (
            .O(N__33891),
            .I(N__33887));
    InMux I__6199 (
            .O(N__33890),
            .I(N__33884));
    LocalMux I__6198 (
            .O(N__33887),
            .I(N__33879));
    LocalMux I__6197 (
            .O(N__33884),
            .I(N__33879));
    Span4Mux_v I__6196 (
            .O(N__33879),
            .I(N__33876));
    Odrv4 I__6195 (
            .O(N__33876),
            .I(sDAC_mem_1Z0Z_2));
    InMux I__6194 (
            .O(N__33873),
            .I(N__33870));
    LocalMux I__6193 (
            .O(N__33870),
            .I(N__33867));
    Odrv4 I__6192 (
            .O(N__33867),
            .I(sDAC_data_RNO_27Z0Z_5));
    InMux I__6191 (
            .O(N__33864),
            .I(N__33861));
    LocalMux I__6190 (
            .O(N__33861),
            .I(N__33858));
    Span4Mux_v I__6189 (
            .O(N__33858),
            .I(N__33855));
    Odrv4 I__6188 (
            .O(N__33855),
            .I(sDAC_mem_33Z0Z_5));
    CascadeMux I__6187 (
            .O(N__33852),
            .I(sDAC_data_RNO_27Z0Z_8_cascade_));
    InMux I__6186 (
            .O(N__33849),
            .I(N__33843));
    InMux I__6185 (
            .O(N__33848),
            .I(N__33843));
    LocalMux I__6184 (
            .O(N__33843),
            .I(sDAC_mem_32Z0Z_5));
    InMux I__6183 (
            .O(N__33840),
            .I(N__33837));
    LocalMux I__6182 (
            .O(N__33837),
            .I(sDAC_data_RNO_26Z0Z_8));
    CascadeMux I__6181 (
            .O(N__33834),
            .I(N__33830));
    CascadeMux I__6180 (
            .O(N__33833),
            .I(N__33827));
    InMux I__6179 (
            .O(N__33830),
            .I(N__33822));
    InMux I__6178 (
            .O(N__33827),
            .I(N__33822));
    LocalMux I__6177 (
            .O(N__33822),
            .I(sDAC_mem_1Z0Z_5));
    InMux I__6176 (
            .O(N__33819),
            .I(N__33816));
    LocalMux I__6175 (
            .O(N__33816),
            .I(N__33813));
    Span4Mux_h I__6174 (
            .O(N__33813),
            .I(N__33810));
    Odrv4 I__6173 (
            .O(N__33810),
            .I(sDAC_mem_33Z0Z_6));
    CascadeMux I__6172 (
            .O(N__33807),
            .I(sDAC_data_RNO_26Z0Z_9_cascade_));
    CascadeMux I__6171 (
            .O(N__33804),
            .I(N__33800));
    CascadeMux I__6170 (
            .O(N__33803),
            .I(N__33797));
    InMux I__6169 (
            .O(N__33800),
            .I(N__33792));
    InMux I__6168 (
            .O(N__33797),
            .I(N__33792));
    LocalMux I__6167 (
            .O(N__33792),
            .I(N__33789));
    Odrv4 I__6166 (
            .O(N__33789),
            .I(sDAC_mem_32Z0Z_6));
    InMux I__6165 (
            .O(N__33786),
            .I(N__33783));
    LocalMux I__6164 (
            .O(N__33783),
            .I(sDAC_data_RNO_27Z0Z_9));
    InMux I__6163 (
            .O(N__33780),
            .I(N__33774));
    InMux I__6162 (
            .O(N__33779),
            .I(N__33774));
    LocalMux I__6161 (
            .O(N__33774),
            .I(sDAC_mem_1Z0Z_6));
    CascadeMux I__6160 (
            .O(N__33771),
            .I(sDAC_data_2_5_cascade_));
    InMux I__6159 (
            .O(N__33768),
            .I(N__33765));
    LocalMux I__6158 (
            .O(N__33765),
            .I(N__33762));
    Span4Mux_v I__6157 (
            .O(N__33762),
            .I(N__33759));
    Odrv4 I__6156 (
            .O(N__33759),
            .I(sDAC_dataZ0Z_5));
    InMux I__6155 (
            .O(N__33756),
            .I(N__33753));
    LocalMux I__6154 (
            .O(N__33753),
            .I(N__33750));
    Odrv4 I__6153 (
            .O(N__33750),
            .I(sDAC_mem_2Z0Z_2));
    CascadeMux I__6152 (
            .O(N__33747),
            .I(sDAC_data_2_6_bm_1_5_cascade_));
    InMux I__6151 (
            .O(N__33744),
            .I(N__33741));
    LocalMux I__6150 (
            .O(N__33741),
            .I(sDAC_mem_3Z0Z_2));
    InMux I__6149 (
            .O(N__33738),
            .I(N__33735));
    LocalMux I__6148 (
            .O(N__33735),
            .I(sDAC_data_RNO_15Z0Z_5));
    CascadeMux I__6147 (
            .O(N__33732),
            .I(sDAC_data_2_20_am_1_7_cascade_));
    CascadeMux I__6146 (
            .O(N__33729),
            .I(sDAC_data_RNO_17Z0Z_7_cascade_));
    CascadeMux I__6145 (
            .O(N__33726),
            .I(sDAC_data_RNO_8Z0Z_7_cascade_));
    InMux I__6144 (
            .O(N__33723),
            .I(N__33720));
    LocalMux I__6143 (
            .O(N__33720),
            .I(sDAC_data_RNO_7Z0Z_7));
    CascadeMux I__6142 (
            .O(N__33717),
            .I(sDAC_data_2_20_am_1_5_cascade_));
    CascadeMux I__6141 (
            .O(N__33714),
            .I(sDAC_data_RNO_7Z0Z_5_cascade_));
    InMux I__6140 (
            .O(N__33711),
            .I(N__33708));
    LocalMux I__6139 (
            .O(N__33708),
            .I(sDAC_data_RNO_8Z0Z_5));
    InMux I__6138 (
            .O(N__33705),
            .I(N__33702));
    LocalMux I__6137 (
            .O(N__33702),
            .I(N__33699));
    Odrv4 I__6136 (
            .O(N__33699),
            .I(sDAC_data_RNO_21Z0Z_5));
    CascadeMux I__6135 (
            .O(N__33696),
            .I(sDAC_data_RNO_10Z0Z_5_cascade_));
    InMux I__6134 (
            .O(N__33693),
            .I(N__33690));
    LocalMux I__6133 (
            .O(N__33690),
            .I(sDAC_data_2_32_ns_1_5));
    InMux I__6132 (
            .O(N__33687),
            .I(N__33684));
    LocalMux I__6131 (
            .O(N__33684),
            .I(N__33681));
    Odrv4 I__6130 (
            .O(N__33681),
            .I(sDAC_data_RNO_5Z0Z_5));
    CascadeMux I__6129 (
            .O(N__33678),
            .I(sDAC_data_2_14_ns_1_5_cascade_));
    InMux I__6128 (
            .O(N__33675),
            .I(N__33672));
    LocalMux I__6127 (
            .O(N__33672),
            .I(N__33669));
    Odrv4 I__6126 (
            .O(N__33669),
            .I(sDAC_data_RNO_4Z0Z_5));
    InMux I__6125 (
            .O(N__33666),
            .I(N__33663));
    LocalMux I__6124 (
            .O(N__33663),
            .I(sDAC_data_RNO_2Z0Z_5));
    CascadeMux I__6123 (
            .O(N__33660),
            .I(sDAC_data_RNO_1Z0Z_5_cascade_));
    InMux I__6122 (
            .O(N__33657),
            .I(N__33654));
    LocalMux I__6121 (
            .O(N__33654),
            .I(sDAC_data_2_41_ns_1_5));
    CascadeMux I__6120 (
            .O(N__33651),
            .I(sDAC_data_2_13_am_1_6_cascade_));
    InMux I__6119 (
            .O(N__33648),
            .I(N__33645));
    LocalMux I__6118 (
            .O(N__33645),
            .I(sDAC_mem_4Z0Z_3));
    InMux I__6117 (
            .O(N__33642),
            .I(N__33639));
    LocalMux I__6116 (
            .O(N__33639),
            .I(N__33636));
    Span4Mux_v I__6115 (
            .O(N__33636),
            .I(N__33633));
    Odrv4 I__6114 (
            .O(N__33633),
            .I(sDAC_mem_4Z0Z_4));
    CascadeMux I__6113 (
            .O(N__33630),
            .I(sDAC_data_2_13_am_1_7_cascade_));
    CascadeMux I__6112 (
            .O(N__33627),
            .I(N__33624));
    InMux I__6111 (
            .O(N__33624),
            .I(N__33621));
    LocalMux I__6110 (
            .O(N__33621),
            .I(sDAC_mem_2Z0Z_0));
    CascadeMux I__6109 (
            .O(N__33618),
            .I(sDAC_data_2_6_bm_1_3_cascade_));
    InMux I__6108 (
            .O(N__33615),
            .I(N__33612));
    LocalMux I__6107 (
            .O(N__33612),
            .I(sDAC_mem_3Z0Z_0));
    CascadeMux I__6106 (
            .O(N__33609),
            .I(sDAC_data_RNO_17Z0Z_5_cascade_));
    InMux I__6105 (
            .O(N__33606),
            .I(N__33603));
    LocalMux I__6104 (
            .O(N__33603),
            .I(sDAC_mem_6Z0Z_0));
    InMux I__6103 (
            .O(N__33600),
            .I(N__33597));
    LocalMux I__6102 (
            .O(N__33597),
            .I(sDAC_mem_38Z0Z_1));
    CascadeMux I__6101 (
            .O(N__33594),
            .I(sDAC_data_2_13_bm_1_4_cascade_));
    InMux I__6100 (
            .O(N__33591),
            .I(N__33588));
    LocalMux I__6099 (
            .O(N__33588),
            .I(sDAC_mem_6Z0Z_1));
    InMux I__6098 (
            .O(N__33585),
            .I(N__33582));
    LocalMux I__6097 (
            .O(N__33582),
            .I(sDAC_mem_6Z0Z_2));
    CascadeMux I__6096 (
            .O(N__33579),
            .I(sDAC_data_2_13_bm_1_5_cascade_));
    CascadeMux I__6095 (
            .O(N__33576),
            .I(sDAC_data_2_13_am_1_5_cascade_));
    InMux I__6094 (
            .O(N__33573),
            .I(N__33570));
    LocalMux I__6093 (
            .O(N__33570),
            .I(sDAC_mem_4Z0Z_2));
    InMux I__6092 (
            .O(N__33567),
            .I(N__33532));
    InMux I__6091 (
            .O(N__33566),
            .I(N__33532));
    InMux I__6090 (
            .O(N__33565),
            .I(N__33532));
    InMux I__6089 (
            .O(N__33564),
            .I(N__33532));
    InMux I__6088 (
            .O(N__33563),
            .I(N__33523));
    InMux I__6087 (
            .O(N__33562),
            .I(N__33523));
    InMux I__6086 (
            .O(N__33561),
            .I(N__33523));
    InMux I__6085 (
            .O(N__33560),
            .I(N__33523));
    InMux I__6084 (
            .O(N__33559),
            .I(N__33514));
    InMux I__6083 (
            .O(N__33558),
            .I(N__33514));
    InMux I__6082 (
            .O(N__33557),
            .I(N__33514));
    InMux I__6081 (
            .O(N__33556),
            .I(N__33514));
    InMux I__6080 (
            .O(N__33555),
            .I(N__33505));
    InMux I__6079 (
            .O(N__33554),
            .I(N__33505));
    InMux I__6078 (
            .O(N__33553),
            .I(N__33505));
    InMux I__6077 (
            .O(N__33552),
            .I(N__33505));
    InMux I__6076 (
            .O(N__33551),
            .I(N__33494));
    InMux I__6075 (
            .O(N__33550),
            .I(N__33494));
    InMux I__6074 (
            .O(N__33549),
            .I(N__33494));
    InMux I__6073 (
            .O(N__33548),
            .I(N__33494));
    InMux I__6072 (
            .O(N__33547),
            .I(N__33485));
    InMux I__6071 (
            .O(N__33546),
            .I(N__33485));
    InMux I__6070 (
            .O(N__33545),
            .I(N__33485));
    InMux I__6069 (
            .O(N__33544),
            .I(N__33485));
    InMux I__6068 (
            .O(N__33543),
            .I(N__33479));
    InMux I__6067 (
            .O(N__33542),
            .I(N__33479));
    InMux I__6066 (
            .O(N__33541),
            .I(N__33476));
    LocalMux I__6065 (
            .O(N__33532),
            .I(N__33470));
    LocalMux I__6064 (
            .O(N__33523),
            .I(N__33470));
    LocalMux I__6063 (
            .O(N__33514),
            .I(N__33465));
    LocalMux I__6062 (
            .O(N__33505),
            .I(N__33465));
    InMux I__6061 (
            .O(N__33504),
            .I(N__33460));
    InMux I__6060 (
            .O(N__33503),
            .I(N__33460));
    LocalMux I__6059 (
            .O(N__33494),
            .I(N__33453));
    LocalMux I__6058 (
            .O(N__33485),
            .I(N__33450));
    InMux I__6057 (
            .O(N__33484),
            .I(N__33447));
    LocalMux I__6056 (
            .O(N__33479),
            .I(N__33438));
    LocalMux I__6055 (
            .O(N__33476),
            .I(N__33438));
    InMux I__6054 (
            .O(N__33475),
            .I(N__33435));
    Span4Mux_h I__6053 (
            .O(N__33470),
            .I(N__33431));
    Span4Mux_h I__6052 (
            .O(N__33465),
            .I(N__33428));
    LocalMux I__6051 (
            .O(N__33460),
            .I(N__33425));
    InMux I__6050 (
            .O(N__33459),
            .I(N__33416));
    InMux I__6049 (
            .O(N__33458),
            .I(N__33416));
    InMux I__6048 (
            .O(N__33457),
            .I(N__33416));
    InMux I__6047 (
            .O(N__33456),
            .I(N__33416));
    Span4Mux_v I__6046 (
            .O(N__33453),
            .I(N__33409));
    Span4Mux_v I__6045 (
            .O(N__33450),
            .I(N__33409));
    LocalMux I__6044 (
            .O(N__33447),
            .I(N__33409));
    InMux I__6043 (
            .O(N__33446),
            .I(N__33400));
    InMux I__6042 (
            .O(N__33445),
            .I(N__33400));
    InMux I__6041 (
            .O(N__33444),
            .I(N__33400));
    InMux I__6040 (
            .O(N__33443),
            .I(N__33400));
    Span4Mux_h I__6039 (
            .O(N__33438),
            .I(N__33395));
    LocalMux I__6038 (
            .O(N__33435),
            .I(N__33395));
    InMux I__6037 (
            .O(N__33434),
            .I(N__33392));
    Span4Mux_v I__6036 (
            .O(N__33431),
            .I(N__33388));
    Span4Mux_h I__6035 (
            .O(N__33428),
            .I(N__33385));
    Span4Mux_v I__6034 (
            .O(N__33425),
            .I(N__33380));
    LocalMux I__6033 (
            .O(N__33416),
            .I(N__33380));
    Span4Mux_v I__6032 (
            .O(N__33409),
            .I(N__33375));
    LocalMux I__6031 (
            .O(N__33400),
            .I(N__33375));
    Span4Mux_v I__6030 (
            .O(N__33395),
            .I(N__33370));
    LocalMux I__6029 (
            .O(N__33392),
            .I(N__33370));
    CascadeMux I__6028 (
            .O(N__33391),
            .I(N__33367));
    Span4Mux_v I__6027 (
            .O(N__33388),
            .I(N__33364));
    Span4Mux_v I__6026 (
            .O(N__33385),
            .I(N__33361));
    Span4Mux_v I__6025 (
            .O(N__33380),
            .I(N__33356));
    Span4Mux_v I__6024 (
            .O(N__33375),
            .I(N__33356));
    Span4Mux_v I__6023 (
            .O(N__33370),
            .I(N__33353));
    InMux I__6022 (
            .O(N__33367),
            .I(N__33350));
    Span4Mux_h I__6021 (
            .O(N__33364),
            .I(N__33347));
    Span4Mux_v I__6020 (
            .O(N__33361),
            .I(N__33344));
    Span4Mux_h I__6019 (
            .O(N__33356),
            .I(N__33339));
    Span4Mux_v I__6018 (
            .O(N__33353),
            .I(N__33339));
    LocalMux I__6017 (
            .O(N__33350),
            .I(sEEPointerResetZ0));
    Odrv4 I__6016 (
            .O(N__33347),
            .I(sEEPointerResetZ0));
    Odrv4 I__6015 (
            .O(N__33344),
            .I(sEEPointerResetZ0));
    Odrv4 I__6014 (
            .O(N__33339),
            .I(sEEPointerResetZ0));
    InMux I__6013 (
            .O(N__33330),
            .I(sRAM_pointer_write_cry_17));
    InMux I__6012 (
            .O(N__33327),
            .I(N__33324));
    LocalMux I__6011 (
            .O(N__33324),
            .I(N__33321));
    Span4Mux_h I__6010 (
            .O(N__33321),
            .I(N__33317));
    InMux I__6009 (
            .O(N__33320),
            .I(N__33314));
    Span4Mux_h I__6008 (
            .O(N__33317),
            .I(N__33311));
    LocalMux I__6007 (
            .O(N__33314),
            .I(sRAM_pointer_writeZ0Z_18));
    Odrv4 I__6006 (
            .O(N__33311),
            .I(sRAM_pointer_writeZ0Z_18));
    CEMux I__6005 (
            .O(N__33306),
            .I(N__33297));
    CEMux I__6004 (
            .O(N__33305),
            .I(N__33297));
    CEMux I__6003 (
            .O(N__33304),
            .I(N__33297));
    GlobalMux I__6002 (
            .O(N__33297),
            .I(N__33294));
    gio2CtrlBuf I__6001 (
            .O(N__33294),
            .I(N_26_g));
    CascadeMux I__6000 (
            .O(N__33291),
            .I(N__33288));
    InMux I__5999 (
            .O(N__33288),
            .I(N__33278));
    InMux I__5998 (
            .O(N__33287),
            .I(N__33278));
    InMux I__5997 (
            .O(N__33286),
            .I(N__33278));
    InMux I__5996 (
            .O(N__33285),
            .I(N__33274));
    LocalMux I__5995 (
            .O(N__33278),
            .I(N__33271));
    InMux I__5994 (
            .O(N__33277),
            .I(N__33268));
    LocalMux I__5993 (
            .O(N__33274),
            .I(N__33265));
    Span4Mux_v I__5992 (
            .O(N__33271),
            .I(N__33262));
    LocalMux I__5991 (
            .O(N__33268),
            .I(N__33259));
    Span4Mux_h I__5990 (
            .O(N__33265),
            .I(N__33256));
    Span4Mux_h I__5989 (
            .O(N__33262),
            .I(N__33251));
    Span4Mux_v I__5988 (
            .O(N__33259),
            .I(N__33251));
    Sp12to4 I__5987 (
            .O(N__33256),
            .I(N__33248));
    Span4Mux_v I__5986 (
            .O(N__33251),
            .I(N__33245));
    Span12Mux_v I__5985 (
            .O(N__33248),
            .I(N__33240));
    Sp12to4 I__5984 (
            .O(N__33245),
            .I(N__33240));
    Span12Mux_h I__5983 (
            .O(N__33240),
            .I(N__33237));
    Odrv12 I__5982 (
            .O(N__33237),
            .I(spi_cs_ft_c));
    CascadeMux I__5981 (
            .O(N__33234),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_ ));
    InMux I__5980 (
            .O(N__33231),
            .I(N__33225));
    InMux I__5979 (
            .O(N__33230),
            .I(N__33225));
    LocalMux I__5978 (
            .O(N__33225),
            .I(N__33218));
    InMux I__5977 (
            .O(N__33224),
            .I(N__33215));
    InMux I__5976 (
            .O(N__33223),
            .I(N__33206));
    InMux I__5975 (
            .O(N__33222),
            .I(N__33206));
    InMux I__5974 (
            .O(N__33221),
            .I(N__33206));
    Span4Mux_v I__5973 (
            .O(N__33218),
            .I(N__33201));
    LocalMux I__5972 (
            .O(N__33215),
            .I(N__33201));
    InMux I__5971 (
            .O(N__33214),
            .I(N__33198));
    InMux I__5970 (
            .O(N__33213),
            .I(N__33195));
    LocalMux I__5969 (
            .O(N__33206),
            .I(N__33191));
    Span4Mux_v I__5968 (
            .O(N__33201),
            .I(N__33186));
    LocalMux I__5967 (
            .O(N__33198),
            .I(N__33186));
    LocalMux I__5966 (
            .O(N__33195),
            .I(N__33183));
    InMux I__5965 (
            .O(N__33194),
            .I(N__33180));
    Span4Mux_v I__5964 (
            .O(N__33191),
            .I(N__33177));
    Span4Mux_v I__5963 (
            .O(N__33186),
            .I(N__33172));
    Span4Mux_v I__5962 (
            .O(N__33183),
            .I(N__33172));
    LocalMux I__5961 (
            .O(N__33180),
            .I(N__33169));
    Odrv4 I__5960 (
            .O(N__33177),
            .I(\spi_slave_inst.spi_csZ0 ));
    Odrv4 I__5959 (
            .O(N__33172),
            .I(\spi_slave_inst.spi_csZ0 ));
    Odrv4 I__5958 (
            .O(N__33169),
            .I(\spi_slave_inst.spi_csZ0 ));
    CascadeMux I__5957 (
            .O(N__33162),
            .I(\spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_ ));
    InMux I__5956 (
            .O(N__33159),
            .I(N__33156));
    LocalMux I__5955 (
            .O(N__33156),
            .I(N__33153));
    Span4Mux_h I__5954 (
            .O(N__33153),
            .I(N__33150));
    Sp12to4 I__5953 (
            .O(N__33150),
            .I(N__33146));
    InMux I__5952 (
            .O(N__33149),
            .I(N__33143));
    Odrv12 I__5951 (
            .O(N__33146),
            .I(\spi_slave_inst.tx_done_neg_sclk_iZ0 ));
    LocalMux I__5950 (
            .O(N__33143),
            .I(\spi_slave_inst.tx_done_neg_sclk_iZ0 ));
    CascadeMux I__5949 (
            .O(N__33138),
            .I(N__33135));
    InMux I__5948 (
            .O(N__33135),
            .I(N__33132));
    LocalMux I__5947 (
            .O(N__33132),
            .I(N__33129));
    Span12Mux_v I__5946 (
            .O(N__33129),
            .I(N__33126));
    Span12Mux_h I__5945 (
            .O(N__33126),
            .I(N__33123));
    Odrv12 I__5944 (
            .O(N__33123),
            .I(spi_miso_flash_c));
    IoInMux I__5943 (
            .O(N__33120),
            .I(N__33117));
    LocalMux I__5942 (
            .O(N__33117),
            .I(N__33114));
    IoSpan4Mux I__5941 (
            .O(N__33114),
            .I(N__33111));
    Span4Mux_s2_h I__5940 (
            .O(N__33111),
            .I(N__33108));
    Sp12to4 I__5939 (
            .O(N__33108),
            .I(N__33105));
    Span12Mux_s8_h I__5938 (
            .O(N__33105),
            .I(N__33102));
    Odrv12 I__5937 (
            .O(N__33102),
            .I(spi_miso_rpi_c));
    CascadeMux I__5936 (
            .O(N__33099),
            .I(sDAC_data_2_13_bm_1_3_cascade_));
    InMux I__5935 (
            .O(N__33096),
            .I(N__33093));
    LocalMux I__5934 (
            .O(N__33093),
            .I(N__33089));
    InMux I__5933 (
            .O(N__33092),
            .I(N__33086));
    Odrv4 I__5932 (
            .O(N__33089),
            .I(sRAM_pointer_writeZ0Z_10));
    LocalMux I__5931 (
            .O(N__33086),
            .I(sRAM_pointer_writeZ0Z_10));
    InMux I__5930 (
            .O(N__33081),
            .I(sRAM_pointer_write_cry_9));
    CascadeMux I__5929 (
            .O(N__33078),
            .I(N__33075));
    InMux I__5928 (
            .O(N__33075),
            .I(N__33072));
    LocalMux I__5927 (
            .O(N__33072),
            .I(N__33068));
    InMux I__5926 (
            .O(N__33071),
            .I(N__33065));
    Odrv4 I__5925 (
            .O(N__33068),
            .I(sRAM_pointer_writeZ0Z_11));
    LocalMux I__5924 (
            .O(N__33065),
            .I(sRAM_pointer_writeZ0Z_11));
    InMux I__5923 (
            .O(N__33060),
            .I(sRAM_pointer_write_cry_10));
    InMux I__5922 (
            .O(N__33057),
            .I(N__33054));
    LocalMux I__5921 (
            .O(N__33054),
            .I(N__33051));
    Span4Mux_h I__5920 (
            .O(N__33051),
            .I(N__33047));
    InMux I__5919 (
            .O(N__33050),
            .I(N__33044));
    Odrv4 I__5918 (
            .O(N__33047),
            .I(sRAM_pointer_writeZ0Z_12));
    LocalMux I__5917 (
            .O(N__33044),
            .I(sRAM_pointer_writeZ0Z_12));
    InMux I__5916 (
            .O(N__33039),
            .I(sRAM_pointer_write_cry_11));
    CascadeMux I__5915 (
            .O(N__33036),
            .I(N__33033));
    InMux I__5914 (
            .O(N__33033),
            .I(N__33030));
    LocalMux I__5913 (
            .O(N__33030),
            .I(N__33026));
    InMux I__5912 (
            .O(N__33029),
            .I(N__33023));
    Odrv4 I__5911 (
            .O(N__33026),
            .I(sRAM_pointer_writeZ0Z_13));
    LocalMux I__5910 (
            .O(N__33023),
            .I(sRAM_pointer_writeZ0Z_13));
    InMux I__5909 (
            .O(N__33018),
            .I(sRAM_pointer_write_cry_12));
    InMux I__5908 (
            .O(N__33015),
            .I(N__33012));
    LocalMux I__5907 (
            .O(N__33012),
            .I(N__33009));
    Span4Mux_h I__5906 (
            .O(N__33009),
            .I(N__33005));
    InMux I__5905 (
            .O(N__33008),
            .I(N__33002));
    Odrv4 I__5904 (
            .O(N__33005),
            .I(sRAM_pointer_writeZ0Z_14));
    LocalMux I__5903 (
            .O(N__33002),
            .I(sRAM_pointer_writeZ0Z_14));
    InMux I__5902 (
            .O(N__32997),
            .I(sRAM_pointer_write_cry_13));
    InMux I__5901 (
            .O(N__32994),
            .I(N__32991));
    LocalMux I__5900 (
            .O(N__32991),
            .I(N__32988));
    Span4Mux_h I__5899 (
            .O(N__32988),
            .I(N__32984));
    InMux I__5898 (
            .O(N__32987),
            .I(N__32981));
    Odrv4 I__5897 (
            .O(N__32984),
            .I(sRAM_pointer_writeZ0Z_15));
    LocalMux I__5896 (
            .O(N__32981),
            .I(sRAM_pointer_writeZ0Z_15));
    InMux I__5895 (
            .O(N__32976),
            .I(sRAM_pointer_write_cry_14));
    InMux I__5894 (
            .O(N__32973),
            .I(N__32970));
    LocalMux I__5893 (
            .O(N__32970),
            .I(N__32966));
    InMux I__5892 (
            .O(N__32969),
            .I(N__32963));
    Span4Mux_v I__5891 (
            .O(N__32966),
            .I(N__32960));
    LocalMux I__5890 (
            .O(N__32963),
            .I(sRAM_pointer_writeZ0Z_16));
    Odrv4 I__5889 (
            .O(N__32960),
            .I(sRAM_pointer_writeZ0Z_16));
    InMux I__5888 (
            .O(N__32955),
            .I(bfn_13_20_0_));
    InMux I__5887 (
            .O(N__32952),
            .I(N__32949));
    LocalMux I__5886 (
            .O(N__32949),
            .I(N__32946));
    Span4Mux_h I__5885 (
            .O(N__32946),
            .I(N__32943));
    Span4Mux_h I__5884 (
            .O(N__32943),
            .I(N__32939));
    InMux I__5883 (
            .O(N__32942),
            .I(N__32936));
    Odrv4 I__5882 (
            .O(N__32939),
            .I(sRAM_pointer_writeZ0Z_17));
    LocalMux I__5881 (
            .O(N__32936),
            .I(sRAM_pointer_writeZ0Z_17));
    InMux I__5880 (
            .O(N__32931),
            .I(sRAM_pointer_write_cry_16));
    InMux I__5879 (
            .O(N__32928),
            .I(sRAM_pointer_write_cry_0));
    InMux I__5878 (
            .O(N__32925),
            .I(N__32922));
    LocalMux I__5877 (
            .O(N__32922),
            .I(N__32919));
    Span4Mux_h I__5876 (
            .O(N__32919),
            .I(N__32915));
    InMux I__5875 (
            .O(N__32918),
            .I(N__32912));
    Odrv4 I__5874 (
            .O(N__32915),
            .I(sRAM_pointer_writeZ0Z_2));
    LocalMux I__5873 (
            .O(N__32912),
            .I(sRAM_pointer_writeZ0Z_2));
    InMux I__5872 (
            .O(N__32907),
            .I(sRAM_pointer_write_cry_1));
    InMux I__5871 (
            .O(N__32904),
            .I(N__32901));
    LocalMux I__5870 (
            .O(N__32901),
            .I(N__32898));
    Span4Mux_h I__5869 (
            .O(N__32898),
            .I(N__32894));
    InMux I__5868 (
            .O(N__32897),
            .I(N__32891));
    Odrv4 I__5867 (
            .O(N__32894),
            .I(sRAM_pointer_writeZ0Z_3));
    LocalMux I__5866 (
            .O(N__32891),
            .I(sRAM_pointer_writeZ0Z_3));
    InMux I__5865 (
            .O(N__32886),
            .I(sRAM_pointer_write_cry_2));
    InMux I__5864 (
            .O(N__32883),
            .I(N__32880));
    LocalMux I__5863 (
            .O(N__32880),
            .I(N__32877));
    Span4Mux_h I__5862 (
            .O(N__32877),
            .I(N__32874));
    Span4Mux_h I__5861 (
            .O(N__32874),
            .I(N__32870));
    InMux I__5860 (
            .O(N__32873),
            .I(N__32867));
    Odrv4 I__5859 (
            .O(N__32870),
            .I(sRAM_pointer_writeZ0Z_4));
    LocalMux I__5858 (
            .O(N__32867),
            .I(sRAM_pointer_writeZ0Z_4));
    InMux I__5857 (
            .O(N__32862),
            .I(sRAM_pointer_write_cry_3));
    CascadeMux I__5856 (
            .O(N__32859),
            .I(N__32856));
    InMux I__5855 (
            .O(N__32856),
            .I(N__32853));
    LocalMux I__5854 (
            .O(N__32853),
            .I(N__32849));
    InMux I__5853 (
            .O(N__32852),
            .I(N__32846));
    Odrv4 I__5852 (
            .O(N__32849),
            .I(sRAM_pointer_writeZ0Z_5));
    LocalMux I__5851 (
            .O(N__32846),
            .I(sRAM_pointer_writeZ0Z_5));
    InMux I__5850 (
            .O(N__32841),
            .I(sRAM_pointer_write_cry_4));
    InMux I__5849 (
            .O(N__32838),
            .I(N__32835));
    LocalMux I__5848 (
            .O(N__32835),
            .I(N__32831));
    InMux I__5847 (
            .O(N__32834),
            .I(N__32828));
    Odrv4 I__5846 (
            .O(N__32831),
            .I(sRAM_pointer_writeZ0Z_6));
    LocalMux I__5845 (
            .O(N__32828),
            .I(sRAM_pointer_writeZ0Z_6));
    InMux I__5844 (
            .O(N__32823),
            .I(sRAM_pointer_write_cry_5));
    InMux I__5843 (
            .O(N__32820),
            .I(N__32817));
    LocalMux I__5842 (
            .O(N__32817),
            .I(N__32813));
    InMux I__5841 (
            .O(N__32816),
            .I(N__32810));
    Odrv4 I__5840 (
            .O(N__32813),
            .I(sRAM_pointer_writeZ0Z_7));
    LocalMux I__5839 (
            .O(N__32810),
            .I(sRAM_pointer_writeZ0Z_7));
    InMux I__5838 (
            .O(N__32805),
            .I(sRAM_pointer_write_cry_6));
    InMux I__5837 (
            .O(N__32802),
            .I(N__32799));
    LocalMux I__5836 (
            .O(N__32799),
            .I(N__32796));
    Span4Mux_v I__5835 (
            .O(N__32796),
            .I(N__32792));
    InMux I__5834 (
            .O(N__32795),
            .I(N__32789));
    Odrv4 I__5833 (
            .O(N__32792),
            .I(sRAM_pointer_writeZ0Z_8));
    LocalMux I__5832 (
            .O(N__32789),
            .I(sRAM_pointer_writeZ0Z_8));
    InMux I__5831 (
            .O(N__32784),
            .I(bfn_13_19_0_));
    InMux I__5830 (
            .O(N__32781),
            .I(N__32778));
    LocalMux I__5829 (
            .O(N__32778),
            .I(N__32775));
    Span4Mux_v I__5828 (
            .O(N__32775),
            .I(N__32772));
    Span4Mux_h I__5827 (
            .O(N__32772),
            .I(N__32768));
    InMux I__5826 (
            .O(N__32771),
            .I(N__32765));
    Odrv4 I__5825 (
            .O(N__32768),
            .I(sRAM_pointer_writeZ0Z_9));
    LocalMux I__5824 (
            .O(N__32765),
            .I(sRAM_pointer_writeZ0Z_9));
    InMux I__5823 (
            .O(N__32760),
            .I(sRAM_pointer_write_cry_8));
    CascadeMux I__5822 (
            .O(N__32757),
            .I(N_107_cascade_));
    IoInMux I__5821 (
            .O(N__32754),
            .I(N__32751));
    LocalMux I__5820 (
            .O(N__32751),
            .I(N__32748));
    IoSpan4Mux I__5819 (
            .O(N__32748),
            .I(N__32745));
    Span4Mux_s3_h I__5818 (
            .O(N__32745),
            .I(N__32742));
    Sp12to4 I__5817 (
            .O(N__32742),
            .I(N__32739));
    Span12Mux_v I__5816 (
            .O(N__32739),
            .I(N__32736));
    Span12Mux_h I__5815 (
            .O(N__32736),
            .I(N__32732));
    InMux I__5814 (
            .O(N__32735),
            .I(N__32729));
    Odrv12 I__5813 (
            .O(N__32732),
            .I(RAM_DATA_cl_5Z0Z_15));
    LocalMux I__5812 (
            .O(N__32729),
            .I(RAM_DATA_cl_5Z0Z_15));
    CascadeMux I__5811 (
            .O(N__32724),
            .I(N_108_cascade_));
    IoInMux I__5810 (
            .O(N__32721),
            .I(N__32718));
    LocalMux I__5809 (
            .O(N__32718),
            .I(N__32715));
    IoSpan4Mux I__5808 (
            .O(N__32715),
            .I(N__32712));
    IoSpan4Mux I__5807 (
            .O(N__32712),
            .I(N__32709));
    Span4Mux_s3_h I__5806 (
            .O(N__32709),
            .I(N__32706));
    Span4Mux_h I__5805 (
            .O(N__32706),
            .I(N__32703));
    Span4Mux_h I__5804 (
            .O(N__32703),
            .I(N__32699));
    InMux I__5803 (
            .O(N__32702),
            .I(N__32696));
    Odrv4 I__5802 (
            .O(N__32699),
            .I(RAM_DATA_cl_6Z0Z_15));
    LocalMux I__5801 (
            .O(N__32696),
            .I(RAM_DATA_cl_6Z0Z_15));
    InMux I__5800 (
            .O(N__32691),
            .I(N__32672));
    InMux I__5799 (
            .O(N__32690),
            .I(N__32665));
    InMux I__5798 (
            .O(N__32689),
            .I(N__32665));
    InMux I__5797 (
            .O(N__32688),
            .I(N__32665));
    InMux I__5796 (
            .O(N__32687),
            .I(N__32658));
    InMux I__5795 (
            .O(N__32686),
            .I(N__32658));
    InMux I__5794 (
            .O(N__32685),
            .I(N__32658));
    InMux I__5793 (
            .O(N__32684),
            .I(N__32649));
    InMux I__5792 (
            .O(N__32683),
            .I(N__32649));
    InMux I__5791 (
            .O(N__32682),
            .I(N__32649));
    InMux I__5790 (
            .O(N__32681),
            .I(N__32649));
    InMux I__5789 (
            .O(N__32680),
            .I(N__32640));
    InMux I__5788 (
            .O(N__32679),
            .I(N__32640));
    InMux I__5787 (
            .O(N__32678),
            .I(N__32640));
    InMux I__5786 (
            .O(N__32677),
            .I(N__32640));
    CascadeMux I__5785 (
            .O(N__32676),
            .I(N__32637));
    CascadeMux I__5784 (
            .O(N__32675),
            .I(N__32628));
    LocalMux I__5783 (
            .O(N__32672),
            .I(N__32625));
    LocalMux I__5782 (
            .O(N__32665),
            .I(N__32614));
    LocalMux I__5781 (
            .O(N__32658),
            .I(N__32614));
    LocalMux I__5780 (
            .O(N__32649),
            .I(N__32614));
    LocalMux I__5779 (
            .O(N__32640),
            .I(N__32614));
    InMux I__5778 (
            .O(N__32637),
            .I(N__32611));
    InMux I__5777 (
            .O(N__32636),
            .I(N__32604));
    InMux I__5776 (
            .O(N__32635),
            .I(N__32604));
    InMux I__5775 (
            .O(N__32634),
            .I(N__32604));
    InMux I__5774 (
            .O(N__32633),
            .I(N__32599));
    InMux I__5773 (
            .O(N__32632),
            .I(N__32599));
    InMux I__5772 (
            .O(N__32631),
            .I(N__32596));
    InMux I__5771 (
            .O(N__32628),
            .I(N__32591));
    Span4Mux_v I__5770 (
            .O(N__32625),
            .I(N__32587));
    InMux I__5769 (
            .O(N__32624),
            .I(N__32584));
    CascadeMux I__5768 (
            .O(N__32623),
            .I(N__32580));
    Span4Mux_v I__5767 (
            .O(N__32614),
            .I(N__32569));
    LocalMux I__5766 (
            .O(N__32611),
            .I(N__32569));
    LocalMux I__5765 (
            .O(N__32604),
            .I(N__32569));
    LocalMux I__5764 (
            .O(N__32599),
            .I(N__32569));
    LocalMux I__5763 (
            .O(N__32596),
            .I(N__32569));
    InMux I__5762 (
            .O(N__32595),
            .I(N__32566));
    CascadeMux I__5761 (
            .O(N__32594),
            .I(N__32563));
    LocalMux I__5760 (
            .O(N__32591),
            .I(N__32559));
    CascadeMux I__5759 (
            .O(N__32590),
            .I(N__32555));
    Span4Mux_h I__5758 (
            .O(N__32587),
            .I(N__32551));
    LocalMux I__5757 (
            .O(N__32584),
            .I(N__32548));
    IoInMux I__5756 (
            .O(N__32583),
            .I(N__32543));
    InMux I__5755 (
            .O(N__32580),
            .I(N__32540));
    Span4Mux_v I__5754 (
            .O(N__32569),
            .I(N__32535));
    LocalMux I__5753 (
            .O(N__32566),
            .I(N__32535));
    InMux I__5752 (
            .O(N__32563),
            .I(N__32532));
    InMux I__5751 (
            .O(N__32562),
            .I(N__32529));
    Span4Mux_v I__5750 (
            .O(N__32559),
            .I(N__32526));
    InMux I__5749 (
            .O(N__32558),
            .I(N__32523));
    InMux I__5748 (
            .O(N__32555),
            .I(N__32520));
    CascadeMux I__5747 (
            .O(N__32554),
            .I(N__32517));
    Span4Mux_h I__5746 (
            .O(N__32551),
            .I(N__32510));
    Span4Mux_v I__5745 (
            .O(N__32548),
            .I(N__32510));
    InMux I__5744 (
            .O(N__32547),
            .I(N__32507));
    CascadeMux I__5743 (
            .O(N__32546),
            .I(N__32490));
    LocalMux I__5742 (
            .O(N__32543),
            .I(N__32487));
    LocalMux I__5741 (
            .O(N__32540),
            .I(N__32484));
    Span4Mux_v I__5740 (
            .O(N__32535),
            .I(N__32479));
    LocalMux I__5739 (
            .O(N__32532),
            .I(N__32479));
    LocalMux I__5738 (
            .O(N__32529),
            .I(N__32476));
    Span4Mux_v I__5737 (
            .O(N__32526),
            .I(N__32471));
    LocalMux I__5736 (
            .O(N__32523),
            .I(N__32471));
    LocalMux I__5735 (
            .O(N__32520),
            .I(N__32463));
    InMux I__5734 (
            .O(N__32517),
            .I(N__32456));
    InMux I__5733 (
            .O(N__32516),
            .I(N__32456));
    CEMux I__5732 (
            .O(N__32515),
            .I(N__32456));
    Span4Mux_v I__5731 (
            .O(N__32510),
            .I(N__32451));
    LocalMux I__5730 (
            .O(N__32507),
            .I(N__32451));
    CascadeMux I__5729 (
            .O(N__32506),
            .I(N__32448));
    CascadeMux I__5728 (
            .O(N__32505),
            .I(N__32445));
    CascadeMux I__5727 (
            .O(N__32504),
            .I(N__32441));
    InMux I__5726 (
            .O(N__32503),
            .I(N__32434));
    InMux I__5725 (
            .O(N__32502),
            .I(N__32434));
    InMux I__5724 (
            .O(N__32501),
            .I(N__32434));
    InMux I__5723 (
            .O(N__32500),
            .I(N__32423));
    InMux I__5722 (
            .O(N__32499),
            .I(N__32423));
    InMux I__5721 (
            .O(N__32498),
            .I(N__32423));
    InMux I__5720 (
            .O(N__32497),
            .I(N__32423));
    InMux I__5719 (
            .O(N__32496),
            .I(N__32423));
    InMux I__5718 (
            .O(N__32495),
            .I(N__32414));
    InMux I__5717 (
            .O(N__32494),
            .I(N__32414));
    InMux I__5716 (
            .O(N__32493),
            .I(N__32414));
    InMux I__5715 (
            .O(N__32490),
            .I(N__32414));
    Span4Mux_s2_h I__5714 (
            .O(N__32487),
            .I(N__32410));
    Span4Mux_v I__5713 (
            .O(N__32484),
            .I(N__32407));
    Span4Mux_v I__5712 (
            .O(N__32479),
            .I(N__32404));
    Span4Mux_h I__5711 (
            .O(N__32476),
            .I(N__32399));
    Span4Mux_v I__5710 (
            .O(N__32471),
            .I(N__32399));
    InMux I__5709 (
            .O(N__32470),
            .I(N__32391));
    InMux I__5708 (
            .O(N__32469),
            .I(N__32391));
    InMux I__5707 (
            .O(N__32468),
            .I(N__32391));
    InMux I__5706 (
            .O(N__32467),
            .I(N__32386));
    InMux I__5705 (
            .O(N__32466),
            .I(N__32386));
    Span4Mux_v I__5704 (
            .O(N__32463),
            .I(N__32383));
    LocalMux I__5703 (
            .O(N__32456),
            .I(N__32380));
    Span4Mux_v I__5702 (
            .O(N__32451),
            .I(N__32377));
    InMux I__5701 (
            .O(N__32448),
            .I(N__32372));
    InMux I__5700 (
            .O(N__32445),
            .I(N__32372));
    InMux I__5699 (
            .O(N__32444),
            .I(N__32367));
    InMux I__5698 (
            .O(N__32441),
            .I(N__32367));
    LocalMux I__5697 (
            .O(N__32434),
            .I(N__32364));
    LocalMux I__5696 (
            .O(N__32423),
            .I(N__32361));
    LocalMux I__5695 (
            .O(N__32414),
            .I(N__32358));
    InMux I__5694 (
            .O(N__32413),
            .I(N__32355));
    Sp12to4 I__5693 (
            .O(N__32410),
            .I(N__32347));
    Span4Mux_h I__5692 (
            .O(N__32407),
            .I(N__32340));
    Span4Mux_h I__5691 (
            .O(N__32404),
            .I(N__32340));
    Span4Mux_v I__5690 (
            .O(N__32399),
            .I(N__32340));
    InMux I__5689 (
            .O(N__32398),
            .I(N__32337));
    LocalMux I__5688 (
            .O(N__32391),
            .I(N__32332));
    LocalMux I__5687 (
            .O(N__32386),
            .I(N__32332));
    Span4Mux_h I__5686 (
            .O(N__32383),
            .I(N__32327));
    Span4Mux_h I__5685 (
            .O(N__32380),
            .I(N__32327));
    Span4Mux_v I__5684 (
            .O(N__32377),
            .I(N__32323));
    LocalMux I__5683 (
            .O(N__32372),
            .I(N__32318));
    LocalMux I__5682 (
            .O(N__32367),
            .I(N__32318));
    Span4Mux_v I__5681 (
            .O(N__32364),
            .I(N__32309));
    Span4Mux_h I__5680 (
            .O(N__32361),
            .I(N__32309));
    Span4Mux_h I__5679 (
            .O(N__32358),
            .I(N__32309));
    LocalMux I__5678 (
            .O(N__32355),
            .I(N__32309));
    InMux I__5677 (
            .O(N__32354),
            .I(N__32302));
    InMux I__5676 (
            .O(N__32353),
            .I(N__32302));
    InMux I__5675 (
            .O(N__32352),
            .I(N__32302));
    InMux I__5674 (
            .O(N__32351),
            .I(N__32299));
    InMux I__5673 (
            .O(N__32350),
            .I(N__32296));
    Span12Mux_v I__5672 (
            .O(N__32347),
            .I(N__32293));
    Span4Mux_v I__5671 (
            .O(N__32340),
            .I(N__32290));
    LocalMux I__5670 (
            .O(N__32337),
            .I(N__32287));
    Span4Mux_v I__5669 (
            .O(N__32332),
            .I(N__32282));
    Span4Mux_v I__5668 (
            .O(N__32327),
            .I(N__32282));
    IoInMux I__5667 (
            .O(N__32326),
            .I(N__32279));
    Sp12to4 I__5666 (
            .O(N__32323),
            .I(N__32276));
    Span12Mux_s9_v I__5665 (
            .O(N__32318),
            .I(N__32265));
    Sp12to4 I__5664 (
            .O(N__32309),
            .I(N__32265));
    LocalMux I__5663 (
            .O(N__32302),
            .I(N__32265));
    LocalMux I__5662 (
            .O(N__32299),
            .I(N__32265));
    LocalMux I__5661 (
            .O(N__32296),
            .I(N__32265));
    Span12Mux_v I__5660 (
            .O(N__32293),
            .I(N__32262));
    Sp12to4 I__5659 (
            .O(N__32290),
            .I(N__32259));
    Sp12to4 I__5658 (
            .O(N__32287),
            .I(N__32254));
    Sp12to4 I__5657 (
            .O(N__32282),
            .I(N__32254));
    LocalMux I__5656 (
            .O(N__32279),
            .I(N__32251));
    Span12Mux_h I__5655 (
            .O(N__32276),
            .I(N__32246));
    Span12Mux_v I__5654 (
            .O(N__32265),
            .I(N__32246));
    Span12Mux_h I__5653 (
            .O(N__32262),
            .I(N__32239));
    Span12Mux_h I__5652 (
            .O(N__32259),
            .I(N__32239));
    Span12Mux_v I__5651 (
            .O(N__32254),
            .I(N__32239));
    IoSpan4Mux I__5650 (
            .O(N__32251),
            .I(N__32236));
    Odrv12 I__5649 (
            .O(N__32246),
            .I(LED3_c));
    Odrv12 I__5648 (
            .O(N__32239),
            .I(LED3_c));
    Odrv4 I__5647 (
            .O(N__32236),
            .I(LED3_c));
    CascadeMux I__5646 (
            .O(N__32229),
            .I(N__32208));
    CascadeMux I__5645 (
            .O(N__32228),
            .I(N__32205));
    CascadeMux I__5644 (
            .O(N__32227),
            .I(N__32202));
    CascadeMux I__5643 (
            .O(N__32226),
            .I(N__32199));
    InMux I__5642 (
            .O(N__32225),
            .I(N__32187));
    InMux I__5641 (
            .O(N__32224),
            .I(N__32187));
    InMux I__5640 (
            .O(N__32223),
            .I(N__32187));
    InMux I__5639 (
            .O(N__32222),
            .I(N__32187));
    CascadeMux I__5638 (
            .O(N__32221),
            .I(N__32172));
    CascadeMux I__5637 (
            .O(N__32220),
            .I(N__32169));
    CascadeMux I__5636 (
            .O(N__32219),
            .I(N__32166));
    CascadeMux I__5635 (
            .O(N__32218),
            .I(N__32160));
    InMux I__5634 (
            .O(N__32217),
            .I(N__32154));
    InMux I__5633 (
            .O(N__32216),
            .I(N__32154));
    InMux I__5632 (
            .O(N__32215),
            .I(N__32148));
    InMux I__5631 (
            .O(N__32214),
            .I(N__32141));
    InMux I__5630 (
            .O(N__32213),
            .I(N__32141));
    InMux I__5629 (
            .O(N__32212),
            .I(N__32141));
    InMux I__5628 (
            .O(N__32211),
            .I(N__32138));
    InMux I__5627 (
            .O(N__32208),
            .I(N__32123));
    InMux I__5626 (
            .O(N__32205),
            .I(N__32123));
    InMux I__5625 (
            .O(N__32202),
            .I(N__32123));
    InMux I__5624 (
            .O(N__32199),
            .I(N__32123));
    InMux I__5623 (
            .O(N__32198),
            .I(N__32123));
    InMux I__5622 (
            .O(N__32197),
            .I(N__32123));
    InMux I__5621 (
            .O(N__32196),
            .I(N__32123));
    LocalMux I__5620 (
            .O(N__32187),
            .I(N__32120));
    InMux I__5619 (
            .O(N__32186),
            .I(N__32103));
    InMux I__5618 (
            .O(N__32185),
            .I(N__32103));
    InMux I__5617 (
            .O(N__32184),
            .I(N__32103));
    InMux I__5616 (
            .O(N__32183),
            .I(N__32103));
    InMux I__5615 (
            .O(N__32182),
            .I(N__32103));
    InMux I__5614 (
            .O(N__32181),
            .I(N__32103));
    InMux I__5613 (
            .O(N__32180),
            .I(N__32103));
    InMux I__5612 (
            .O(N__32179),
            .I(N__32103));
    CascadeMux I__5611 (
            .O(N__32178),
            .I(N__32099));
    InMux I__5610 (
            .O(N__32177),
            .I(N__32094));
    InMux I__5609 (
            .O(N__32176),
            .I(N__32094));
    InMux I__5608 (
            .O(N__32175),
            .I(N__32091));
    InMux I__5607 (
            .O(N__32172),
            .I(N__32088));
    InMux I__5606 (
            .O(N__32169),
            .I(N__32077));
    InMux I__5605 (
            .O(N__32166),
            .I(N__32077));
    InMux I__5604 (
            .O(N__32165),
            .I(N__32077));
    InMux I__5603 (
            .O(N__32164),
            .I(N__32077));
    InMux I__5602 (
            .O(N__32163),
            .I(N__32077));
    InMux I__5601 (
            .O(N__32160),
            .I(N__32072));
    InMux I__5600 (
            .O(N__32159),
            .I(N__32072));
    LocalMux I__5599 (
            .O(N__32154),
            .I(N__32069));
    InMux I__5598 (
            .O(N__32153),
            .I(N__32063));
    InMux I__5597 (
            .O(N__32152),
            .I(N__32058));
    InMux I__5596 (
            .O(N__32151),
            .I(N__32058));
    LocalMux I__5595 (
            .O(N__32148),
            .I(N__32055));
    LocalMux I__5594 (
            .O(N__32141),
            .I(N__32052));
    LocalMux I__5593 (
            .O(N__32138),
            .I(N__32049));
    LocalMux I__5592 (
            .O(N__32123),
            .I(N__32042));
    Span4Mux_h I__5591 (
            .O(N__32120),
            .I(N__32042));
    LocalMux I__5590 (
            .O(N__32103),
            .I(N__32042));
    InMux I__5589 (
            .O(N__32102),
            .I(N__32037));
    InMux I__5588 (
            .O(N__32099),
            .I(N__32037));
    LocalMux I__5587 (
            .O(N__32094),
            .I(N__32032));
    LocalMux I__5586 (
            .O(N__32091),
            .I(N__32032));
    LocalMux I__5585 (
            .O(N__32088),
            .I(N__32023));
    LocalMux I__5584 (
            .O(N__32077),
            .I(N__32023));
    LocalMux I__5583 (
            .O(N__32072),
            .I(N__32023));
    Span4Mux_v I__5582 (
            .O(N__32069),
            .I(N__32023));
    InMux I__5581 (
            .O(N__32068),
            .I(N__32016));
    InMux I__5580 (
            .O(N__32067),
            .I(N__32016));
    InMux I__5579 (
            .O(N__32066),
            .I(N__32016));
    LocalMux I__5578 (
            .O(N__32063),
            .I(N__32009));
    LocalMux I__5577 (
            .O(N__32058),
            .I(N__32009));
    Span12Mux_v I__5576 (
            .O(N__32055),
            .I(N__32009));
    Span4Mux_h I__5575 (
            .O(N__32052),
            .I(N__32004));
    Span4Mux_h I__5574 (
            .O(N__32049),
            .I(N__32004));
    Span4Mux_h I__5573 (
            .O(N__32042),
            .I(N__32001));
    LocalMux I__5572 (
            .O(N__32037),
            .I(N__31998));
    Span4Mux_v I__5571 (
            .O(N__32032),
            .I(N__31993));
    Span4Mux_v I__5570 (
            .O(N__32023),
            .I(N__31993));
    LocalMux I__5569 (
            .O(N__32016),
            .I(un4_sacqtime_cry_23_THRU_CO));
    Odrv12 I__5568 (
            .O(N__32009),
            .I(un4_sacqtime_cry_23_THRU_CO));
    Odrv4 I__5567 (
            .O(N__32004),
            .I(un4_sacqtime_cry_23_THRU_CO));
    Odrv4 I__5566 (
            .O(N__32001),
            .I(un4_sacqtime_cry_23_THRU_CO));
    Odrv4 I__5565 (
            .O(N__31998),
            .I(un4_sacqtime_cry_23_THRU_CO));
    Odrv4 I__5564 (
            .O(N__31993),
            .I(un4_sacqtime_cry_23_THRU_CO));
    CascadeMux I__5563 (
            .O(N__31980),
            .I(N_95_cascade_));
    InMux I__5562 (
            .O(N__31977),
            .I(N__31974));
    LocalMux I__5561 (
            .O(N__31974),
            .I(N__31970));
    InMux I__5560 (
            .O(N__31973),
            .I(N__31952));
    Span4Mux_h I__5559 (
            .O(N__31970),
            .I(N__31949));
    InMux I__5558 (
            .O(N__31969),
            .I(N__31927));
    InMux I__5557 (
            .O(N__31968),
            .I(N__31927));
    InMux I__5556 (
            .O(N__31967),
            .I(N__31927));
    InMux I__5555 (
            .O(N__31966),
            .I(N__31922));
    InMux I__5554 (
            .O(N__31965),
            .I(N__31922));
    InMux I__5553 (
            .O(N__31964),
            .I(N__31917));
    InMux I__5552 (
            .O(N__31963),
            .I(N__31917));
    InMux I__5551 (
            .O(N__31962),
            .I(N__31897));
    InMux I__5550 (
            .O(N__31961),
            .I(N__31897));
    InMux I__5549 (
            .O(N__31960),
            .I(N__31897));
    InMux I__5548 (
            .O(N__31959),
            .I(N__31897));
    InMux I__5547 (
            .O(N__31958),
            .I(N__31897));
    InMux I__5546 (
            .O(N__31957),
            .I(N__31897));
    InMux I__5545 (
            .O(N__31956),
            .I(N__31892));
    InMux I__5544 (
            .O(N__31955),
            .I(N__31892));
    LocalMux I__5543 (
            .O(N__31952),
            .I(N__31889));
    Span4Mux_v I__5542 (
            .O(N__31949),
            .I(N__31886));
    InMux I__5541 (
            .O(N__31948),
            .I(N__31873));
    InMux I__5540 (
            .O(N__31947),
            .I(N__31873));
    InMux I__5539 (
            .O(N__31946),
            .I(N__31873));
    InMux I__5538 (
            .O(N__31945),
            .I(N__31873));
    InMux I__5537 (
            .O(N__31944),
            .I(N__31866));
    InMux I__5536 (
            .O(N__31943),
            .I(N__31866));
    InMux I__5535 (
            .O(N__31942),
            .I(N__31866));
    InMux I__5534 (
            .O(N__31941),
            .I(N__31849));
    InMux I__5533 (
            .O(N__31940),
            .I(N__31849));
    InMux I__5532 (
            .O(N__31939),
            .I(N__31849));
    InMux I__5531 (
            .O(N__31938),
            .I(N__31849));
    InMux I__5530 (
            .O(N__31937),
            .I(N__31849));
    InMux I__5529 (
            .O(N__31936),
            .I(N__31849));
    InMux I__5528 (
            .O(N__31935),
            .I(N__31849));
    InMux I__5527 (
            .O(N__31934),
            .I(N__31849));
    LocalMux I__5526 (
            .O(N__31927),
            .I(N__31840));
    LocalMux I__5525 (
            .O(N__31922),
            .I(N__31840));
    LocalMux I__5524 (
            .O(N__31917),
            .I(N__31840));
    InMux I__5523 (
            .O(N__31916),
            .I(N__31835));
    InMux I__5522 (
            .O(N__31915),
            .I(N__31835));
    InMux I__5521 (
            .O(N__31914),
            .I(N__31824));
    InMux I__5520 (
            .O(N__31913),
            .I(N__31824));
    InMux I__5519 (
            .O(N__31912),
            .I(N__31824));
    InMux I__5518 (
            .O(N__31911),
            .I(N__31824));
    InMux I__5517 (
            .O(N__31910),
            .I(N__31824));
    LocalMux I__5516 (
            .O(N__31897),
            .I(N__31817));
    LocalMux I__5515 (
            .O(N__31892),
            .I(N__31817));
    Span4Mux_v I__5514 (
            .O(N__31889),
            .I(N__31817));
    Span4Mux_h I__5513 (
            .O(N__31886),
            .I(N__31814));
    InMux I__5512 (
            .O(N__31885),
            .I(N__31805));
    InMux I__5511 (
            .O(N__31884),
            .I(N__31805));
    InMux I__5510 (
            .O(N__31883),
            .I(N__31805));
    InMux I__5509 (
            .O(N__31882),
            .I(N__31805));
    LocalMux I__5508 (
            .O(N__31873),
            .I(N__31798));
    LocalMux I__5507 (
            .O(N__31866),
            .I(N__31798));
    LocalMux I__5506 (
            .O(N__31849),
            .I(N__31798));
    InMux I__5505 (
            .O(N__31848),
            .I(N__31793));
    InMux I__5504 (
            .O(N__31847),
            .I(N__31793));
    Span4Mux_v I__5503 (
            .O(N__31840),
            .I(N__31788));
    LocalMux I__5502 (
            .O(N__31835),
            .I(N__31788));
    LocalMux I__5501 (
            .O(N__31824),
            .I(un1_sacqtime_cry_23_THRU_CO));
    Odrv4 I__5500 (
            .O(N__31817),
            .I(un1_sacqtime_cry_23_THRU_CO));
    Odrv4 I__5499 (
            .O(N__31814),
            .I(un1_sacqtime_cry_23_THRU_CO));
    LocalMux I__5498 (
            .O(N__31805),
            .I(un1_sacqtime_cry_23_THRU_CO));
    Odrv12 I__5497 (
            .O(N__31798),
            .I(un1_sacqtime_cry_23_THRU_CO));
    LocalMux I__5496 (
            .O(N__31793),
            .I(un1_sacqtime_cry_23_THRU_CO));
    Odrv4 I__5495 (
            .O(N__31788),
            .I(un1_sacqtime_cry_23_THRU_CO));
    IoInMux I__5494 (
            .O(N__31773),
            .I(N__31770));
    LocalMux I__5493 (
            .O(N__31770),
            .I(N__31767));
    IoSpan4Mux I__5492 (
            .O(N__31767),
            .I(N__31764));
    Span4Mux_s2_h I__5491 (
            .O(N__31764),
            .I(N__31761));
    Sp12to4 I__5490 (
            .O(N__31761),
            .I(N__31758));
    Span12Mux_h I__5489 (
            .O(N__31758),
            .I(N__31754));
    InMux I__5488 (
            .O(N__31757),
            .I(N__31751));
    Odrv12 I__5487 (
            .O(N__31754),
            .I(RAM_DATA_cl_7Z0Z_15));
    LocalMux I__5486 (
            .O(N__31751),
            .I(RAM_DATA_cl_7Z0Z_15));
    IoInMux I__5485 (
            .O(N__31746),
            .I(N__31743));
    LocalMux I__5484 (
            .O(N__31743),
            .I(N__31740));
    IoSpan4Mux I__5483 (
            .O(N__31740),
            .I(N__31737));
    IoSpan4Mux I__5482 (
            .O(N__31737),
            .I(N__31734));
    Span4Mux_s2_h I__5481 (
            .O(N__31734),
            .I(N__31731));
    Sp12to4 I__5480 (
            .O(N__31731),
            .I(N__31728));
    Span12Mux_h I__5479 (
            .O(N__31728),
            .I(N__31725));
    Span12Mux_v I__5478 (
            .O(N__31725),
            .I(N__31721));
    InMux I__5477 (
            .O(N__31724),
            .I(N__31718));
    Odrv12 I__5476 (
            .O(N__31721),
            .I(RAM_DATA_cl_4Z0Z_15));
    LocalMux I__5475 (
            .O(N__31718),
            .I(RAM_DATA_cl_4Z0Z_15));
    InMux I__5474 (
            .O(N__31713),
            .I(N__31698));
    InMux I__5473 (
            .O(N__31712),
            .I(N__31698));
    InMux I__5472 (
            .O(N__31711),
            .I(N__31698));
    InMux I__5471 (
            .O(N__31710),
            .I(N__31698));
    InMux I__5470 (
            .O(N__31709),
            .I(N__31686));
    InMux I__5469 (
            .O(N__31708),
            .I(N__31686));
    InMux I__5468 (
            .O(N__31707),
            .I(N__31686));
    LocalMux I__5467 (
            .O(N__31698),
            .I(N__31680));
    InMux I__5466 (
            .O(N__31697),
            .I(N__31671));
    InMux I__5465 (
            .O(N__31696),
            .I(N__31671));
    InMux I__5464 (
            .O(N__31695),
            .I(N__31671));
    InMux I__5463 (
            .O(N__31694),
            .I(N__31671));
    InMux I__5462 (
            .O(N__31693),
            .I(N__31666));
    LocalMux I__5461 (
            .O(N__31686),
            .I(N__31663));
    InMux I__5460 (
            .O(N__31685),
            .I(N__31656));
    InMux I__5459 (
            .O(N__31684),
            .I(N__31656));
    InMux I__5458 (
            .O(N__31683),
            .I(N__31656));
    Span4Mux_h I__5457 (
            .O(N__31680),
            .I(N__31653));
    LocalMux I__5456 (
            .O(N__31671),
            .I(N__31650));
    InMux I__5455 (
            .O(N__31670),
            .I(N__31645));
    InMux I__5454 (
            .O(N__31669),
            .I(N__31645));
    LocalMux I__5453 (
            .O(N__31666),
            .I(N__31642));
    Odrv4 I__5452 (
            .O(N__31663),
            .I(N_71));
    LocalMux I__5451 (
            .O(N__31656),
            .I(N_71));
    Odrv4 I__5450 (
            .O(N__31653),
            .I(N_71));
    Odrv4 I__5449 (
            .O(N__31650),
            .I(N_71));
    LocalMux I__5448 (
            .O(N__31645),
            .I(N_71));
    Odrv4 I__5447 (
            .O(N__31642),
            .I(N_71));
    InMux I__5446 (
            .O(N__31629),
            .I(N__31626));
    LocalMux I__5445 (
            .O(N__31626),
            .I(N_105));
    CascadeMux I__5444 (
            .O(N__31623),
            .I(N__31620));
    InMux I__5443 (
            .O(N__31620),
            .I(N__31616));
    InMux I__5442 (
            .O(N__31619),
            .I(N__31613));
    LocalMux I__5441 (
            .O(N__31616),
            .I(sRAM_pointer_writeZ0Z_0));
    LocalMux I__5440 (
            .O(N__31613),
            .I(sRAM_pointer_writeZ0Z_0));
    InMux I__5439 (
            .O(N__31608),
            .I(bfn_13_18_0_));
    CascadeMux I__5438 (
            .O(N__31605),
            .I(N__31602));
    InMux I__5437 (
            .O(N__31602),
            .I(N__31598));
    InMux I__5436 (
            .O(N__31601),
            .I(N__31595));
    LocalMux I__5435 (
            .O(N__31598),
            .I(sRAM_pointer_writeZ0Z_1));
    LocalMux I__5434 (
            .O(N__31595),
            .I(sRAM_pointer_writeZ0Z_1));
    InMux I__5433 (
            .O(N__31590),
            .I(N__31587));
    LocalMux I__5432 (
            .O(N__31587),
            .I(N__31584));
    Sp12to4 I__5431 (
            .O(N__31584),
            .I(N__31581));
    Span12Mux_v I__5430 (
            .O(N__31581),
            .I(N__31578));
    Span12Mux_h I__5429 (
            .O(N__31578),
            .I(N__31575));
    Odrv12 I__5428 (
            .O(N__31575),
            .I(ADC4_c));
    IoInMux I__5427 (
            .O(N__31572),
            .I(N__31569));
    LocalMux I__5426 (
            .O(N__31569),
            .I(N__31566));
    Span4Mux_s2_v I__5425 (
            .O(N__31566),
            .I(N__31563));
    Sp12to4 I__5424 (
            .O(N__31563),
            .I(N__31560));
    Span12Mux_h I__5423 (
            .O(N__31560),
            .I(N__31557));
    Odrv12 I__5422 (
            .O(N__31557),
            .I(RAM_DATA_1Z0Z_4));
    InMux I__5421 (
            .O(N__31554),
            .I(N__31551));
    LocalMux I__5420 (
            .O(N__31551),
            .I(N__31548));
    Span12Mux_s11_v I__5419 (
            .O(N__31548),
            .I(N__31545));
    Span12Mux_h I__5418 (
            .O(N__31545),
            .I(N__31542));
    Odrv12 I__5417 (
            .O(N__31542),
            .I(ADC6_c));
    IoInMux I__5416 (
            .O(N__31539),
            .I(N__31536));
    LocalMux I__5415 (
            .O(N__31536),
            .I(N__31533));
    Span4Mux_s1_v I__5414 (
            .O(N__31533),
            .I(N__31530));
    Sp12to4 I__5413 (
            .O(N__31530),
            .I(N__31527));
    Span12Mux_h I__5412 (
            .O(N__31527),
            .I(N__31524));
    Odrv12 I__5411 (
            .O(N__31524),
            .I(RAM_DATA_1Z0Z_6));
    InMux I__5410 (
            .O(N__31521),
            .I(N__31518));
    LocalMux I__5409 (
            .O(N__31518),
            .I(N__31515));
    Span4Mux_v I__5408 (
            .O(N__31515),
            .I(N__31512));
    Sp12to4 I__5407 (
            .O(N__31512),
            .I(N__31509));
    Span12Mux_h I__5406 (
            .O(N__31509),
            .I(N__31506));
    Span12Mux_h I__5405 (
            .O(N__31506),
            .I(N__31503));
    Odrv12 I__5404 (
            .O(N__31503),
            .I(ADC9_c));
    IoInMux I__5403 (
            .O(N__31500),
            .I(N__31497));
    LocalMux I__5402 (
            .O(N__31497),
            .I(N__31494));
    Span4Mux_s3_h I__5401 (
            .O(N__31494),
            .I(N__31491));
    Sp12to4 I__5400 (
            .O(N__31491),
            .I(N__31488));
    Span12Mux_s7_v I__5399 (
            .O(N__31488),
            .I(N__31485));
    Span12Mux_h I__5398 (
            .O(N__31485),
            .I(N__31482));
    Span12Mux_v I__5397 (
            .O(N__31482),
            .I(N__31479));
    Odrv12 I__5396 (
            .O(N__31479),
            .I(RAM_DATA_1Z0Z_10));
    InMux I__5395 (
            .O(N__31476),
            .I(N__31473));
    LocalMux I__5394 (
            .O(N__31473),
            .I(N__31470));
    Span4Mux_v I__5393 (
            .O(N__31470),
            .I(N__31467));
    Sp12to4 I__5392 (
            .O(N__31467),
            .I(N__31464));
    Span12Mux_h I__5391 (
            .O(N__31464),
            .I(N__31461));
    Span12Mux_v I__5390 (
            .O(N__31461),
            .I(N__31458));
    Odrv12 I__5389 (
            .O(N__31458),
            .I(top_tour1_c));
    IoInMux I__5388 (
            .O(N__31455),
            .I(N__31452));
    LocalMux I__5387 (
            .O(N__31452),
            .I(N__31449));
    IoSpan4Mux I__5386 (
            .O(N__31449),
            .I(N__31446));
    Span4Mux_s1_h I__5385 (
            .O(N__31446),
            .I(N__31443));
    Sp12to4 I__5384 (
            .O(N__31443),
            .I(N__31440));
    Span12Mux_h I__5383 (
            .O(N__31440),
            .I(N__31437));
    Odrv12 I__5382 (
            .O(N__31437),
            .I(RAM_DATA_1Z0Z_11));
    InMux I__5381 (
            .O(N__31434),
            .I(N__31431));
    LocalMux I__5380 (
            .O(N__31431),
            .I(N__31428));
    Sp12to4 I__5379 (
            .O(N__31428),
            .I(N__31425));
    Span12Mux_s9_v I__5378 (
            .O(N__31425),
            .I(N__31422));
    Span12Mux_v I__5377 (
            .O(N__31422),
            .I(N__31419));
    Span12Mux_h I__5376 (
            .O(N__31419),
            .I(N__31416));
    Odrv12 I__5375 (
            .O(N__31416),
            .I(top_tour2_c));
    IoInMux I__5374 (
            .O(N__31413),
            .I(N__31410));
    LocalMux I__5373 (
            .O(N__31410),
            .I(N__31407));
    IoSpan4Mux I__5372 (
            .O(N__31407),
            .I(N__31404));
    IoSpan4Mux I__5371 (
            .O(N__31404),
            .I(N__31401));
    Span4Mux_s2_h I__5370 (
            .O(N__31401),
            .I(N__31398));
    Sp12to4 I__5369 (
            .O(N__31398),
            .I(N__31395));
    Odrv12 I__5368 (
            .O(N__31395),
            .I(RAM_DATA_1Z0Z_12));
    InMux I__5367 (
            .O(N__31392),
            .I(N__31380));
    InMux I__5366 (
            .O(N__31391),
            .I(N__31380));
    InMux I__5365 (
            .O(N__31390),
            .I(N__31380));
    InMux I__5364 (
            .O(N__31389),
            .I(N__31376));
    InMux I__5363 (
            .O(N__31388),
            .I(N__31373));
    InMux I__5362 (
            .O(N__31387),
            .I(N__31370));
    LocalMux I__5361 (
            .O(N__31380),
            .I(N__31367));
    InMux I__5360 (
            .O(N__31379),
            .I(N__31364));
    LocalMux I__5359 (
            .O(N__31376),
            .I(N__31360));
    LocalMux I__5358 (
            .O(N__31373),
            .I(N__31351));
    LocalMux I__5357 (
            .O(N__31370),
            .I(N__31351));
    Span4Mux_v I__5356 (
            .O(N__31367),
            .I(N__31351));
    LocalMux I__5355 (
            .O(N__31364),
            .I(N__31351));
    InMux I__5354 (
            .O(N__31363),
            .I(N__31346));
    Span4Mux_h I__5353 (
            .O(N__31360),
            .I(N__31343));
    Span4Mux_h I__5352 (
            .O(N__31351),
            .I(N__31340));
    InMux I__5351 (
            .O(N__31350),
            .I(N__31337));
    InMux I__5350 (
            .O(N__31349),
            .I(N__31334));
    LocalMux I__5349 (
            .O(N__31346),
            .I(N__31331));
    Span4Mux_h I__5348 (
            .O(N__31343),
            .I(N__31326));
    Span4Mux_v I__5347 (
            .O(N__31340),
            .I(N__31326));
    LocalMux I__5346 (
            .O(N__31337),
            .I(sTrigCounterZ0Z_0));
    LocalMux I__5345 (
            .O(N__31334),
            .I(sTrigCounterZ0Z_0));
    Odrv4 I__5344 (
            .O(N__31331),
            .I(sTrigCounterZ0Z_0));
    Odrv4 I__5343 (
            .O(N__31326),
            .I(sTrigCounterZ0Z_0));
    IoInMux I__5342 (
            .O(N__31317),
            .I(N__31314));
    LocalMux I__5341 (
            .O(N__31314),
            .I(N__31311));
    Span12Mux_s3_h I__5340 (
            .O(N__31311),
            .I(N__31308));
    Span12Mux_h I__5339 (
            .O(N__31308),
            .I(N__31305));
    Odrv12 I__5338 (
            .O(N__31305),
            .I(RAM_DATA_1Z0Z_13));
    CascadeMux I__5337 (
            .O(N__31302),
            .I(N__31294));
    InMux I__5336 (
            .O(N__31301),
            .I(N__31290));
    InMux I__5335 (
            .O(N__31300),
            .I(N__31287));
    InMux I__5334 (
            .O(N__31299),
            .I(N__31284));
    InMux I__5333 (
            .O(N__31298),
            .I(N__31281));
    InMux I__5332 (
            .O(N__31297),
            .I(N__31273));
    InMux I__5331 (
            .O(N__31294),
            .I(N__31273));
    InMux I__5330 (
            .O(N__31293),
            .I(N__31273));
    LocalMux I__5329 (
            .O(N__31290),
            .I(N__31270));
    LocalMux I__5328 (
            .O(N__31287),
            .I(N__31263));
    LocalMux I__5327 (
            .O(N__31284),
            .I(N__31263));
    LocalMux I__5326 (
            .O(N__31281),
            .I(N__31263));
    InMux I__5325 (
            .O(N__31280),
            .I(N__31259));
    LocalMux I__5324 (
            .O(N__31273),
            .I(N__31256));
    Span4Mux_h I__5323 (
            .O(N__31270),
            .I(N__31253));
    Span4Mux_h I__5322 (
            .O(N__31263),
            .I(N__31250));
    InMux I__5321 (
            .O(N__31262),
            .I(N__31247));
    LocalMux I__5320 (
            .O(N__31259),
            .I(N__31242));
    Span4Mux_h I__5319 (
            .O(N__31256),
            .I(N__31242));
    Span4Mux_h I__5318 (
            .O(N__31253),
            .I(N__31237));
    Span4Mux_v I__5317 (
            .O(N__31250),
            .I(N__31237));
    LocalMux I__5316 (
            .O(N__31247),
            .I(sTrigCounterZ0Z_1));
    Odrv4 I__5315 (
            .O(N__31242),
            .I(sTrigCounterZ0Z_1));
    Odrv4 I__5314 (
            .O(N__31237),
            .I(sTrigCounterZ0Z_1));
    IoInMux I__5313 (
            .O(N__31230),
            .I(N__31227));
    LocalMux I__5312 (
            .O(N__31227),
            .I(N__31224));
    Span12Mux_s3_h I__5311 (
            .O(N__31224),
            .I(N__31221));
    Span12Mux_h I__5310 (
            .O(N__31221),
            .I(N__31218));
    Odrv12 I__5309 (
            .O(N__31218),
            .I(RAM_DATA_1Z0Z_14));
    InMux I__5308 (
            .O(N__31215),
            .I(N__31212));
    LocalMux I__5307 (
            .O(N__31212),
            .I(N__31209));
    Span4Mux_v I__5306 (
            .O(N__31209),
            .I(N__31206));
    Sp12to4 I__5305 (
            .O(N__31206),
            .I(N__31203));
    Span12Mux_h I__5304 (
            .O(N__31203),
            .I(N__31200));
    Odrv12 I__5303 (
            .O(N__31200),
            .I(ADC2_c));
    IoInMux I__5302 (
            .O(N__31197),
            .I(N__31194));
    LocalMux I__5301 (
            .O(N__31194),
            .I(N__31191));
    Span12Mux_s3_v I__5300 (
            .O(N__31191),
            .I(N__31188));
    Span12Mux_h I__5299 (
            .O(N__31188),
            .I(N__31185));
    Odrv12 I__5298 (
            .O(N__31185),
            .I(RAM_DATA_1Z0Z_2));
    CEMux I__5297 (
            .O(N__31182),
            .I(N__31178));
    CEMux I__5296 (
            .O(N__31181),
            .I(N__31175));
    LocalMux I__5295 (
            .O(N__31178),
            .I(N_31_i));
    LocalMux I__5294 (
            .O(N__31175),
            .I(N_31_i));
    CEMux I__5293 (
            .O(N__31170),
            .I(N__31167));
    LocalMux I__5292 (
            .O(N__31167),
            .I(N__31164));
    Span12Mux_v I__5291 (
            .O(N__31164),
            .I(N__31161));
    Odrv12 I__5290 (
            .O(N__31161),
            .I(sAddress_RNIA6242Z0Z_2));
    InMux I__5289 (
            .O(N__31158),
            .I(N__31155));
    LocalMux I__5288 (
            .O(N__31155),
            .I(sDAC_mem_19Z0Z_4));
    InMux I__5287 (
            .O(N__31152),
            .I(N__31149));
    LocalMux I__5286 (
            .O(N__31149),
            .I(sDAC_mem_18Z0Z_4));
    InMux I__5285 (
            .O(N__31146),
            .I(N__31143));
    LocalMux I__5284 (
            .O(N__31143),
            .I(sDAC_mem_19Z0Z_5));
    InMux I__5283 (
            .O(N__31140),
            .I(N__31137));
    LocalMux I__5282 (
            .O(N__31137),
            .I(sDAC_mem_18Z0Z_5));
    InMux I__5281 (
            .O(N__31134),
            .I(N__31131));
    LocalMux I__5280 (
            .O(N__31131),
            .I(sDAC_mem_19Z0Z_6));
    InMux I__5279 (
            .O(N__31128),
            .I(N__31125));
    LocalMux I__5278 (
            .O(N__31125),
            .I(sDAC_mem_18Z0Z_6));
    CEMux I__5277 (
            .O(N__31122),
            .I(N__31119));
    LocalMux I__5276 (
            .O(N__31119),
            .I(N__31116));
    Odrv4 I__5275 (
            .O(N__31116),
            .I(sDAC_mem_19_1_sqmuxa));
    CEMux I__5274 (
            .O(N__31113),
            .I(N__31110));
    LocalMux I__5273 (
            .O(N__31110),
            .I(sDAC_mem_32_1_sqmuxa));
    InMux I__5272 (
            .O(N__31107),
            .I(N__31101));
    InMux I__5271 (
            .O(N__31106),
            .I(N__31098));
    InMux I__5270 (
            .O(N__31105),
            .I(N__31095));
    InMux I__5269 (
            .O(N__31104),
            .I(N__31091));
    LocalMux I__5268 (
            .O(N__31101),
            .I(N__31087));
    LocalMux I__5267 (
            .O(N__31098),
            .I(N__31084));
    LocalMux I__5266 (
            .O(N__31095),
            .I(N__31081));
    InMux I__5265 (
            .O(N__31094),
            .I(N__31078));
    LocalMux I__5264 (
            .O(N__31091),
            .I(N__31075));
    InMux I__5263 (
            .O(N__31090),
            .I(N__31067));
    Span4Mux_h I__5262 (
            .O(N__31087),
            .I(N__31064));
    Span4Mux_v I__5261 (
            .O(N__31084),
            .I(N__31059));
    Span4Mux_v I__5260 (
            .O(N__31081),
            .I(N__31059));
    LocalMux I__5259 (
            .O(N__31078),
            .I(N__31056));
    Span4Mux_h I__5258 (
            .O(N__31075),
            .I(N__31053));
    InMux I__5257 (
            .O(N__31074),
            .I(N__31048));
    InMux I__5256 (
            .O(N__31073),
            .I(N__31048));
    InMux I__5255 (
            .O(N__31072),
            .I(N__31045));
    InMux I__5254 (
            .O(N__31071),
            .I(N__31040));
    InMux I__5253 (
            .O(N__31070),
            .I(N__31040));
    LocalMux I__5252 (
            .O(N__31067),
            .I(N__31037));
    Odrv4 I__5251 (
            .O(N__31064),
            .I(N_141));
    Odrv4 I__5250 (
            .O(N__31059),
            .I(N_141));
    Odrv4 I__5249 (
            .O(N__31056),
            .I(N_141));
    Odrv4 I__5248 (
            .O(N__31053),
            .I(N_141));
    LocalMux I__5247 (
            .O(N__31048),
            .I(N_141));
    LocalMux I__5246 (
            .O(N__31045),
            .I(N_141));
    LocalMux I__5245 (
            .O(N__31040),
            .I(N_141));
    Odrv4 I__5244 (
            .O(N__31037),
            .I(N_141));
    CEMux I__5243 (
            .O(N__31020),
            .I(N__31017));
    LocalMux I__5242 (
            .O(N__31017),
            .I(N__31013));
    CEMux I__5241 (
            .O(N__31016),
            .I(N__31010));
    Span4Mux_h I__5240 (
            .O(N__31013),
            .I(N__31005));
    LocalMux I__5239 (
            .O(N__31010),
            .I(N__31005));
    Span4Mux_h I__5238 (
            .O(N__31005),
            .I(N__31002));
    Odrv4 I__5237 (
            .O(N__31002),
            .I(sEETrigCounter_1_sqmuxa));
    CascadeMux I__5236 (
            .O(N__30999),
            .I(N_1480_cascade_));
    InMux I__5235 (
            .O(N__30996),
            .I(N__30993));
    LocalMux I__5234 (
            .O(N__30993),
            .I(N__30988));
    InMux I__5233 (
            .O(N__30992),
            .I(N__30985));
    InMux I__5232 (
            .O(N__30991),
            .I(N__30982));
    Odrv4 I__5231 (
            .O(N__30988),
            .I(un1_spointer11_5_0_2));
    LocalMux I__5230 (
            .O(N__30985),
            .I(un1_spointer11_5_0_2));
    LocalMux I__5229 (
            .O(N__30982),
            .I(un1_spointer11_5_0_2));
    CEMux I__5228 (
            .O(N__30975),
            .I(N__30972));
    LocalMux I__5227 (
            .O(N__30972),
            .I(N__30969));
    Span4Mux_v I__5226 (
            .O(N__30969),
            .I(N__30966));
    Odrv4 I__5225 (
            .O(N__30966),
            .I(sAddress_RNIA6242_2Z0Z_2));
    CascadeMux I__5224 (
            .O(N__30963),
            .I(N_280_cascade_));
    CEMux I__5223 (
            .O(N__30960),
            .I(N__30957));
    LocalMux I__5222 (
            .O(N__30957),
            .I(sDAC_mem_17_1_sqmuxa));
    InMux I__5221 (
            .O(N__30954),
            .I(N__30951));
    LocalMux I__5220 (
            .O(N__30951),
            .I(N__30948));
    Span4Mux_v I__5219 (
            .O(N__30948),
            .I(N__30943));
    InMux I__5218 (
            .O(N__30947),
            .I(N__30938));
    InMux I__5217 (
            .O(N__30946),
            .I(N__30938));
    Odrv4 I__5216 (
            .O(N__30943),
            .I(sAddressZ0Z_6));
    LocalMux I__5215 (
            .O(N__30938),
            .I(sAddressZ0Z_6));
    CascadeMux I__5214 (
            .O(N__30933),
            .I(N__30930));
    InMux I__5213 (
            .O(N__30930),
            .I(N__30927));
    LocalMux I__5212 (
            .O(N__30927),
            .I(N__30923));
    CascadeMux I__5211 (
            .O(N__30926),
            .I(N__30919));
    Span4Mux_h I__5210 (
            .O(N__30923),
            .I(N__30916));
    InMux I__5209 (
            .O(N__30922),
            .I(N__30911));
    InMux I__5208 (
            .O(N__30919),
            .I(N__30911));
    Odrv4 I__5207 (
            .O(N__30916),
            .I(sAddressZ0Z_7));
    LocalMux I__5206 (
            .O(N__30911),
            .I(sAddressZ0Z_7));
    InMux I__5205 (
            .O(N__30906),
            .I(N__30903));
    LocalMux I__5204 (
            .O(N__30903),
            .I(sEEPonPoff_1_sqmuxa_0_a2_1));
    CEMux I__5203 (
            .O(N__30900),
            .I(N__30897));
    LocalMux I__5202 (
            .O(N__30897),
            .I(N__30893));
    CEMux I__5201 (
            .O(N__30896),
            .I(N__30890));
    Span4Mux_h I__5200 (
            .O(N__30893),
            .I(N__30887));
    LocalMux I__5199 (
            .O(N__30890),
            .I(N__30884));
    Span4Mux_h I__5198 (
            .O(N__30887),
            .I(N__30881));
    Sp12to4 I__5197 (
            .O(N__30884),
            .I(N__30878));
    Odrv4 I__5196 (
            .O(N__30881),
            .I(sEEPon_1_sqmuxa));
    Odrv12 I__5195 (
            .O(N__30878),
            .I(sEEPon_1_sqmuxa));
    InMux I__5194 (
            .O(N__30873),
            .I(N__30861));
    InMux I__5193 (
            .O(N__30872),
            .I(N__30861));
    InMux I__5192 (
            .O(N__30871),
            .I(N__30861));
    InMux I__5191 (
            .O(N__30870),
            .I(N__30861));
    LocalMux I__5190 (
            .O(N__30861),
            .I(N_291));
    CEMux I__5189 (
            .O(N__30858),
            .I(N__30855));
    LocalMux I__5188 (
            .O(N__30855),
            .I(N__30852));
    Odrv4 I__5187 (
            .O(N__30852),
            .I(sDAC_mem_33_1_sqmuxa));
    InMux I__5186 (
            .O(N__30849),
            .I(N__30846));
    LocalMux I__5185 (
            .O(N__30846),
            .I(sDAC_mem_23Z0Z_2));
    InMux I__5184 (
            .O(N__30843),
            .I(N__30840));
    LocalMux I__5183 (
            .O(N__30840),
            .I(sDAC_mem_22Z0Z_2));
    InMux I__5182 (
            .O(N__30837),
            .I(N__30834));
    LocalMux I__5181 (
            .O(N__30834),
            .I(sDAC_mem_23Z0Z_3));
    InMux I__5180 (
            .O(N__30831),
            .I(N__30828));
    LocalMux I__5179 (
            .O(N__30828),
            .I(sDAC_mem_22Z0Z_3));
    InMux I__5178 (
            .O(N__30825),
            .I(N__30822));
    LocalMux I__5177 (
            .O(N__30822),
            .I(sDAC_mem_23Z0Z_4));
    InMux I__5176 (
            .O(N__30819),
            .I(N__30816));
    LocalMux I__5175 (
            .O(N__30816),
            .I(sDAC_mem_22Z0Z_4));
    CascadeMux I__5174 (
            .O(N__30813),
            .I(N_291_cascade_));
    CEMux I__5173 (
            .O(N__30810),
            .I(N__30807));
    LocalMux I__5172 (
            .O(N__30807),
            .I(N__30804));
    Span4Mux_h I__5171 (
            .O(N__30804),
            .I(N__30801));
    Span4Mux_h I__5170 (
            .O(N__30801),
            .I(N__30798));
    Odrv4 I__5169 (
            .O(N__30798),
            .I(sEEPonPoff_1_sqmuxa));
    InMux I__5168 (
            .O(N__30795),
            .I(N__30791));
    InMux I__5167 (
            .O(N__30794),
            .I(N__30788));
    LocalMux I__5166 (
            .O(N__30791),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0 ));
    LocalMux I__5165 (
            .O(N__30788),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0 ));
    InMux I__5164 (
            .O(N__30783),
            .I(N__30779));
    InMux I__5163 (
            .O(N__30782),
            .I(N__30776));
    LocalMux I__5162 (
            .O(N__30779),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1 ));
    LocalMux I__5161 (
            .O(N__30776),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1 ));
    InMux I__5160 (
            .O(N__30771),
            .I(N__30767));
    InMux I__5159 (
            .O(N__30770),
            .I(N__30764));
    LocalMux I__5158 (
            .O(N__30767),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2 ));
    LocalMux I__5157 (
            .O(N__30764),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2 ));
    InMux I__5156 (
            .O(N__30759),
            .I(N__30755));
    InMux I__5155 (
            .O(N__30758),
            .I(N__30752));
    LocalMux I__5154 (
            .O(N__30755),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3 ));
    LocalMux I__5153 (
            .O(N__30752),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3 ));
    InMux I__5152 (
            .O(N__30747),
            .I(N__30743));
    InMux I__5151 (
            .O(N__30746),
            .I(N__30740));
    LocalMux I__5150 (
            .O(N__30743),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4 ));
    LocalMux I__5149 (
            .O(N__30740),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4 ));
    InMux I__5148 (
            .O(N__30735),
            .I(N__30731));
    InMux I__5147 (
            .O(N__30734),
            .I(N__30728));
    LocalMux I__5146 (
            .O(N__30731),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5 ));
    LocalMux I__5145 (
            .O(N__30728),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5 ));
    InMux I__5144 (
            .O(N__30723),
            .I(N__30719));
    InMux I__5143 (
            .O(N__30722),
            .I(N__30716));
    LocalMux I__5142 (
            .O(N__30719),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6 ));
    LocalMux I__5141 (
            .O(N__30716),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6 ));
    InMux I__5140 (
            .O(N__30711),
            .I(N__30708));
    LocalMux I__5139 (
            .O(N__30708),
            .I(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7 ));
    ClkMux I__5138 (
            .O(N__30705),
            .I(N__30678));
    ClkMux I__5137 (
            .O(N__30704),
            .I(N__30678));
    ClkMux I__5136 (
            .O(N__30703),
            .I(N__30678));
    ClkMux I__5135 (
            .O(N__30702),
            .I(N__30678));
    ClkMux I__5134 (
            .O(N__30701),
            .I(N__30678));
    ClkMux I__5133 (
            .O(N__30700),
            .I(N__30678));
    ClkMux I__5132 (
            .O(N__30699),
            .I(N__30678));
    ClkMux I__5131 (
            .O(N__30698),
            .I(N__30678));
    ClkMux I__5130 (
            .O(N__30697),
            .I(N__30678));
    GlobalMux I__5129 (
            .O(N__30678),
            .I(N__30675));
    gio2CtrlBuf I__5128 (
            .O(N__30675),
            .I(spi_sclk_g));
    CEMux I__5127 (
            .O(N__30672),
            .I(N__30668));
    CEMux I__5126 (
            .O(N__30671),
            .I(N__30665));
    LocalMux I__5125 (
            .O(N__30668),
            .I(N__30661));
    LocalMux I__5124 (
            .O(N__30665),
            .I(N__30658));
    CEMux I__5123 (
            .O(N__30664),
            .I(N__30655));
    Span4Mux_h I__5122 (
            .O(N__30661),
            .I(N__30652));
    Span4Mux_h I__5121 (
            .O(N__30658),
            .I(N__30649));
    LocalMux I__5120 (
            .O(N__30655),
            .I(N__30646));
    Odrv4 I__5119 (
            .O(N__30652),
            .I(\spi_slave_inst.spi_cs_iZ0 ));
    Odrv4 I__5118 (
            .O(N__30649),
            .I(\spi_slave_inst.spi_cs_iZ0 ));
    Odrv4 I__5117 (
            .O(N__30646),
            .I(\spi_slave_inst.spi_cs_iZ0 ));
    InMux I__5116 (
            .O(N__30639),
            .I(N__30636));
    LocalMux I__5115 (
            .O(N__30636),
            .I(N__30633));
    Span12Mux_s11_v I__5114 (
            .O(N__30633),
            .I(N__30630));
    Span12Mux_h I__5113 (
            .O(N__30630),
            .I(N__30627));
    Odrv12 I__5112 (
            .O(N__30627),
            .I(ADC8_c));
    IoInMux I__5111 (
            .O(N__30624),
            .I(N__30621));
    LocalMux I__5110 (
            .O(N__30621),
            .I(N__30618));
    IoSpan4Mux I__5109 (
            .O(N__30618),
            .I(N__30615));
    Span4Mux_s3_h I__5108 (
            .O(N__30615),
            .I(N__30612));
    Sp12to4 I__5107 (
            .O(N__30612),
            .I(N__30609));
    Span12Mux_h I__5106 (
            .O(N__30609),
            .I(N__30606));
    Span12Mux_v I__5105 (
            .O(N__30606),
            .I(N__30603));
    Odrv12 I__5104 (
            .O(N__30603),
            .I(RAM_DATA_1Z0Z_9));
    IoInMux I__5103 (
            .O(N__30600),
            .I(N__30597));
    LocalMux I__5102 (
            .O(N__30597),
            .I(N__30594));
    Span4Mux_s2_h I__5101 (
            .O(N__30594),
            .I(N__30591));
    Sp12to4 I__5100 (
            .O(N__30591),
            .I(N__30588));
    Span12Mux_v I__5099 (
            .O(N__30588),
            .I(N__30585));
    Span12Mux_h I__5098 (
            .O(N__30585),
            .I(N__30582));
    Odrv12 I__5097 (
            .O(N__30582),
            .I(RAM_DATA_1Z0Z_15));
    IoInMux I__5096 (
            .O(N__30579),
            .I(N__30576));
    LocalMux I__5095 (
            .O(N__30576),
            .I(N__30573));
    IoSpan4Mux I__5094 (
            .O(N__30573),
            .I(N__30570));
    Span4Mux_s1_v I__5093 (
            .O(N__30570),
            .I(N__30567));
    Sp12to4 I__5092 (
            .O(N__30567),
            .I(N__30564));
    Span12Mux_h I__5091 (
            .O(N__30564),
            .I(N__30561));
    Odrv12 I__5090 (
            .O(N__30561),
            .I(RAM_DATA_1Z0Z_7));
    IoInMux I__5089 (
            .O(N__30558),
            .I(N__30555));
    LocalMux I__5088 (
            .O(N__30555),
            .I(N__30552));
    Span4Mux_s2_v I__5087 (
            .O(N__30552),
            .I(N__30549));
    Span4Mux_h I__5086 (
            .O(N__30549),
            .I(N__30546));
    Span4Mux_h I__5085 (
            .O(N__30546),
            .I(N__30543));
    Span4Mux_h I__5084 (
            .O(N__30543),
            .I(N__30540));
    Span4Mux_v I__5083 (
            .O(N__30540),
            .I(N__30536));
    InMux I__5082 (
            .O(N__30539),
            .I(N__30533));
    Odrv4 I__5081 (
            .O(N__30536),
            .I(RAM_DATA_cl_1Z0Z_15));
    LocalMux I__5080 (
            .O(N__30533),
            .I(RAM_DATA_cl_1Z0Z_15));
    InMux I__5079 (
            .O(N__30528),
            .I(N__30525));
    LocalMux I__5078 (
            .O(N__30525),
            .I(N_100));
    IoInMux I__5077 (
            .O(N__30522),
            .I(N__30519));
    LocalMux I__5076 (
            .O(N__30519),
            .I(N__30516));
    IoSpan4Mux I__5075 (
            .O(N__30516),
            .I(N__30513));
    IoSpan4Mux I__5074 (
            .O(N__30513),
            .I(N__30510));
    Span4Mux_s3_h I__5073 (
            .O(N__30510),
            .I(N__30507));
    Sp12to4 I__5072 (
            .O(N__30507),
            .I(N__30504));
    Span12Mux_h I__5071 (
            .O(N__30504),
            .I(N__30500));
    InMux I__5070 (
            .O(N__30503),
            .I(N__30497));
    Odrv12 I__5069 (
            .O(N__30500),
            .I(RAM_DATA_cl_13Z0Z_15));
    LocalMux I__5068 (
            .O(N__30497),
            .I(RAM_DATA_cl_13Z0Z_15));
    InMux I__5067 (
            .O(N__30492),
            .I(N__30489));
    LocalMux I__5066 (
            .O(N__30489),
            .I(N_97));
    IoInMux I__5065 (
            .O(N__30486),
            .I(N__30483));
    LocalMux I__5064 (
            .O(N__30483),
            .I(N__30480));
    IoSpan4Mux I__5063 (
            .O(N__30480),
            .I(N__30477));
    IoSpan4Mux I__5062 (
            .O(N__30477),
            .I(N__30474));
    Sp12to4 I__5061 (
            .O(N__30474),
            .I(N__30471));
    Span12Mux_s7_h I__5060 (
            .O(N__30471),
            .I(N__30467));
    InMux I__5059 (
            .O(N__30470),
            .I(N__30464));
    Odrv12 I__5058 (
            .O(N__30467),
            .I(RAM_DATA_cl_2Z0Z_15));
    LocalMux I__5057 (
            .O(N__30464),
            .I(RAM_DATA_cl_2Z0Z_15));
    InMux I__5056 (
            .O(N__30459),
            .I(N__30456));
    LocalMux I__5055 (
            .O(N__30456),
            .I(N_101));
    InMux I__5054 (
            .O(N__30453),
            .I(N__30450));
    LocalMux I__5053 (
            .O(N__30450),
            .I(N_103));
    IoInMux I__5052 (
            .O(N__30447),
            .I(N__30444));
    LocalMux I__5051 (
            .O(N__30444),
            .I(N__30441));
    Span4Mux_s3_v I__5050 (
            .O(N__30441),
            .I(N__30438));
    Span4Mux_h I__5049 (
            .O(N__30438),
            .I(N__30435));
    Span4Mux_h I__5048 (
            .O(N__30435),
            .I(N__30432));
    Span4Mux_h I__5047 (
            .O(N__30432),
            .I(N__30428));
    InMux I__5046 (
            .O(N__30431),
            .I(N__30425));
    Odrv4 I__5045 (
            .O(N__30428),
            .I(RAM_DATA_cl_3Z0Z_15));
    LocalMux I__5044 (
            .O(N__30425),
            .I(RAM_DATA_cl_3Z0Z_15));
    InMux I__5043 (
            .O(N__30420),
            .I(N__30417));
    LocalMux I__5042 (
            .O(N__30417),
            .I(N__30414));
    Span12Mux_v I__5041 (
            .O(N__30414),
            .I(N__30411));
    Span12Mux_h I__5040 (
            .O(N__30411),
            .I(N__30408));
    Odrv12 I__5039 (
            .O(N__30408),
            .I(spi_mosi_ft_c));
    InMux I__5038 (
            .O(N__30405),
            .I(N__30402));
    LocalMux I__5037 (
            .O(N__30402),
            .I(N__30399));
    Span4Mux_v I__5036 (
            .O(N__30399),
            .I(N__30396));
    Sp12to4 I__5035 (
            .O(N__30396),
            .I(N__30393));
    Span12Mux_h I__5034 (
            .O(N__30393),
            .I(N__30389));
    InMux I__5033 (
            .O(N__30392),
            .I(N__30386));
    Odrv12 I__5032 (
            .O(N__30389),
            .I(sRAM_pointer_readZ0Z_11));
    LocalMux I__5031 (
            .O(N__30386),
            .I(sRAM_pointer_readZ0Z_11));
    IoInMux I__5030 (
            .O(N__30381),
            .I(N__30378));
    LocalMux I__5029 (
            .O(N__30378),
            .I(N__30375));
    IoSpan4Mux I__5028 (
            .O(N__30375),
            .I(N__30372));
    Span4Mux_s1_h I__5027 (
            .O(N__30372),
            .I(N__30369));
    Span4Mux_v I__5026 (
            .O(N__30369),
            .I(N__30366));
    Sp12to4 I__5025 (
            .O(N__30366),
            .I(N__30363));
    Span12Mux_v I__5024 (
            .O(N__30363),
            .I(N__30360));
    Span12Mux_h I__5023 (
            .O(N__30360),
            .I(N__30357));
    Odrv12 I__5022 (
            .O(N__30357),
            .I(RAM_ADD_c_11));
    CascadeMux I__5021 (
            .O(N__30354),
            .I(N__30351));
    InMux I__5020 (
            .O(N__30351),
            .I(N__30348));
    LocalMux I__5019 (
            .O(N__30348),
            .I(N__30345));
    Span4Mux_v I__5018 (
            .O(N__30345),
            .I(N__30342));
    Span4Mux_v I__5017 (
            .O(N__30342),
            .I(N__30339));
    Sp12to4 I__5016 (
            .O(N__30339),
            .I(N__30335));
    InMux I__5015 (
            .O(N__30338),
            .I(N__30332));
    Odrv12 I__5014 (
            .O(N__30335),
            .I(sRAM_pointer_readZ0Z_12));
    LocalMux I__5013 (
            .O(N__30332),
            .I(sRAM_pointer_readZ0Z_12));
    IoInMux I__5012 (
            .O(N__30327),
            .I(N__30324));
    LocalMux I__5011 (
            .O(N__30324),
            .I(N__30321));
    Span12Mux_s4_h I__5010 (
            .O(N__30321),
            .I(N__30318));
    Span12Mux_v I__5009 (
            .O(N__30318),
            .I(N__30315));
    Span12Mux_h I__5008 (
            .O(N__30315),
            .I(N__30312));
    Odrv12 I__5007 (
            .O(N__30312),
            .I(RAM_ADD_c_12));
    InMux I__5006 (
            .O(N__30309),
            .I(N__30306));
    LocalMux I__5005 (
            .O(N__30306),
            .I(N__30303));
    Span12Mux_h I__5004 (
            .O(N__30303),
            .I(N__30299));
    InMux I__5003 (
            .O(N__30302),
            .I(N__30296));
    Odrv12 I__5002 (
            .O(N__30299),
            .I(sRAM_pointer_readZ0Z_13));
    LocalMux I__5001 (
            .O(N__30296),
            .I(sRAM_pointer_readZ0Z_13));
    IoInMux I__5000 (
            .O(N__30291),
            .I(N__30288));
    LocalMux I__4999 (
            .O(N__30288),
            .I(N__30285));
    Span4Mux_s3_h I__4998 (
            .O(N__30285),
            .I(N__30282));
    Sp12to4 I__4997 (
            .O(N__30282),
            .I(N__30279));
    Span12Mux_s10_v I__4996 (
            .O(N__30279),
            .I(N__30276));
    Span12Mux_h I__4995 (
            .O(N__30276),
            .I(N__30273));
    Span12Mux_v I__4994 (
            .O(N__30273),
            .I(N__30270));
    Odrv12 I__4993 (
            .O(N__30270),
            .I(RAM_ADD_c_13));
    CEMux I__4992 (
            .O(N__30267),
            .I(N__30264));
    LocalMux I__4991 (
            .O(N__30264),
            .I(N__30259));
    CEMux I__4990 (
            .O(N__30263),
            .I(N__30256));
    CEMux I__4989 (
            .O(N__30262),
            .I(N__30253));
    Span4Mux_v I__4988 (
            .O(N__30259),
            .I(N__30248));
    LocalMux I__4987 (
            .O(N__30256),
            .I(N__30248));
    LocalMux I__4986 (
            .O(N__30253),
            .I(N__30243));
    Span4Mux_v I__4985 (
            .O(N__30248),
            .I(N__30243));
    Odrv4 I__4984 (
            .O(N__30243),
            .I(N_67_i));
    InMux I__4983 (
            .O(N__30240),
            .I(N__30237));
    LocalMux I__4982 (
            .O(N__30237),
            .I(N__30234));
    Span4Mux_v I__4981 (
            .O(N__30234),
            .I(N__30231));
    Sp12to4 I__4980 (
            .O(N__30231),
            .I(N__30228));
    Span12Mux_h I__4979 (
            .O(N__30228),
            .I(N__30225));
    Odrv12 I__4978 (
            .O(N__30225),
            .I(ADC3_c));
    IoInMux I__4977 (
            .O(N__30222),
            .I(N__30219));
    LocalMux I__4976 (
            .O(N__30219),
            .I(N__30216));
    Span4Mux_s0_v I__4975 (
            .O(N__30216),
            .I(N__30213));
    Sp12to4 I__4974 (
            .O(N__30213),
            .I(N__30210));
    Span12Mux_h I__4973 (
            .O(N__30210),
            .I(N__30207));
    Odrv12 I__4972 (
            .O(N__30207),
            .I(RAM_DATA_1Z0Z_3));
    InMux I__4971 (
            .O(N__30204),
            .I(N__30201));
    LocalMux I__4970 (
            .O(N__30201),
            .I(N__30198));
    Span4Mux_v I__4969 (
            .O(N__30198),
            .I(N__30195));
    Sp12to4 I__4968 (
            .O(N__30195),
            .I(N__30192));
    Span12Mux_h I__4967 (
            .O(N__30192),
            .I(N__30189));
    Odrv12 I__4966 (
            .O(N__30189),
            .I(ADC0_c));
    IoInMux I__4965 (
            .O(N__30186),
            .I(N__30183));
    LocalMux I__4964 (
            .O(N__30183),
            .I(N__30180));
    Span4Mux_s3_v I__4963 (
            .O(N__30180),
            .I(N__30177));
    Span4Mux_h I__4962 (
            .O(N__30177),
            .I(N__30174));
    Sp12to4 I__4961 (
            .O(N__30174),
            .I(N__30171));
    Span12Mux_s8_v I__4960 (
            .O(N__30171),
            .I(N__30168));
    Odrv12 I__4959 (
            .O(N__30168),
            .I(RAM_DATA_1Z0Z_0));
    InMux I__4958 (
            .O(N__30165),
            .I(N__30162));
    LocalMux I__4957 (
            .O(N__30162),
            .I(N__30159));
    Span4Mux_v I__4956 (
            .O(N__30159),
            .I(N__30156));
    Sp12to4 I__4955 (
            .O(N__30156),
            .I(N__30153));
    Span12Mux_h I__4954 (
            .O(N__30153),
            .I(N__30150));
    Odrv12 I__4953 (
            .O(N__30150),
            .I(ADC5_c));
    IoInMux I__4952 (
            .O(N__30147),
            .I(N__30144));
    LocalMux I__4951 (
            .O(N__30144),
            .I(N__30141));
    IoSpan4Mux I__4950 (
            .O(N__30141),
            .I(N__30138));
    Span4Mux_s2_v I__4949 (
            .O(N__30138),
            .I(N__30135));
    Sp12to4 I__4948 (
            .O(N__30135),
            .I(N__30132));
    Span12Mux_s10_v I__4947 (
            .O(N__30132),
            .I(N__30129));
    Span12Mux_h I__4946 (
            .O(N__30129),
            .I(N__30126));
    Odrv12 I__4945 (
            .O(N__30126),
            .I(RAM_DATA_1Z0Z_5));
    InMux I__4944 (
            .O(N__30123),
            .I(N__30120));
    LocalMux I__4943 (
            .O(N__30120),
            .I(N__30117));
    Span4Mux_v I__4942 (
            .O(N__30117),
            .I(N__30114));
    Sp12to4 I__4941 (
            .O(N__30114),
            .I(N__30111));
    Span12Mux_h I__4940 (
            .O(N__30111),
            .I(N__30108));
    Odrv12 I__4939 (
            .O(N__30108),
            .I(ADC1_c));
    IoInMux I__4938 (
            .O(N__30105),
            .I(N__30102));
    LocalMux I__4937 (
            .O(N__30102),
            .I(N__30099));
    Span12Mux_s9_v I__4936 (
            .O(N__30099),
            .I(N__30096));
    Span12Mux_h I__4935 (
            .O(N__30096),
            .I(N__30093));
    Odrv12 I__4934 (
            .O(N__30093),
            .I(RAM_DATA_1Z0Z_1));
    InMux I__4933 (
            .O(N__30090),
            .I(N__30087));
    LocalMux I__4932 (
            .O(N__30087),
            .I(N__30084));
    Span12Mux_s9_v I__4931 (
            .O(N__30084),
            .I(N__30081));
    Span12Mux_h I__4930 (
            .O(N__30081),
            .I(N__30078));
    Odrv12 I__4929 (
            .O(N__30078),
            .I(ADC7_c));
    IoInMux I__4928 (
            .O(N__30075),
            .I(N__30072));
    LocalMux I__4927 (
            .O(N__30072),
            .I(N__30069));
    Span4Mux_s0_h I__4926 (
            .O(N__30069),
            .I(N__30066));
    Span4Mux_v I__4925 (
            .O(N__30066),
            .I(N__30063));
    Sp12to4 I__4924 (
            .O(N__30063),
            .I(N__30060));
    Span12Mux_v I__4923 (
            .O(N__30060),
            .I(N__30057));
    Span12Mux_h I__4922 (
            .O(N__30057),
            .I(N__30054));
    Odrv12 I__4921 (
            .O(N__30054),
            .I(RAM_DATA_1Z0Z_8));
    InMux I__4920 (
            .O(N__30051),
            .I(N__30048));
    LocalMux I__4919 (
            .O(N__30048),
            .I(N__30045));
    Span4Mux_h I__4918 (
            .O(N__30045),
            .I(N__30042));
    Sp12to4 I__4917 (
            .O(N__30042),
            .I(N__30039));
    Span12Mux_v I__4916 (
            .O(N__30039),
            .I(N__30036));
    Span12Mux_h I__4915 (
            .O(N__30036),
            .I(N__30033));
    Odrv12 I__4914 (
            .O(N__30033),
            .I(RAM_DATA_in_11));
    InMux I__4913 (
            .O(N__30030),
            .I(N__30027));
    LocalMux I__4912 (
            .O(N__30027),
            .I(N__30024));
    Span4Mux_v I__4911 (
            .O(N__30024),
            .I(N__30021));
    Span4Mux_v I__4910 (
            .O(N__30021),
            .I(N__30018));
    Sp12to4 I__4909 (
            .O(N__30018),
            .I(N__30015));
    Span12Mux_h I__4908 (
            .O(N__30015),
            .I(N__30012));
    Odrv12 I__4907 (
            .O(N__30012),
            .I(RAM_DATA_in_3));
    InMux I__4906 (
            .O(N__30009),
            .I(N__30006));
    LocalMux I__4905 (
            .O(N__30006),
            .I(N__30003));
    Span4Mux_h I__4904 (
            .O(N__30003),
            .I(N__30000));
    Odrv4 I__4903 (
            .O(N__30000),
            .I(spi_data_misoZ0Z_3));
    InMux I__4902 (
            .O(N__29997),
            .I(N__29994));
    LocalMux I__4901 (
            .O(N__29994),
            .I(N__29991));
    Span4Mux_v I__4900 (
            .O(N__29991),
            .I(N__29988));
    Sp12to4 I__4899 (
            .O(N__29988),
            .I(N__29985));
    Span12Mux_v I__4898 (
            .O(N__29985),
            .I(N__29982));
    Span12Mux_h I__4897 (
            .O(N__29982),
            .I(N__29979));
    Odrv12 I__4896 (
            .O(N__29979),
            .I(RAM_DATA_in_12));
    CascadeMux I__4895 (
            .O(N__29976),
            .I(N__29973));
    InMux I__4894 (
            .O(N__29973),
            .I(N__29970));
    LocalMux I__4893 (
            .O(N__29970),
            .I(N__29967));
    Span4Mux_v I__4892 (
            .O(N__29967),
            .I(N__29964));
    Span4Mux_v I__4891 (
            .O(N__29964),
            .I(N__29961));
    Sp12to4 I__4890 (
            .O(N__29961),
            .I(N__29958));
    Span12Mux_h I__4889 (
            .O(N__29958),
            .I(N__29955));
    Odrv12 I__4888 (
            .O(N__29955),
            .I(RAM_DATA_in_4));
    InMux I__4887 (
            .O(N__29952),
            .I(N__29949));
    LocalMux I__4886 (
            .O(N__29949),
            .I(N__29946));
    Span4Mux_v I__4885 (
            .O(N__29946),
            .I(N__29943));
    Odrv4 I__4884 (
            .O(N__29943),
            .I(spi_data_misoZ0Z_4));
    CEMux I__4883 (
            .O(N__29940),
            .I(N__29934));
    InMux I__4882 (
            .O(N__29939),
            .I(N__29926));
    InMux I__4881 (
            .O(N__29938),
            .I(N__29926));
    InMux I__4880 (
            .O(N__29937),
            .I(N__29926));
    LocalMux I__4879 (
            .O(N__29934),
            .I(N__29917));
    InMux I__4878 (
            .O(N__29933),
            .I(N__29914));
    LocalMux I__4877 (
            .O(N__29926),
            .I(N__29911));
    InMux I__4876 (
            .O(N__29925),
            .I(N__29898));
    InMux I__4875 (
            .O(N__29924),
            .I(N__29898));
    InMux I__4874 (
            .O(N__29923),
            .I(N__29898));
    InMux I__4873 (
            .O(N__29922),
            .I(N__29898));
    InMux I__4872 (
            .O(N__29921),
            .I(N__29898));
    InMux I__4871 (
            .O(N__29920),
            .I(N__29898));
    Odrv4 I__4870 (
            .O(N__29917),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    LocalMux I__4869 (
            .O(N__29914),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    Odrv4 I__4868 (
            .O(N__29911),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    LocalMux I__4867 (
            .O(N__29898),
            .I(un4_sacqtime_cry_23_c_RNITTSZ0Z3));
    InMux I__4866 (
            .O(N__29889),
            .I(N__29886));
    LocalMux I__4865 (
            .O(N__29886),
            .I(N__29883));
    Span4Mux_v I__4864 (
            .O(N__29883),
            .I(N__29880));
    Sp12to4 I__4863 (
            .O(N__29880),
            .I(N__29877));
    Span12Mux_h I__4862 (
            .O(N__29877),
            .I(N__29874));
    Odrv12 I__4861 (
            .O(N__29874),
            .I(RAM_DATA_in_5));
    CascadeMux I__4860 (
            .O(N__29871),
            .I(N__29865));
    CascadeMux I__4859 (
            .O(N__29870),
            .I(N__29861));
    CascadeMux I__4858 (
            .O(N__29869),
            .I(N__29857));
    CascadeMux I__4857 (
            .O(N__29868),
            .I(N__29853));
    InMux I__4856 (
            .O(N__29865),
            .I(N__29838));
    InMux I__4855 (
            .O(N__29864),
            .I(N__29838));
    InMux I__4854 (
            .O(N__29861),
            .I(N__29838));
    InMux I__4853 (
            .O(N__29860),
            .I(N__29838));
    InMux I__4852 (
            .O(N__29857),
            .I(N__29838));
    InMux I__4851 (
            .O(N__29856),
            .I(N__29838));
    InMux I__4850 (
            .O(N__29853),
            .I(N__29833));
    InMux I__4849 (
            .O(N__29852),
            .I(N__29833));
    InMux I__4848 (
            .O(N__29851),
            .I(N__29830));
    LocalMux I__4847 (
            .O(N__29838),
            .I(N_75));
    LocalMux I__4846 (
            .O(N__29833),
            .I(N_75));
    LocalMux I__4845 (
            .O(N__29830),
            .I(N_75));
    InMux I__4844 (
            .O(N__29823),
            .I(N__29820));
    LocalMux I__4843 (
            .O(N__29820),
            .I(N__29817));
    Span4Mux_v I__4842 (
            .O(N__29817),
            .I(N__29814));
    Span4Mux_h I__4841 (
            .O(N__29814),
            .I(N__29811));
    Span4Mux_h I__4840 (
            .O(N__29811),
            .I(N__29808));
    Span4Mux_h I__4839 (
            .O(N__29808),
            .I(N__29805));
    IoSpan4Mux I__4838 (
            .O(N__29805),
            .I(N__29802));
    Odrv4 I__4837 (
            .O(N__29802),
            .I(RAM_DATA_in_13));
    InMux I__4836 (
            .O(N__29799),
            .I(N__29796));
    LocalMux I__4835 (
            .O(N__29796),
            .I(N__29793));
    Span4Mux_v I__4834 (
            .O(N__29793),
            .I(N__29790));
    Odrv4 I__4833 (
            .O(N__29790),
            .I(spi_data_misoZ0Z_5));
    CEMux I__4832 (
            .O(N__29787),
            .I(N__29784));
    LocalMux I__4831 (
            .O(N__29784),
            .I(N__29781));
    Span4Mux_v I__4830 (
            .O(N__29781),
            .I(N__29777));
    CEMux I__4829 (
            .O(N__29780),
            .I(N__29774));
    Span4Mux_h I__4828 (
            .O(N__29777),
            .I(N__29771));
    LocalMux I__4827 (
            .O(N__29774),
            .I(N__29768));
    Odrv4 I__4826 (
            .O(N__29771),
            .I(N_6));
    Odrv12 I__4825 (
            .O(N__29768),
            .I(N_6));
    InMux I__4824 (
            .O(N__29763),
            .I(N__29760));
    LocalMux I__4823 (
            .O(N__29760),
            .I(N__29757));
    Span4Mux_h I__4822 (
            .O(N__29757),
            .I(N__29754));
    Sp12to4 I__4821 (
            .O(N__29754),
            .I(N__29751));
    Span12Mux_v I__4820 (
            .O(N__29751),
            .I(N__29747));
    InMux I__4819 (
            .O(N__29750),
            .I(N__29744));
    Odrv12 I__4818 (
            .O(N__29747),
            .I(sRAM_pointer_readZ0Z_0));
    LocalMux I__4817 (
            .O(N__29744),
            .I(sRAM_pointer_readZ0Z_0));
    IoInMux I__4816 (
            .O(N__29739),
            .I(N__29736));
    LocalMux I__4815 (
            .O(N__29736),
            .I(N__29733));
    Span4Mux_s1_v I__4814 (
            .O(N__29733),
            .I(N__29730));
    Span4Mux_v I__4813 (
            .O(N__29730),
            .I(N__29727));
    Span4Mux_h I__4812 (
            .O(N__29727),
            .I(N__29724));
    Span4Mux_v I__4811 (
            .O(N__29724),
            .I(N__29721));
    Odrv4 I__4810 (
            .O(N__29721),
            .I(RAM_ADD_c_0));
    InMux I__4809 (
            .O(N__29718),
            .I(N__29715));
    LocalMux I__4808 (
            .O(N__29715),
            .I(N__29712));
    Span4Mux_h I__4807 (
            .O(N__29712),
            .I(N__29709));
    Span4Mux_v I__4806 (
            .O(N__29709),
            .I(N__29706));
    Odrv4 I__4805 (
            .O(N__29706),
            .I(reset_rpi_ibuf_RNI7JCVZ0));
    CascadeMux I__4804 (
            .O(N__29703),
            .I(N__29700));
    InMux I__4803 (
            .O(N__29700),
            .I(N__29694));
    InMux I__4802 (
            .O(N__29699),
            .I(N__29694));
    LocalMux I__4801 (
            .O(N__29694),
            .I(N__29691));
    Odrv4 I__4800 (
            .O(N__29691),
            .I(sRAM_ADD_0_sqmuxa_i_0));
    InMux I__4799 (
            .O(N__29688),
            .I(N__29685));
    LocalMux I__4798 (
            .O(N__29685),
            .I(N__29682));
    Span4Mux_v I__4797 (
            .O(N__29682),
            .I(N__29679));
    Sp12to4 I__4796 (
            .O(N__29679),
            .I(N__29676));
    Span12Mux_h I__4795 (
            .O(N__29676),
            .I(N__29672));
    InMux I__4794 (
            .O(N__29675),
            .I(N__29669));
    Odrv12 I__4793 (
            .O(N__29672),
            .I(sRAM_pointer_readZ0Z_1));
    LocalMux I__4792 (
            .O(N__29669),
            .I(sRAM_pointer_readZ0Z_1));
    IoInMux I__4791 (
            .O(N__29664),
            .I(N__29661));
    LocalMux I__4790 (
            .O(N__29661),
            .I(N__29658));
    Span4Mux_s3_v I__4789 (
            .O(N__29658),
            .I(N__29655));
    Span4Mux_h I__4788 (
            .O(N__29655),
            .I(N__29652));
    Sp12to4 I__4787 (
            .O(N__29652),
            .I(N__29649));
    Odrv12 I__4786 (
            .O(N__29649),
            .I(RAM_ADD_c_1));
    CascadeMux I__4785 (
            .O(N__29646),
            .I(N__29643));
    InMux I__4784 (
            .O(N__29643),
            .I(N__29640));
    LocalMux I__4783 (
            .O(N__29640),
            .I(N__29637));
    Span4Mux_h I__4782 (
            .O(N__29637),
            .I(N__29634));
    Span4Mux_h I__4781 (
            .O(N__29634),
            .I(N__29631));
    Span4Mux_h I__4780 (
            .O(N__29631),
            .I(N__29627));
    InMux I__4779 (
            .O(N__29630),
            .I(N__29624));
    Span4Mux_v I__4778 (
            .O(N__29627),
            .I(N__29621));
    LocalMux I__4777 (
            .O(N__29624),
            .I(sRAM_pointer_readZ0Z_10));
    Odrv4 I__4776 (
            .O(N__29621),
            .I(sRAM_pointer_readZ0Z_10));
    IoInMux I__4775 (
            .O(N__29616),
            .I(N__29613));
    LocalMux I__4774 (
            .O(N__29613),
            .I(N__29610));
    IoSpan4Mux I__4773 (
            .O(N__29610),
            .I(N__29607));
    Span4Mux_s0_h I__4772 (
            .O(N__29607),
            .I(N__29604));
    Span4Mux_v I__4771 (
            .O(N__29604),
            .I(N__29601));
    Sp12to4 I__4770 (
            .O(N__29601),
            .I(N__29598));
    Span12Mux_v I__4769 (
            .O(N__29598),
            .I(N__29595));
    Span12Mux_h I__4768 (
            .O(N__29595),
            .I(N__29592));
    Odrv12 I__4767 (
            .O(N__29592),
            .I(RAM_ADD_c_10));
    InMux I__4766 (
            .O(N__29589),
            .I(sCounterADC_cry_1));
    InMux I__4765 (
            .O(N__29586),
            .I(sCounterADC_cry_2));
    InMux I__4764 (
            .O(N__29583),
            .I(sCounterADC_cry_3));
    InMux I__4763 (
            .O(N__29580),
            .I(sCounterADC_cry_4));
    InMux I__4762 (
            .O(N__29577),
            .I(sCounterADC_cry_5));
    InMux I__4761 (
            .O(N__29574),
            .I(sCounterADC_cry_6));
    InMux I__4760 (
            .O(N__29571),
            .I(N__29568));
    LocalMux I__4759 (
            .O(N__29568),
            .I(N__29565));
    Span4Mux_h I__4758 (
            .O(N__29565),
            .I(N__29562));
    Span4Mux_v I__4757 (
            .O(N__29562),
            .I(N__29559));
    Sp12to4 I__4756 (
            .O(N__29559),
            .I(N__29556));
    Span12Mux_v I__4755 (
            .O(N__29556),
            .I(N__29553));
    Span12Mux_h I__4754 (
            .O(N__29553),
            .I(N__29550));
    Odrv12 I__4753 (
            .O(N__29550),
            .I(RAM_DATA_in_8));
    CascadeMux I__4752 (
            .O(N__29547),
            .I(N__29544));
    InMux I__4751 (
            .O(N__29544),
            .I(N__29541));
    LocalMux I__4750 (
            .O(N__29541),
            .I(N__29538));
    Span4Mux_v I__4749 (
            .O(N__29538),
            .I(N__29535));
    Sp12to4 I__4748 (
            .O(N__29535),
            .I(N__29532));
    Span12Mux_h I__4747 (
            .O(N__29532),
            .I(N__29529));
    Odrv12 I__4746 (
            .O(N__29529),
            .I(RAM_DATA_in_0));
    InMux I__4745 (
            .O(N__29526),
            .I(N__29523));
    LocalMux I__4744 (
            .O(N__29523),
            .I(N__29520));
    Sp12to4 I__4743 (
            .O(N__29520),
            .I(N__29517));
    Odrv12 I__4742 (
            .O(N__29517),
            .I(spi_data_misoZ0Z_0));
    InMux I__4741 (
            .O(N__29514),
            .I(N__29511));
    LocalMux I__4740 (
            .O(N__29511),
            .I(N__29508));
    Span12Mux_h I__4739 (
            .O(N__29508),
            .I(N__29505));
    Span12Mux_v I__4738 (
            .O(N__29505),
            .I(N__29502));
    Odrv12 I__4737 (
            .O(N__29502),
            .I(RAM_DATA_in_9));
    InMux I__4736 (
            .O(N__29499),
            .I(N__29496));
    LocalMux I__4735 (
            .O(N__29496),
            .I(N__29493));
    Sp12to4 I__4734 (
            .O(N__29493),
            .I(N__29490));
    Span12Mux_v I__4733 (
            .O(N__29490),
            .I(N__29487));
    Span12Mux_h I__4732 (
            .O(N__29487),
            .I(N__29484));
    Odrv12 I__4731 (
            .O(N__29484),
            .I(RAM_DATA_in_1));
    InMux I__4730 (
            .O(N__29481),
            .I(N__29478));
    LocalMux I__4729 (
            .O(N__29478),
            .I(N__29475));
    Span4Mux_h I__4728 (
            .O(N__29475),
            .I(N__29472));
    Odrv4 I__4727 (
            .O(N__29472),
            .I(spi_data_misoZ0Z_1));
    InMux I__4726 (
            .O(N__29469),
            .I(N__29466));
    LocalMux I__4725 (
            .O(N__29466),
            .I(N__29463));
    Span4Mux_h I__4724 (
            .O(N__29463),
            .I(N__29460));
    Span4Mux_h I__4723 (
            .O(N__29460),
            .I(N__29457));
    Sp12to4 I__4722 (
            .O(N__29457),
            .I(N__29454));
    Span12Mux_v I__4721 (
            .O(N__29454),
            .I(N__29451));
    Span12Mux_v I__4720 (
            .O(N__29451),
            .I(N__29448));
    Odrv12 I__4719 (
            .O(N__29448),
            .I(RAM_DATA_in_10));
    CascadeMux I__4718 (
            .O(N__29445),
            .I(N__29442));
    InMux I__4717 (
            .O(N__29442),
            .I(N__29439));
    LocalMux I__4716 (
            .O(N__29439),
            .I(N__29436));
    Span4Mux_v I__4715 (
            .O(N__29436),
            .I(N__29433));
    Span4Mux_v I__4714 (
            .O(N__29433),
            .I(N__29430));
    Sp12to4 I__4713 (
            .O(N__29430),
            .I(N__29427));
    Span12Mux_h I__4712 (
            .O(N__29427),
            .I(N__29424));
    Odrv12 I__4711 (
            .O(N__29424),
            .I(RAM_DATA_in_2));
    InMux I__4710 (
            .O(N__29421),
            .I(N__29418));
    LocalMux I__4709 (
            .O(N__29418),
            .I(N__29415));
    Span4Mux_h I__4708 (
            .O(N__29415),
            .I(N__29412));
    Odrv4 I__4707 (
            .O(N__29412),
            .I(spi_data_misoZ0Z_2));
    InMux I__4706 (
            .O(N__29409),
            .I(N__29406));
    LocalMux I__4705 (
            .O(N__29406),
            .I(N__29403));
    Span4Mux_h I__4704 (
            .O(N__29403),
            .I(N__29400));
    Odrv4 I__4703 (
            .O(N__29400),
            .I(sEEPoffZ0Z_11));
    InMux I__4702 (
            .O(N__29397),
            .I(N__29394));
    LocalMux I__4701 (
            .O(N__29394),
            .I(N__29391));
    Span4Mux_v I__4700 (
            .O(N__29391),
            .I(N__29388));
    Odrv4 I__4699 (
            .O(N__29388),
            .I(sEEPoffZ0Z_12));
    InMux I__4698 (
            .O(N__29385),
            .I(N__29382));
    LocalMux I__4697 (
            .O(N__29382),
            .I(N__29379));
    Odrv4 I__4696 (
            .O(N__29379),
            .I(sEEPoffZ0Z_13));
    InMux I__4695 (
            .O(N__29376),
            .I(N__29373));
    LocalMux I__4694 (
            .O(N__29373),
            .I(N__29370));
    Odrv4 I__4693 (
            .O(N__29370),
            .I(sEEPoffZ0Z_14));
    CascadeMux I__4692 (
            .O(N__29367),
            .I(N__29364));
    InMux I__4691 (
            .O(N__29364),
            .I(N__29361));
    LocalMux I__4690 (
            .O(N__29361),
            .I(N__29358));
    Odrv4 I__4689 (
            .O(N__29358),
            .I(sEEPoffZ0Z_15));
    InMux I__4688 (
            .O(N__29355),
            .I(N__29352));
    LocalMux I__4687 (
            .O(N__29352),
            .I(N__29349));
    Odrv4 I__4686 (
            .O(N__29349),
            .I(sEEPoffZ0Z_8));
    InMux I__4685 (
            .O(N__29346),
            .I(N__29343));
    LocalMux I__4684 (
            .O(N__29343),
            .I(N__29340));
    Odrv12 I__4683 (
            .O(N__29340),
            .I(sEEPoffZ0Z_9));
    CEMux I__4682 (
            .O(N__29337),
            .I(N__29334));
    LocalMux I__4681 (
            .O(N__29334),
            .I(N__29331));
    Span4Mux_v I__4680 (
            .O(N__29331),
            .I(N__29328));
    Span4Mux_h I__4679 (
            .O(N__29328),
            .I(N__29325));
    Odrv4 I__4678 (
            .O(N__29325),
            .I(sAddress_RNIA6242_1Z0Z_2));
    InMux I__4677 (
            .O(N__29322),
            .I(bfn_12_15_0_));
    InMux I__4676 (
            .O(N__29319),
            .I(sCounterADC_cry_0));
    InMux I__4675 (
            .O(N__29316),
            .I(N__29313));
    LocalMux I__4674 (
            .O(N__29313),
            .I(N__29310));
    Odrv12 I__4673 (
            .O(N__29310),
            .I(sEEPoffZ0Z_0));
    CascadeMux I__4672 (
            .O(N__29307),
            .I(N__29304));
    InMux I__4671 (
            .O(N__29304),
            .I(N__29301));
    LocalMux I__4670 (
            .O(N__29301),
            .I(N__29298));
    Span4Mux_h I__4669 (
            .O(N__29298),
            .I(N__29295));
    Odrv4 I__4668 (
            .O(N__29295),
            .I(sEEPoffZ0Z_1));
    InMux I__4667 (
            .O(N__29292),
            .I(N__29289));
    LocalMux I__4666 (
            .O(N__29289),
            .I(N__29286));
    Odrv4 I__4665 (
            .O(N__29286),
            .I(sEEPoffZ0Z_2));
    InMux I__4664 (
            .O(N__29283),
            .I(N__29280));
    LocalMux I__4663 (
            .O(N__29280),
            .I(N__29277));
    Odrv4 I__4662 (
            .O(N__29277),
            .I(sEEPoffZ0Z_3));
    InMux I__4661 (
            .O(N__29274),
            .I(N__29271));
    LocalMux I__4660 (
            .O(N__29271),
            .I(N__29268));
    Odrv4 I__4659 (
            .O(N__29268),
            .I(sEEPoffZ0Z_4));
    InMux I__4658 (
            .O(N__29265),
            .I(N__29262));
    LocalMux I__4657 (
            .O(N__29262),
            .I(N__29259));
    Odrv12 I__4656 (
            .O(N__29259),
            .I(sEEPoffZ0Z_5));
    InMux I__4655 (
            .O(N__29256),
            .I(N__29253));
    LocalMux I__4654 (
            .O(N__29253),
            .I(N__29250));
    Odrv12 I__4653 (
            .O(N__29250),
            .I(sEEPoffZ0Z_6));
    InMux I__4652 (
            .O(N__29247),
            .I(N__29244));
    LocalMux I__4651 (
            .O(N__29244),
            .I(N__29241));
    Odrv12 I__4650 (
            .O(N__29241),
            .I(sEEPoffZ0Z_7));
    InMux I__4649 (
            .O(N__29238),
            .I(N__29235));
    LocalMux I__4648 (
            .O(N__29235),
            .I(N__29232));
    Odrv12 I__4647 (
            .O(N__29232),
            .I(sEEPoffZ0Z_10));
    InMux I__4646 (
            .O(N__29229),
            .I(N__29226));
    LocalMux I__4645 (
            .O(N__29226),
            .I(N__29223));
    Odrv12 I__4644 (
            .O(N__29223),
            .I(\spi_slave_inst.un1_spointer11_2_0_a2_0_6_4 ));
    CascadeMux I__4643 (
            .O(N__29220),
            .I(\spi_slave_inst.un1_spointer11_2_0_a2_0_6_5_cascade_ ));
    InMux I__4642 (
            .O(N__29217),
            .I(N__29214));
    LocalMux I__4641 (
            .O(N__29214),
            .I(N__29210));
    InMux I__4640 (
            .O(N__29213),
            .I(N__29207));
    Span4Mux_h I__4639 (
            .O(N__29210),
            .I(N__29202));
    LocalMux I__4638 (
            .O(N__29207),
            .I(N__29202));
    Odrv4 I__4637 (
            .O(N__29202),
            .I(un1_spointer11_2_0));
    CascadeMux I__4636 (
            .O(N__29199),
            .I(N_285_cascade_));
    CascadeMux I__4635 (
            .O(N__29196),
            .I(N__29193));
    InMux I__4634 (
            .O(N__29193),
            .I(N__29185));
    InMux I__4633 (
            .O(N__29192),
            .I(N__29180));
    InMux I__4632 (
            .O(N__29191),
            .I(N__29180));
    InMux I__4631 (
            .O(N__29190),
            .I(N__29177));
    InMux I__4630 (
            .O(N__29189),
            .I(N__29173));
    InMux I__4629 (
            .O(N__29188),
            .I(N__29170));
    LocalMux I__4628 (
            .O(N__29185),
            .I(N__29167));
    LocalMux I__4627 (
            .O(N__29180),
            .I(N__29162));
    LocalMux I__4626 (
            .O(N__29177),
            .I(N__29162));
    InMux I__4625 (
            .O(N__29176),
            .I(N__29159));
    LocalMux I__4624 (
            .O(N__29173),
            .I(sPointerZ0Z_0));
    LocalMux I__4623 (
            .O(N__29170),
            .I(sPointerZ0Z_0));
    Odrv4 I__4622 (
            .O(N__29167),
            .I(sPointerZ0Z_0));
    Odrv4 I__4621 (
            .O(N__29162),
            .I(sPointerZ0Z_0));
    LocalMux I__4620 (
            .O(N__29159),
            .I(sPointerZ0Z_0));
    CascadeMux I__4619 (
            .O(N__29148),
            .I(N_116_cascade_));
    InMux I__4618 (
            .O(N__29145),
            .I(N__29141));
    InMux I__4617 (
            .O(N__29144),
            .I(N__29138));
    LocalMux I__4616 (
            .O(N__29141),
            .I(N_159));
    LocalMux I__4615 (
            .O(N__29138),
            .I(N_159));
    CascadeMux I__4614 (
            .O(N__29133),
            .I(N_117_cascade_));
    InMux I__4613 (
            .O(N__29130),
            .I(N__29124));
    InMux I__4612 (
            .O(N__29129),
            .I(N__29121));
    InMux I__4611 (
            .O(N__29128),
            .I(N__29118));
    InMux I__4610 (
            .O(N__29127),
            .I(N__29115));
    LocalMux I__4609 (
            .O(N__29124),
            .I(spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1));
    LocalMux I__4608 (
            .O(N__29121),
            .I(spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1));
    LocalMux I__4607 (
            .O(N__29118),
            .I(spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1));
    LocalMux I__4606 (
            .O(N__29115),
            .I(spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1));
    InMux I__4605 (
            .O(N__29106),
            .I(N__29090));
    InMux I__4604 (
            .O(N__29105),
            .I(N__29085));
    InMux I__4603 (
            .O(N__29104),
            .I(N__29085));
    InMux I__4602 (
            .O(N__29103),
            .I(N__29073));
    InMux I__4601 (
            .O(N__29102),
            .I(N__29073));
    InMux I__4600 (
            .O(N__29101),
            .I(N__29073));
    InMux I__4599 (
            .O(N__29100),
            .I(N__29073));
    InMux I__4598 (
            .O(N__29099),
            .I(N__29073));
    InMux I__4597 (
            .O(N__29098),
            .I(N__29064));
    InMux I__4596 (
            .O(N__29097),
            .I(N__29064));
    InMux I__4595 (
            .O(N__29096),
            .I(N__29064));
    InMux I__4594 (
            .O(N__29095),
            .I(N__29064));
    InMux I__4593 (
            .O(N__29094),
            .I(N__29061));
    InMux I__4592 (
            .O(N__29093),
            .I(N__29057));
    LocalMux I__4591 (
            .O(N__29090),
            .I(N__29054));
    LocalMux I__4590 (
            .O(N__29085),
            .I(N__29051));
    InMux I__4589 (
            .O(N__29084),
            .I(N__29048));
    LocalMux I__4588 (
            .O(N__29073),
            .I(N__29045));
    LocalMux I__4587 (
            .O(N__29064),
            .I(N__29042));
    LocalMux I__4586 (
            .O(N__29061),
            .I(N__29037));
    InMux I__4585 (
            .O(N__29060),
            .I(N__29034));
    LocalMux I__4584 (
            .O(N__29057),
            .I(N__29031));
    Span4Mux_v I__4583 (
            .O(N__29054),
            .I(N__29024));
    Span4Mux_v I__4582 (
            .O(N__29051),
            .I(N__29024));
    LocalMux I__4581 (
            .O(N__29048),
            .I(N__29024));
    Span4Mux_v I__4580 (
            .O(N__29045),
            .I(N__29019));
    Span4Mux_h I__4579 (
            .O(N__29042),
            .I(N__29019));
    InMux I__4578 (
            .O(N__29041),
            .I(N__29014));
    InMux I__4577 (
            .O(N__29040),
            .I(N__29014));
    Span12Mux_h I__4576 (
            .O(N__29037),
            .I(N__29011));
    LocalMux I__4575 (
            .O(N__29034),
            .I(N__29006));
    Span12Mux_v I__4574 (
            .O(N__29031),
            .I(N__29006));
    Span4Mux_h I__4573 (
            .O(N__29024),
            .I(N__29003));
    Span4Mux_h I__4572 (
            .O(N__29019),
            .I(N__29000));
    LocalMux I__4571 (
            .O(N__29014),
            .I(sEETrigInternalZ0));
    Odrv12 I__4570 (
            .O(N__29011),
            .I(sEETrigInternalZ0));
    Odrv12 I__4569 (
            .O(N__29006),
            .I(sEETrigInternalZ0));
    Odrv4 I__4568 (
            .O(N__29003),
            .I(sEETrigInternalZ0));
    Odrv4 I__4567 (
            .O(N__29000),
            .I(sEETrigInternalZ0));
    CEMux I__4566 (
            .O(N__28989),
            .I(N__28985));
    CEMux I__4565 (
            .O(N__28988),
            .I(N__28982));
    LocalMux I__4564 (
            .O(N__28985),
            .I(N__28977));
    LocalMux I__4563 (
            .O(N__28982),
            .I(N__28977));
    Sp12to4 I__4562 (
            .O(N__28977),
            .I(N__28974));
    Odrv12 I__4561 (
            .O(N__28974),
            .I(sDAC_mem_23_1_sqmuxa));
    CascadeMux I__4560 (
            .O(N__28971),
            .I(N_275_cascade_));
    CascadeMux I__4559 (
            .O(N__28968),
            .I(N_360_cascade_));
    InMux I__4558 (
            .O(N__28965),
            .I(N__28962));
    LocalMux I__4557 (
            .O(N__28962),
            .I(N_269));
    InMux I__4556 (
            .O(N__28959),
            .I(N__28956));
    LocalMux I__4555 (
            .O(N__28956),
            .I(N__28953));
    Span4Mux_h I__4554 (
            .O(N__28953),
            .I(N__28950));
    Span4Mux_h I__4553 (
            .O(N__28950),
            .I(N__28947));
    Odrv4 I__4552 (
            .O(N__28947),
            .I(N_132));
    CEMux I__4551 (
            .O(N__28944),
            .I(N__28941));
    LocalMux I__4550 (
            .O(N__28941),
            .I(N__28938));
    Odrv12 I__4549 (
            .O(N__28938),
            .I(sAddress_RNIA6242_0Z0Z_0));
    CascadeMux I__4548 (
            .O(N__28935),
            .I(N__28932));
    InMux I__4547 (
            .O(N__28932),
            .I(N__28929));
    LocalMux I__4546 (
            .O(N__28929),
            .I(un1_spointer11_7_0_tz));
    CascadeMux I__4545 (
            .O(N__28926),
            .I(un1_spointer11_7_0_tz_cascade_));
    CEMux I__4544 (
            .O(N__28923),
            .I(N__28920));
    LocalMux I__4543 (
            .O(N__28920),
            .I(N__28917));
    Odrv12 I__4542 (
            .O(N__28917),
            .I(sAddress_RNID9242Z0Z_3));
    CascadeMux I__4541 (
            .O(N__28914),
            .I(un1_spointer11_5_0_2_cascade_));
    CEMux I__4540 (
            .O(N__28911),
            .I(N__28908));
    LocalMux I__4539 (
            .O(N__28908),
            .I(N__28905));
    Span4Mux_v I__4538 (
            .O(N__28905),
            .I(N__28902));
    Odrv4 I__4537 (
            .O(N__28902),
            .I(sAddress_RNIA6242_0Z0Z_2));
    InMux I__4536 (
            .O(N__28899),
            .I(N__28896));
    LocalMux I__4535 (
            .O(N__28896),
            .I(N__28893));
    Odrv4 I__4534 (
            .O(N__28893),
            .I(sDAC_dataZ0Z_0));
    InMux I__4533 (
            .O(N__28890),
            .I(N__28887));
    LocalMux I__4532 (
            .O(N__28887),
            .I(N__28884));
    Span4Mux_h I__4531 (
            .O(N__28884),
            .I(N__28881));
    Odrv4 I__4530 (
            .O(N__28881),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_0 ));
    InMux I__4529 (
            .O(N__28878),
            .I(N__28875));
    LocalMux I__4528 (
            .O(N__28875),
            .I(N__28872));
    Span4Mux_h I__4527 (
            .O(N__28872),
            .I(N__28869));
    Odrv4 I__4526 (
            .O(N__28869),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_7 ));
    InMux I__4525 (
            .O(N__28866),
            .I(N__28863));
    LocalMux I__4524 (
            .O(N__28863),
            .I(N__28860));
    Span4Mux_h I__4523 (
            .O(N__28860),
            .I(N__28857));
    Odrv4 I__4522 (
            .O(N__28857),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_8 ));
    InMux I__4521 (
            .O(N__28854),
            .I(N__28851));
    LocalMux I__4520 (
            .O(N__28851),
            .I(N__28848));
    Span4Mux_v I__4519 (
            .O(N__28848),
            .I(N__28845));
    Odrv4 I__4518 (
            .O(N__28845),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_9 ));
    CEMux I__4517 (
            .O(N__28842),
            .I(N__28838));
    CEMux I__4516 (
            .O(N__28841),
            .I(N__28834));
    LocalMux I__4515 (
            .O(N__28838),
            .I(N__28831));
    CascadeMux I__4514 (
            .O(N__28837),
            .I(N__28828));
    LocalMux I__4513 (
            .O(N__28834),
            .I(N__28825));
    Span4Mux_v I__4512 (
            .O(N__28831),
            .I(N__28822));
    InMux I__4511 (
            .O(N__28828),
            .I(N__28819));
    Odrv12 I__4510 (
            .O(N__28825),
            .I(\spi_master_inst.spi_data_path_u1.tx_ready_iZ0 ));
    Odrv4 I__4509 (
            .O(N__28822),
            .I(\spi_master_inst.spi_data_path_u1.tx_ready_iZ0 ));
    LocalMux I__4508 (
            .O(N__28819),
            .I(\spi_master_inst.spi_data_path_u1.tx_ready_iZ0 ));
    InMux I__4507 (
            .O(N__28812),
            .I(N__28809));
    LocalMux I__4506 (
            .O(N__28809),
            .I(N__28806));
    Span4Mux_h I__4505 (
            .O(N__28806),
            .I(N__28802));
    InMux I__4504 (
            .O(N__28805),
            .I(N__28799));
    Odrv4 I__4503 (
            .O(N__28802),
            .I(\spi_slave_inst.rx_done_reg1_iZ0 ));
    LocalMux I__4502 (
            .O(N__28799),
            .I(\spi_slave_inst.rx_done_reg1_iZ0 ));
    InMux I__4501 (
            .O(N__28794),
            .I(N__28789));
    InMux I__4500 (
            .O(N__28793),
            .I(N__28784));
    InMux I__4499 (
            .O(N__28792),
            .I(N__28784));
    LocalMux I__4498 (
            .O(N__28789),
            .I(N__28781));
    LocalMux I__4497 (
            .O(N__28784),
            .I(N__28778));
    Span4Mux_h I__4496 (
            .O(N__28781),
            .I(N__28775));
    Span12Mux_v I__4495 (
            .O(N__28778),
            .I(N__28772));
    Odrv4 I__4494 (
            .O(N__28775),
            .I(\spi_slave_inst.rx_done_reg2_iZ0 ));
    Odrv12 I__4493 (
            .O(N__28772),
            .I(\spi_slave_inst.rx_done_reg2_iZ0 ));
    CEMux I__4492 (
            .O(N__28767),
            .I(N__28764));
    LocalMux I__4491 (
            .O(N__28764),
            .I(\spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541 ));
    InMux I__4490 (
            .O(N__28761),
            .I(N__28758));
    LocalMux I__4489 (
            .O(N__28758),
            .I(N__28755));
    Odrv12 I__4488 (
            .O(N__28755),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_10 ));
    InMux I__4487 (
            .O(N__28752),
            .I(N__28749));
    LocalMux I__4486 (
            .O(N__28749),
            .I(N__28746));
    Span4Mux_v I__4485 (
            .O(N__28746),
            .I(N__28743));
    Span4Mux_h I__4484 (
            .O(N__28743),
            .I(N__28740));
    Odrv4 I__4483 (
            .O(N__28740),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_13 ));
    InMux I__4482 (
            .O(N__28737),
            .I(N__28734));
    LocalMux I__4481 (
            .O(N__28734),
            .I(N__28731));
    Odrv4 I__4480 (
            .O(N__28731),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_4 ));
    InMux I__4479 (
            .O(N__28728),
            .I(N__28725));
    LocalMux I__4478 (
            .O(N__28725),
            .I(N__28722));
    Odrv12 I__4477 (
            .O(N__28722),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_5 ));
    InMux I__4476 (
            .O(N__28719),
            .I(N__28716));
    LocalMux I__4475 (
            .O(N__28716),
            .I(N__28713));
    Sp12to4 I__4474 (
            .O(N__28713),
            .I(N__28710));
    Span12Mux_v I__4473 (
            .O(N__28710),
            .I(N__28707));
    Span12Mux_h I__4472 (
            .O(N__28707),
            .I(N__28704));
    Odrv12 I__4471 (
            .O(N__28704),
            .I(spi_sclk_ft_c));
    IoInMux I__4470 (
            .O(N__28701),
            .I(N__28698));
    LocalMux I__4469 (
            .O(N__28698),
            .I(N__28695));
    Span4Mux_s3_v I__4468 (
            .O(N__28695),
            .I(N__28692));
    Odrv4 I__4467 (
            .O(N__28692),
            .I(spi_sclk));
    CascadeMux I__4466 (
            .O(N__28689),
            .I(N__28686));
    InMux I__4465 (
            .O(N__28686),
            .I(N__28683));
    LocalMux I__4464 (
            .O(N__28683),
            .I(N__28680));
    Span4Mux_v I__4463 (
            .O(N__28680),
            .I(N__28677));
    Span4Mux_h I__4462 (
            .O(N__28677),
            .I(N__28674));
    Span4Mux_h I__4461 (
            .O(N__28674),
            .I(N__28670));
    InMux I__4460 (
            .O(N__28673),
            .I(N__28667));
    Odrv4 I__4459 (
            .O(N__28670),
            .I(sRAM_pointer_readZ0Z_3));
    LocalMux I__4458 (
            .O(N__28667),
            .I(sRAM_pointer_readZ0Z_3));
    IoInMux I__4457 (
            .O(N__28662),
            .I(N__28659));
    LocalMux I__4456 (
            .O(N__28659),
            .I(N__28656));
    Span12Mux_s9_v I__4455 (
            .O(N__28656),
            .I(N__28653));
    Odrv12 I__4454 (
            .O(N__28653),
            .I(RAM_ADD_c_3));
    InMux I__4453 (
            .O(N__28650),
            .I(N__28647));
    LocalMux I__4452 (
            .O(N__28647),
            .I(N__28644));
    Span4Mux_v I__4451 (
            .O(N__28644),
            .I(N__28641));
    Span4Mux_h I__4450 (
            .O(N__28641),
            .I(N__28638));
    Span4Mux_h I__4449 (
            .O(N__28638),
            .I(N__28634));
    InMux I__4448 (
            .O(N__28637),
            .I(N__28631));
    Odrv4 I__4447 (
            .O(N__28634),
            .I(sRAM_pointer_readZ0Z_4));
    LocalMux I__4446 (
            .O(N__28631),
            .I(sRAM_pointer_readZ0Z_4));
    IoInMux I__4445 (
            .O(N__28626),
            .I(N__28623));
    LocalMux I__4444 (
            .O(N__28623),
            .I(N__28620));
    Span4Mux_s1_v I__4443 (
            .O(N__28620),
            .I(N__28617));
    Span4Mux_v I__4442 (
            .O(N__28617),
            .I(N__28614));
    Span4Mux_v I__4441 (
            .O(N__28614),
            .I(N__28611));
    Sp12to4 I__4440 (
            .O(N__28611),
            .I(N__28608));
    Odrv12 I__4439 (
            .O(N__28608),
            .I(RAM_ADD_c_4));
    InMux I__4438 (
            .O(N__28605),
            .I(N__28602));
    LocalMux I__4437 (
            .O(N__28602),
            .I(N__28599));
    Span4Mux_v I__4436 (
            .O(N__28599),
            .I(N__28596));
    Span4Mux_h I__4435 (
            .O(N__28596),
            .I(N__28593));
    Span4Mux_h I__4434 (
            .O(N__28593),
            .I(N__28589));
    InMux I__4433 (
            .O(N__28592),
            .I(N__28586));
    Odrv4 I__4432 (
            .O(N__28589),
            .I(sRAM_pointer_readZ0Z_5));
    LocalMux I__4431 (
            .O(N__28586),
            .I(sRAM_pointer_readZ0Z_5));
    IoInMux I__4430 (
            .O(N__28581),
            .I(N__28578));
    LocalMux I__4429 (
            .O(N__28578),
            .I(N__28575));
    Span4Mux_s2_h I__4428 (
            .O(N__28575),
            .I(N__28572));
    Span4Mux_v I__4427 (
            .O(N__28572),
            .I(N__28569));
    Sp12to4 I__4426 (
            .O(N__28569),
            .I(N__28566));
    Span12Mux_s9_h I__4425 (
            .O(N__28566),
            .I(N__28563));
    Odrv12 I__4424 (
            .O(N__28563),
            .I(RAM_ADD_c_5));
    InMux I__4423 (
            .O(N__28560),
            .I(N__28557));
    LocalMux I__4422 (
            .O(N__28557),
            .I(N__28554));
    Span4Mux_v I__4421 (
            .O(N__28554),
            .I(N__28551));
    Span4Mux_h I__4420 (
            .O(N__28551),
            .I(N__28548));
    Span4Mux_h I__4419 (
            .O(N__28548),
            .I(N__28544));
    InMux I__4418 (
            .O(N__28547),
            .I(N__28541));
    Odrv4 I__4417 (
            .O(N__28544),
            .I(sRAM_pointer_readZ0Z_6));
    LocalMux I__4416 (
            .O(N__28541),
            .I(sRAM_pointer_readZ0Z_6));
    IoInMux I__4415 (
            .O(N__28536),
            .I(N__28533));
    LocalMux I__4414 (
            .O(N__28533),
            .I(N__28530));
    Span4Mux_s2_h I__4413 (
            .O(N__28530),
            .I(N__28527));
    Span4Mux_h I__4412 (
            .O(N__28527),
            .I(N__28524));
    Span4Mux_h I__4411 (
            .O(N__28524),
            .I(N__28521));
    Sp12to4 I__4410 (
            .O(N__28521),
            .I(N__28518));
    Span12Mux_s8_v I__4409 (
            .O(N__28518),
            .I(N__28515));
    Odrv12 I__4408 (
            .O(N__28515),
            .I(RAM_ADD_c_6));
    CascadeMux I__4407 (
            .O(N__28512),
            .I(N__28509));
    InMux I__4406 (
            .O(N__28509),
            .I(N__28506));
    LocalMux I__4405 (
            .O(N__28506),
            .I(N__28503));
    Sp12to4 I__4404 (
            .O(N__28503),
            .I(N__28500));
    Span12Mux_v I__4403 (
            .O(N__28500),
            .I(N__28496));
    InMux I__4402 (
            .O(N__28499),
            .I(N__28493));
    Odrv12 I__4401 (
            .O(N__28496),
            .I(sRAM_pointer_readZ0Z_7));
    LocalMux I__4400 (
            .O(N__28493),
            .I(sRAM_pointer_readZ0Z_7));
    IoInMux I__4399 (
            .O(N__28488),
            .I(N__28485));
    LocalMux I__4398 (
            .O(N__28485),
            .I(N__28482));
    Span4Mux_s3_h I__4397 (
            .O(N__28482),
            .I(N__28479));
    Span4Mux_h I__4396 (
            .O(N__28479),
            .I(N__28476));
    Span4Mux_h I__4395 (
            .O(N__28476),
            .I(N__28473));
    Sp12to4 I__4394 (
            .O(N__28473),
            .I(N__28470));
    Span12Mux_s8_v I__4393 (
            .O(N__28470),
            .I(N__28467));
    Odrv12 I__4392 (
            .O(N__28467),
            .I(RAM_ADD_c_7));
    InMux I__4391 (
            .O(N__28464),
            .I(N__28461));
    LocalMux I__4390 (
            .O(N__28461),
            .I(N__28458));
    Span4Mux_v I__4389 (
            .O(N__28458),
            .I(N__28455));
    Span4Mux_h I__4388 (
            .O(N__28455),
            .I(N__28452));
    Span4Mux_h I__4387 (
            .O(N__28452),
            .I(N__28448));
    InMux I__4386 (
            .O(N__28451),
            .I(N__28445));
    Odrv4 I__4385 (
            .O(N__28448),
            .I(sRAM_pointer_readZ0Z_8));
    LocalMux I__4384 (
            .O(N__28445),
            .I(sRAM_pointer_readZ0Z_8));
    IoInMux I__4383 (
            .O(N__28440),
            .I(N__28437));
    LocalMux I__4382 (
            .O(N__28437),
            .I(N__28434));
    IoSpan4Mux I__4381 (
            .O(N__28434),
            .I(N__28431));
    Span4Mux_s3_h I__4380 (
            .O(N__28431),
            .I(N__28428));
    Sp12to4 I__4379 (
            .O(N__28428),
            .I(N__28425));
    Span12Mux_h I__4378 (
            .O(N__28425),
            .I(N__28422));
    Odrv12 I__4377 (
            .O(N__28422),
            .I(RAM_ADD_c_8));
    CascadeMux I__4376 (
            .O(N__28419),
            .I(N__28416));
    InMux I__4375 (
            .O(N__28416),
            .I(N__28413));
    LocalMux I__4374 (
            .O(N__28413),
            .I(N__28410));
    Span4Mux_v I__4373 (
            .O(N__28410),
            .I(N__28407));
    Sp12to4 I__4372 (
            .O(N__28407),
            .I(N__28404));
    Span12Mux_h I__4371 (
            .O(N__28404),
            .I(N__28400));
    InMux I__4370 (
            .O(N__28403),
            .I(N__28397));
    Odrv12 I__4369 (
            .O(N__28400),
            .I(sRAM_pointer_readZ0Z_9));
    LocalMux I__4368 (
            .O(N__28397),
            .I(sRAM_pointer_readZ0Z_9));
    IoInMux I__4367 (
            .O(N__28392),
            .I(N__28389));
    LocalMux I__4366 (
            .O(N__28389),
            .I(N__28386));
    IoSpan4Mux I__4365 (
            .O(N__28386),
            .I(N__28383));
    IoSpan4Mux I__4364 (
            .O(N__28383),
            .I(N__28380));
    Sp12to4 I__4363 (
            .O(N__28380),
            .I(N__28377));
    Span12Mux_s7_h I__4362 (
            .O(N__28377),
            .I(N__28374));
    Odrv12 I__4361 (
            .O(N__28374),
            .I(RAM_ADD_c_9));
    InMux I__4360 (
            .O(N__28371),
            .I(N__28368));
    LocalMux I__4359 (
            .O(N__28368),
            .I(N__28365));
    Odrv4 I__4358 (
            .O(N__28365),
            .I(N_102));
    IoInMux I__4357 (
            .O(N__28362),
            .I(N__28359));
    LocalMux I__4356 (
            .O(N__28359),
            .I(N__28356));
    IoSpan4Mux I__4355 (
            .O(N__28356),
            .I(N__28353));
    Sp12to4 I__4354 (
            .O(N__28353),
            .I(N__28349));
    InMux I__4353 (
            .O(N__28352),
            .I(N__28346));
    Span12Mux_s7_h I__4352 (
            .O(N__28349),
            .I(N__28343));
    LocalMux I__4351 (
            .O(N__28346),
            .I(N__28340));
    Span12Mux_v I__4350 (
            .O(N__28343),
            .I(N__28337));
    Span4Mux_h I__4349 (
            .O(N__28340),
            .I(N__28334));
    Odrv12 I__4348 (
            .O(N__28337),
            .I(RAM_DATA_cl_15Z0Z_15));
    Odrv4 I__4347 (
            .O(N__28334),
            .I(RAM_DATA_cl_15Z0Z_15));
    CascadeMux I__4346 (
            .O(N__28329),
            .I(N_96_cascade_));
    IoInMux I__4345 (
            .O(N__28326),
            .I(N__28323));
    LocalMux I__4344 (
            .O(N__28323),
            .I(N__28320));
    IoSpan4Mux I__4343 (
            .O(N__28320),
            .I(N__28317));
    Span4Mux_s2_v I__4342 (
            .O(N__28317),
            .I(N__28314));
    Sp12to4 I__4341 (
            .O(N__28314),
            .I(N__28311));
    Span12Mux_s10_v I__4340 (
            .O(N__28311),
            .I(N__28307));
    InMux I__4339 (
            .O(N__28310),
            .I(N__28304));
    Odrv12 I__4338 (
            .O(N__28307),
            .I(RAM_DATA_cl_8Z0Z_15));
    LocalMux I__4337 (
            .O(N__28304),
            .I(RAM_DATA_cl_8Z0Z_15));
    CascadeMux I__4336 (
            .O(N__28299),
            .I(N__28296));
    InMux I__4335 (
            .O(N__28296),
            .I(N__28293));
    LocalMux I__4334 (
            .O(N__28293),
            .I(N__28290));
    Sp12to4 I__4333 (
            .O(N__28290),
            .I(N__28286));
    InMux I__4332 (
            .O(N__28289),
            .I(N__28283));
    Span12Mux_v I__4331 (
            .O(N__28286),
            .I(N__28280));
    LocalMux I__4330 (
            .O(N__28283),
            .I(sRAM_pointer_readZ0Z_14));
    Odrv12 I__4329 (
            .O(N__28280),
            .I(sRAM_pointer_readZ0Z_14));
    IoInMux I__4328 (
            .O(N__28275),
            .I(N__28272));
    LocalMux I__4327 (
            .O(N__28272),
            .I(N__28269));
    IoSpan4Mux I__4326 (
            .O(N__28269),
            .I(N__28266));
    Span4Mux_s1_h I__4325 (
            .O(N__28266),
            .I(N__28263));
    Span4Mux_h I__4324 (
            .O(N__28263),
            .I(N__28260));
    Sp12to4 I__4323 (
            .O(N__28260),
            .I(N__28257));
    Span12Mux_v I__4322 (
            .O(N__28257),
            .I(N__28254));
    Span12Mux_h I__4321 (
            .O(N__28254),
            .I(N__28251));
    Odrv12 I__4320 (
            .O(N__28251),
            .I(RAM_ADD_c_14));
    InMux I__4319 (
            .O(N__28248),
            .I(N__28245));
    LocalMux I__4318 (
            .O(N__28245),
            .I(N__28242));
    Span12Mux_v I__4317 (
            .O(N__28242),
            .I(N__28238));
    InMux I__4316 (
            .O(N__28241),
            .I(N__28235));
    Odrv12 I__4315 (
            .O(N__28238),
            .I(sRAM_pointer_readZ0Z_15));
    LocalMux I__4314 (
            .O(N__28235),
            .I(sRAM_pointer_readZ0Z_15));
    IoInMux I__4313 (
            .O(N__28230),
            .I(N__28227));
    LocalMux I__4312 (
            .O(N__28227),
            .I(N__28224));
    IoSpan4Mux I__4311 (
            .O(N__28224),
            .I(N__28221));
    Span4Mux_s2_h I__4310 (
            .O(N__28221),
            .I(N__28218));
    Sp12to4 I__4309 (
            .O(N__28218),
            .I(N__28215));
    Span12Mux_s10_h I__4308 (
            .O(N__28215),
            .I(N__28212));
    Odrv12 I__4307 (
            .O(N__28212),
            .I(RAM_ADD_c_15));
    InMux I__4306 (
            .O(N__28209),
            .I(N__28206));
    LocalMux I__4305 (
            .O(N__28206),
            .I(N__28203));
    Span4Mux_h I__4304 (
            .O(N__28203),
            .I(N__28200));
    Span4Mux_h I__4303 (
            .O(N__28200),
            .I(N__28196));
    InMux I__4302 (
            .O(N__28199),
            .I(N__28193));
    Span4Mux_v I__4301 (
            .O(N__28196),
            .I(N__28190));
    LocalMux I__4300 (
            .O(N__28193),
            .I(sRAM_pointer_readZ0Z_16));
    Odrv4 I__4299 (
            .O(N__28190),
            .I(sRAM_pointer_readZ0Z_16));
    IoInMux I__4298 (
            .O(N__28185),
            .I(N__28182));
    LocalMux I__4297 (
            .O(N__28182),
            .I(N__28179));
    Span12Mux_s5_h I__4296 (
            .O(N__28179),
            .I(N__28176));
    Span12Mux_v I__4295 (
            .O(N__28176),
            .I(N__28173));
    Span12Mux_h I__4294 (
            .O(N__28173),
            .I(N__28170));
    Span12Mux_v I__4293 (
            .O(N__28170),
            .I(N__28167));
    Odrv12 I__4292 (
            .O(N__28167),
            .I(RAM_ADD_c_16));
    InMux I__4291 (
            .O(N__28164),
            .I(N__28161));
    LocalMux I__4290 (
            .O(N__28161),
            .I(N__28158));
    Span4Mux_h I__4289 (
            .O(N__28158),
            .I(N__28155));
    Span4Mux_h I__4288 (
            .O(N__28155),
            .I(N__28152));
    Span4Mux_v I__4287 (
            .O(N__28152),
            .I(N__28148));
    InMux I__4286 (
            .O(N__28151),
            .I(N__28145));
    Odrv4 I__4285 (
            .O(N__28148),
            .I(sRAM_pointer_readZ0Z_17));
    LocalMux I__4284 (
            .O(N__28145),
            .I(sRAM_pointer_readZ0Z_17));
    IoInMux I__4283 (
            .O(N__28140),
            .I(N__28137));
    LocalMux I__4282 (
            .O(N__28137),
            .I(N__28134));
    Sp12to4 I__4281 (
            .O(N__28134),
            .I(N__28131));
    Span12Mux_h I__4280 (
            .O(N__28131),
            .I(N__28128));
    Odrv12 I__4279 (
            .O(N__28128),
            .I(RAM_ADD_c_17));
    CascadeMux I__4278 (
            .O(N__28125),
            .I(N__28122));
    InMux I__4277 (
            .O(N__28122),
            .I(N__28119));
    LocalMux I__4276 (
            .O(N__28119),
            .I(N__28116));
    Span4Mux_v I__4275 (
            .O(N__28116),
            .I(N__28113));
    Span4Mux_h I__4274 (
            .O(N__28113),
            .I(N__28110));
    Span4Mux_h I__4273 (
            .O(N__28110),
            .I(N__28106));
    InMux I__4272 (
            .O(N__28109),
            .I(N__28103));
    Odrv4 I__4271 (
            .O(N__28106),
            .I(sRAM_pointer_readZ0Z_18));
    LocalMux I__4270 (
            .O(N__28103),
            .I(sRAM_pointer_readZ0Z_18));
    IoInMux I__4269 (
            .O(N__28098),
            .I(N__28095));
    LocalMux I__4268 (
            .O(N__28095),
            .I(N__28092));
    Span12Mux_s5_h I__4267 (
            .O(N__28092),
            .I(N__28089));
    Span12Mux_h I__4266 (
            .O(N__28089),
            .I(N__28086));
    Span12Mux_v I__4265 (
            .O(N__28086),
            .I(N__28083));
    Odrv12 I__4264 (
            .O(N__28083),
            .I(RAM_ADD_c_18));
    InMux I__4263 (
            .O(N__28080),
            .I(N__28077));
    LocalMux I__4262 (
            .O(N__28077),
            .I(N__28074));
    Span4Mux_v I__4261 (
            .O(N__28074),
            .I(N__28071));
    Span4Mux_h I__4260 (
            .O(N__28071),
            .I(N__28068));
    Span4Mux_h I__4259 (
            .O(N__28068),
            .I(N__28064));
    InMux I__4258 (
            .O(N__28067),
            .I(N__28061));
    Odrv4 I__4257 (
            .O(N__28064),
            .I(sRAM_pointer_readZ0Z_2));
    LocalMux I__4256 (
            .O(N__28061),
            .I(sRAM_pointer_readZ0Z_2));
    IoInMux I__4255 (
            .O(N__28056),
            .I(N__28053));
    LocalMux I__4254 (
            .O(N__28053),
            .I(N__28050));
    Span4Mux_s2_v I__4253 (
            .O(N__28050),
            .I(N__28047));
    Span4Mux_h I__4252 (
            .O(N__28047),
            .I(N__28044));
    Span4Mux_v I__4251 (
            .O(N__28044),
            .I(N__28041));
    Odrv4 I__4250 (
            .O(N__28041),
            .I(RAM_ADD_c_2));
    InMux I__4249 (
            .O(N__28038),
            .I(N__28035));
    LocalMux I__4248 (
            .O(N__28035),
            .I(N__28031));
    InMux I__4247 (
            .O(N__28034),
            .I(N__28028));
    Span4Mux_h I__4246 (
            .O(N__28031),
            .I(N__28025));
    LocalMux I__4245 (
            .O(N__28028),
            .I(sCounterRAMZ0Z_2));
    Odrv4 I__4244 (
            .O(N__28025),
            .I(sCounterRAMZ0Z_2));
    InMux I__4243 (
            .O(N__28020),
            .I(N__28017));
    LocalMux I__4242 (
            .O(N__28017),
            .I(N__28014));
    Span4Mux_v I__4241 (
            .O(N__28014),
            .I(N__28010));
    InMux I__4240 (
            .O(N__28013),
            .I(N__28007));
    Span4Mux_h I__4239 (
            .O(N__28010),
            .I(N__28004));
    LocalMux I__4238 (
            .O(N__28007),
            .I(sCounterRAMZ0Z_1));
    Odrv4 I__4237 (
            .O(N__28004),
            .I(sCounterRAMZ0Z_1));
    CascadeMux I__4236 (
            .O(N__27999),
            .I(spi_data_miso_0_sqmuxa_2_i_o2_5_cascade_));
    InMux I__4235 (
            .O(N__27996),
            .I(N__27993));
    LocalMux I__4234 (
            .O(N__27993),
            .I(N__27990));
    Span4Mux_v I__4233 (
            .O(N__27990),
            .I(N__27987));
    Odrv4 I__4232 (
            .O(N__27987),
            .I(spi_data_miso_0_sqmuxa_2_i_o2_4));
    CascadeMux I__4231 (
            .O(N__27984),
            .I(N_75_cascade_));
    InMux I__4230 (
            .O(N__27981),
            .I(N__27975));
    CascadeMux I__4229 (
            .O(N__27980),
            .I(N__27972));
    InMux I__4228 (
            .O(N__27979),
            .I(N__27969));
    InMux I__4227 (
            .O(N__27978),
            .I(N__27966));
    LocalMux I__4226 (
            .O(N__27975),
            .I(N__27963));
    InMux I__4225 (
            .O(N__27972),
            .I(N__27960));
    LocalMux I__4224 (
            .O(N__27969),
            .I(N__27957));
    LocalMux I__4223 (
            .O(N__27966),
            .I(N__27953));
    Span4Mux_h I__4222 (
            .O(N__27963),
            .I(N__27948));
    LocalMux I__4221 (
            .O(N__27960),
            .I(N__27948));
    Span4Mux_h I__4220 (
            .O(N__27957),
            .I(N__27945));
    CascadeMux I__4219 (
            .O(N__27956),
            .I(N__27942));
    Span4Mux_h I__4218 (
            .O(N__27953),
            .I(N__27939));
    Span4Mux_v I__4217 (
            .O(N__27948),
            .I(N__27936));
    Span4Mux_h I__4216 (
            .O(N__27945),
            .I(N__27933));
    InMux I__4215 (
            .O(N__27942),
            .I(N__27930));
    Span4Mux_h I__4214 (
            .O(N__27939),
            .I(N__27927));
    Span4Mux_v I__4213 (
            .O(N__27936),
            .I(N__27924));
    Span4Mux_v I__4212 (
            .O(N__27933),
            .I(N__27921));
    LocalMux I__4211 (
            .O(N__27930),
            .I(sSPI_MSB0LSBZ0Z1));
    Odrv4 I__4210 (
            .O(N__27927),
            .I(sSPI_MSB0LSBZ0Z1));
    Odrv4 I__4209 (
            .O(N__27924),
            .I(sSPI_MSB0LSBZ0Z1));
    Odrv4 I__4208 (
            .O(N__27921),
            .I(sSPI_MSB0LSBZ0Z1));
    CascadeMux I__4207 (
            .O(N__27912),
            .I(N__27908));
    InMux I__4206 (
            .O(N__27911),
            .I(N__27904));
    InMux I__4205 (
            .O(N__27908),
            .I(N__27901));
    InMux I__4204 (
            .O(N__27907),
            .I(N__27898));
    LocalMux I__4203 (
            .O(N__27904),
            .I(N__27894));
    LocalMux I__4202 (
            .O(N__27901),
            .I(N__27889));
    LocalMux I__4201 (
            .O(N__27898),
            .I(N__27889));
    InMux I__4200 (
            .O(N__27897),
            .I(N__27886));
    Span4Mux_h I__4199 (
            .O(N__27894),
            .I(N__27883));
    Span4Mux_v I__4198 (
            .O(N__27889),
            .I(N__27879));
    LocalMux I__4197 (
            .O(N__27886),
            .I(N__27876));
    Span4Mux_h I__4196 (
            .O(N__27883),
            .I(N__27873));
    InMux I__4195 (
            .O(N__27882),
            .I(N__27870));
    Span4Mux_h I__4194 (
            .O(N__27879),
            .I(N__27865));
    Span4Mux_v I__4193 (
            .O(N__27876),
            .I(N__27865));
    Odrv4 I__4192 (
            .O(N__27873),
            .I(spi_mosi_ready_prev3_RNILKERZ0));
    LocalMux I__4191 (
            .O(N__27870),
            .I(spi_mosi_ready_prev3_RNILKERZ0));
    Odrv4 I__4190 (
            .O(N__27865),
            .I(spi_mosi_ready_prev3_RNILKERZ0));
    InMux I__4189 (
            .O(N__27858),
            .I(N__27855));
    LocalMux I__4188 (
            .O(N__27855),
            .I(N_88));
    CascadeMux I__4187 (
            .O(N__27852),
            .I(N_88_cascade_));
    IoInMux I__4186 (
            .O(N__27849),
            .I(N__27846));
    LocalMux I__4185 (
            .O(N__27846),
            .I(N__27843));
    Span4Mux_s1_h I__4184 (
            .O(N__27843),
            .I(N__27840));
    Span4Mux_h I__4183 (
            .O(N__27840),
            .I(N__27837));
    Span4Mux_h I__4182 (
            .O(N__27837),
            .I(N__27834));
    Span4Mux_h I__4181 (
            .O(N__27834),
            .I(N__27831));
    Span4Mux_v I__4180 (
            .O(N__27831),
            .I(N__27828));
    Odrv4 I__4179 (
            .O(N__27828),
            .I(N_28));
    CascadeMux I__4178 (
            .O(N__27825),
            .I(N_93_cascade_));
    IoInMux I__4177 (
            .O(N__27822),
            .I(N__27819));
    LocalMux I__4176 (
            .O(N__27819),
            .I(N__27816));
    Span4Mux_s0_v I__4175 (
            .O(N__27816),
            .I(N__27813));
    Span4Mux_h I__4174 (
            .O(N__27813),
            .I(N__27810));
    Sp12to4 I__4173 (
            .O(N__27810),
            .I(N__27807));
    Span12Mux_h I__4172 (
            .O(N__27807),
            .I(N__27803));
    InMux I__4171 (
            .O(N__27806),
            .I(N__27800));
    Odrv12 I__4170 (
            .O(N__27803),
            .I(RAM_DATA_cl_9Z0Z_15));
    LocalMux I__4169 (
            .O(N__27800),
            .I(RAM_DATA_cl_9Z0Z_15));
    CascadeMux I__4168 (
            .O(N__27795),
            .I(N_98_cascade_));
    IoInMux I__4167 (
            .O(N__27792),
            .I(N__27789));
    LocalMux I__4166 (
            .O(N__27789),
            .I(N__27786));
    IoSpan4Mux I__4165 (
            .O(N__27786),
            .I(N__27783));
    Span4Mux_s2_v I__4164 (
            .O(N__27783),
            .I(N__27780));
    Sp12to4 I__4163 (
            .O(N__27780),
            .I(N__27777));
    Span12Mux_s10_v I__4162 (
            .O(N__27777),
            .I(N__27773));
    InMux I__4161 (
            .O(N__27776),
            .I(N__27770));
    Odrv12 I__4160 (
            .O(N__27773),
            .I(RAM_DATA_clZ0Z_15));
    LocalMux I__4159 (
            .O(N__27770),
            .I(RAM_DATA_clZ0Z_15));
    InMux I__4158 (
            .O(N__27765),
            .I(N__27762));
    LocalMux I__4157 (
            .O(N__27762),
            .I(N__27759));
    Span4Mux_v I__4156 (
            .O(N__27759),
            .I(N__27756));
    Span4Mux_h I__4155 (
            .O(N__27756),
            .I(N__27753));
    Sp12to4 I__4154 (
            .O(N__27753),
            .I(N__27750));
    Span12Mux_v I__4153 (
            .O(N__27750),
            .I(N__27747));
    Span12Mux_h I__4152 (
            .O(N__27747),
            .I(N__27744));
    Odrv12 I__4151 (
            .O(N__27744),
            .I(RAM_DATA_in_6));
    CascadeMux I__4150 (
            .O(N__27741),
            .I(N__27738));
    InMux I__4149 (
            .O(N__27738),
            .I(N__27735));
    LocalMux I__4148 (
            .O(N__27735),
            .I(N__27732));
    Span4Mux_v I__4147 (
            .O(N__27732),
            .I(N__27729));
    Sp12to4 I__4146 (
            .O(N__27729),
            .I(N__27726));
    Span12Mux_h I__4145 (
            .O(N__27726),
            .I(N__27723));
    Odrv12 I__4144 (
            .O(N__27723),
            .I(RAM_DATA_in_14));
    InMux I__4143 (
            .O(N__27720),
            .I(N__27717));
    LocalMux I__4142 (
            .O(N__27717),
            .I(N__27714));
    Odrv4 I__4141 (
            .O(N__27714),
            .I(spi_data_misoZ0Z_6));
    InMux I__4140 (
            .O(N__27711),
            .I(N__27708));
    LocalMux I__4139 (
            .O(N__27708),
            .I(N__27705));
    Span4Mux_v I__4138 (
            .O(N__27705),
            .I(N__27702));
    Span4Mux_h I__4137 (
            .O(N__27702),
            .I(N__27699));
    Sp12to4 I__4136 (
            .O(N__27699),
            .I(N__27696));
    Span12Mux_v I__4135 (
            .O(N__27696),
            .I(N__27693));
    Span12Mux_h I__4134 (
            .O(N__27693),
            .I(N__27690));
    Odrv12 I__4133 (
            .O(N__27690),
            .I(RAM_DATA_in_7));
    InMux I__4132 (
            .O(N__27687),
            .I(N__27684));
    LocalMux I__4131 (
            .O(N__27684),
            .I(N__27681));
    Span4Mux_v I__4130 (
            .O(N__27681),
            .I(N__27678));
    Sp12to4 I__4129 (
            .O(N__27678),
            .I(N__27675));
    Span12Mux_h I__4128 (
            .O(N__27675),
            .I(N__27672));
    Odrv12 I__4127 (
            .O(N__27672),
            .I(RAM_DATA_in_15));
    InMux I__4126 (
            .O(N__27669),
            .I(N__27666));
    LocalMux I__4125 (
            .O(N__27666),
            .I(N__27663));
    Odrv4 I__4124 (
            .O(N__27663),
            .I(spi_data_misoZ0Z_7));
    IoInMux I__4123 (
            .O(N__27660),
            .I(N__27657));
    LocalMux I__4122 (
            .O(N__27657),
            .I(N__27654));
    IoSpan4Mux I__4121 (
            .O(N__27654),
            .I(N__27651));
    Span4Mux_s2_h I__4120 (
            .O(N__27651),
            .I(N__27648));
    Span4Mux_h I__4119 (
            .O(N__27648),
            .I(N__27645));
    Sp12to4 I__4118 (
            .O(N__27645),
            .I(N__27642));
    Span12Mux_h I__4117 (
            .O(N__27642),
            .I(N__27639));
    Odrv12 I__4116 (
            .O(N__27639),
            .I(RAM_nWE_0_i));
    InMux I__4115 (
            .O(N__27636),
            .I(N__27632));
    InMux I__4114 (
            .O(N__27635),
            .I(N__27629));
    LocalMux I__4113 (
            .O(N__27632),
            .I(N__27626));
    LocalMux I__4112 (
            .O(N__27629),
            .I(sADC_clk_prevZ0));
    Odrv12 I__4111 (
            .O(N__27626),
            .I(sADC_clk_prevZ0));
    InMux I__4110 (
            .O(N__27621),
            .I(N__27618));
    LocalMux I__4109 (
            .O(N__27618),
            .I(N__27612));
    InMux I__4108 (
            .O(N__27617),
            .I(N__27607));
    InMux I__4107 (
            .O(N__27616),
            .I(N__27607));
    IoInMux I__4106 (
            .O(N__27615),
            .I(N__27603));
    Span4Mux_h I__4105 (
            .O(N__27612),
            .I(N__27597));
    LocalMux I__4104 (
            .O(N__27607),
            .I(N__27597));
    InMux I__4103 (
            .O(N__27606),
            .I(N__27594));
    LocalMux I__4102 (
            .O(N__27603),
            .I(N__27591));
    InMux I__4101 (
            .O(N__27602),
            .I(N__27588));
    Span4Mux_v I__4100 (
            .O(N__27597),
            .I(N__27583));
    LocalMux I__4099 (
            .O(N__27594),
            .I(N__27583));
    Odrv12 I__4098 (
            .O(N__27591),
            .I(ADC_clk_c));
    LocalMux I__4097 (
            .O(N__27588),
            .I(ADC_clk_c));
    Odrv4 I__4096 (
            .O(N__27583),
            .I(ADC_clk_c));
    CascadeMux I__4095 (
            .O(N__27576),
            .I(N__27572));
    InMux I__4094 (
            .O(N__27575),
            .I(N__27569));
    InMux I__4093 (
            .O(N__27572),
            .I(N__27565));
    LocalMux I__4092 (
            .O(N__27569),
            .I(N__27562));
    InMux I__4091 (
            .O(N__27568),
            .I(N__27559));
    LocalMux I__4090 (
            .O(N__27565),
            .I(N__27556));
    Span4Mux_h I__4089 (
            .O(N__27562),
            .I(N__27553));
    LocalMux I__4088 (
            .O(N__27559),
            .I(N__27546));
    Span4Mux_v I__4087 (
            .O(N__27556),
            .I(N__27546));
    Span4Mux_v I__4086 (
            .O(N__27553),
            .I(N__27546));
    Odrv4 I__4085 (
            .O(N__27546),
            .I(N_127));
    SRMux I__4084 (
            .O(N__27543),
            .I(N__27537));
    SRMux I__4083 (
            .O(N__27542),
            .I(N__27533));
    SRMux I__4082 (
            .O(N__27541),
            .I(N__27530));
    SRMux I__4081 (
            .O(N__27540),
            .I(N__27527));
    LocalMux I__4080 (
            .O(N__27537),
            .I(N__27524));
    SRMux I__4079 (
            .O(N__27536),
            .I(N__27521));
    LocalMux I__4078 (
            .O(N__27533),
            .I(N__27518));
    LocalMux I__4077 (
            .O(N__27530),
            .I(N__27515));
    LocalMux I__4076 (
            .O(N__27527),
            .I(N__27512));
    Span4Mux_h I__4075 (
            .O(N__27524),
            .I(N__27505));
    LocalMux I__4074 (
            .O(N__27521),
            .I(N__27505));
    Span4Mux_v I__4073 (
            .O(N__27518),
            .I(N__27505));
    Span4Mux_v I__4072 (
            .O(N__27515),
            .I(N__27502));
    Span4Mux_h I__4071 (
            .O(N__27512),
            .I(N__27499));
    Span4Mux_v I__4070 (
            .O(N__27505),
            .I(N__27496));
    Span4Mux_h I__4069 (
            .O(N__27502),
            .I(N__27491));
    Span4Mux_v I__4068 (
            .O(N__27499),
            .I(N__27491));
    Odrv4 I__4067 (
            .O(N__27496),
            .I(N_1470_i));
    Odrv4 I__4066 (
            .O(N__27491),
            .I(N_1470_i));
    CascadeMux I__4065 (
            .O(N__27486),
            .I(N__27483));
    InMux I__4064 (
            .O(N__27483),
            .I(N__27480));
    LocalMux I__4063 (
            .O(N__27480),
            .I(N__27477));
    Odrv4 I__4062 (
            .O(N__27477),
            .I(N_86));
    InMux I__4061 (
            .O(N__27474),
            .I(N__27471));
    LocalMux I__4060 (
            .O(N__27471),
            .I(N__27467));
    InMux I__4059 (
            .O(N__27470),
            .I(N__27464));
    Span4Mux_h I__4058 (
            .O(N__27467),
            .I(N__27461));
    LocalMux I__4057 (
            .O(N__27464),
            .I(sRead_dataZ0));
    Odrv4 I__4056 (
            .O(N__27461),
            .I(sRead_dataZ0));
    InMux I__4055 (
            .O(N__27456),
            .I(N__27453));
    LocalMux I__4054 (
            .O(N__27453),
            .I(N__27449));
    InMux I__4053 (
            .O(N__27452),
            .I(N__27446));
    Span4Mux_h I__4052 (
            .O(N__27449),
            .I(N__27443));
    LocalMux I__4051 (
            .O(N__27446),
            .I(sCounterRAMZ0Z_5));
    Odrv4 I__4050 (
            .O(N__27443),
            .I(sCounterRAMZ0Z_5));
    InMux I__4049 (
            .O(N__27438),
            .I(N__27434));
    CascadeMux I__4048 (
            .O(N__27437),
            .I(N__27431));
    LocalMux I__4047 (
            .O(N__27434),
            .I(N__27428));
    InMux I__4046 (
            .O(N__27431),
            .I(N__27425));
    Span4Mux_h I__4045 (
            .O(N__27428),
            .I(N__27422));
    LocalMux I__4044 (
            .O(N__27425),
            .I(sCounterRAMZ0Z_4));
    Odrv4 I__4043 (
            .O(N__27422),
            .I(sCounterRAMZ0Z_4));
    CascadeMux I__4042 (
            .O(N__27417),
            .I(N__27414));
    InMux I__4041 (
            .O(N__27414),
            .I(N__27411));
    LocalMux I__4040 (
            .O(N__27411),
            .I(N__27407));
    InMux I__4039 (
            .O(N__27410),
            .I(N__27404));
    Span4Mux_h I__4038 (
            .O(N__27407),
            .I(N__27401));
    LocalMux I__4037 (
            .O(N__27404),
            .I(sCounterRAMZ0Z_7));
    Odrv4 I__4036 (
            .O(N__27401),
            .I(sCounterRAMZ0Z_7));
    InMux I__4035 (
            .O(N__27396),
            .I(N__27393));
    LocalMux I__4034 (
            .O(N__27393),
            .I(N__27389));
    InMux I__4033 (
            .O(N__27392),
            .I(N__27386));
    Span4Mux_v I__4032 (
            .O(N__27389),
            .I(N__27383));
    LocalMux I__4031 (
            .O(N__27386),
            .I(sCounterRAMZ0Z_0));
    Odrv4 I__4030 (
            .O(N__27383),
            .I(sCounterRAMZ0Z_0));
    InMux I__4029 (
            .O(N__27378),
            .I(N__27375));
    LocalMux I__4028 (
            .O(N__27375),
            .I(N__27372));
    Span12Mux_s10_v I__4027 (
            .O(N__27372),
            .I(N__27369));
    Odrv12 I__4026 (
            .O(N__27369),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_5 ));
    InMux I__4025 (
            .O(N__27366),
            .I(N__27363));
    LocalMux I__4024 (
            .O(N__27363),
            .I(N__27360));
    Odrv12 I__4023 (
            .O(N__27360),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_6 ));
    InMux I__4022 (
            .O(N__27357),
            .I(N__27354));
    LocalMux I__4021 (
            .O(N__27354),
            .I(N__27351));
    Odrv12 I__4020 (
            .O(N__27351),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_7 ));
    CEMux I__4019 (
            .O(N__27348),
            .I(N__27345));
    LocalMux I__4018 (
            .O(N__27345),
            .I(\spi_slave_inst.un4_i_wr ));
    InMux I__4017 (
            .O(N__27342),
            .I(N__27336));
    InMux I__4016 (
            .O(N__27341),
            .I(N__27336));
    LocalMux I__4015 (
            .O(N__27336),
            .I(spi_mosi_ready64_prevZ0Z2));
    InMux I__4014 (
            .O(N__27333),
            .I(N__27327));
    InMux I__4013 (
            .O(N__27332),
            .I(N__27327));
    LocalMux I__4012 (
            .O(N__27327),
            .I(spi_mosi_ready64_prevZ0));
    CascadeMux I__4011 (
            .O(N__27324),
            .I(N__27321));
    InMux I__4010 (
            .O(N__27321),
            .I(N__27318));
    LocalMux I__4009 (
            .O(N__27318),
            .I(spi_mosi_ready64_prevZ0Z3));
    InMux I__4008 (
            .O(N__27315),
            .I(N__27306));
    InMux I__4007 (
            .O(N__27314),
            .I(N__27306));
    InMux I__4006 (
            .O(N__27313),
            .I(N__27303));
    InMux I__4005 (
            .O(N__27312),
            .I(N__27298));
    InMux I__4004 (
            .O(N__27311),
            .I(N__27298));
    LocalMux I__4003 (
            .O(N__27306),
            .I(spi_mosi_ready));
    LocalMux I__4002 (
            .O(N__27303),
            .I(spi_mosi_ready));
    LocalMux I__4001 (
            .O(N__27298),
            .I(spi_mosi_ready));
    CascadeMux I__4000 (
            .O(N__27291),
            .I(spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_));
    IoInMux I__3999 (
            .O(N__27288),
            .I(N__27285));
    LocalMux I__3998 (
            .O(N__27285),
            .I(N__27282));
    Span12Mux_s3_v I__3997 (
            .O(N__27282),
            .I(N__27279));
    Span12Mux_v I__3996 (
            .O(N__27279),
            .I(N__27276));
    Odrv12 I__3995 (
            .O(N__27276),
            .I(LED3_c_i));
    InMux I__3994 (
            .O(N__27273),
            .I(N__27270));
    LocalMux I__3993 (
            .O(N__27270),
            .I(N__27267));
    Odrv12 I__3992 (
            .O(N__27267),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_0 ));
    InMux I__3991 (
            .O(N__27264),
            .I(N__27261));
    LocalMux I__3990 (
            .O(N__27261),
            .I(N__27258));
    Odrv4 I__3989 (
            .O(N__27258),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_1 ));
    InMux I__3988 (
            .O(N__27255),
            .I(N__27252));
    LocalMux I__3987 (
            .O(N__27252),
            .I(N__27249));
    Odrv4 I__3986 (
            .O(N__27249),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_2 ));
    InMux I__3985 (
            .O(N__27246),
            .I(N__27243));
    LocalMux I__3984 (
            .O(N__27243),
            .I(N__27240));
    Odrv12 I__3983 (
            .O(N__27240),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_3 ));
    InMux I__3982 (
            .O(N__27237),
            .I(N__27234));
    LocalMux I__3981 (
            .O(N__27234),
            .I(N__27231));
    Span4Mux_h I__3980 (
            .O(N__27231),
            .I(N__27228));
    Span4Mux_v I__3979 (
            .O(N__27228),
            .I(N__27225));
    Odrv4 I__3978 (
            .O(N__27225),
            .I(\spi_slave_inst.data_in_reg_iZ0Z_4 ));
    CascadeMux I__3977 (
            .O(N__27222),
            .I(N_206_cascade_));
    CEMux I__3976 (
            .O(N__27219),
            .I(N__27216));
    LocalMux I__3975 (
            .O(N__27216),
            .I(N__27213));
    Span4Mux_v I__3974 (
            .O(N__27213),
            .I(N__27210));
    Span4Mux_v I__3973 (
            .O(N__27210),
            .I(N__27207));
    Odrv4 I__3972 (
            .O(N__27207),
            .I(sAddress_RNIA6242_1Z0Z_0));
    InMux I__3971 (
            .O(N__27204),
            .I(N__27201));
    LocalMux I__3970 (
            .O(N__27201),
            .I(N__27198));
    Odrv4 I__3969 (
            .O(N__27198),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_3 ));
    InMux I__3968 (
            .O(N__27195),
            .I(N__27192));
    LocalMux I__3967 (
            .O(N__27192),
            .I(N__27189));
    Odrv4 I__3966 (
            .O(N__27189),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_7 ));
    InMux I__3965 (
            .O(N__27186),
            .I(N__27183));
    LocalMux I__3964 (
            .O(N__27183),
            .I(N__27180));
    Odrv12 I__3963 (
            .O(N__27180),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_5 ));
    InMux I__3962 (
            .O(N__27177),
            .I(N__27174));
    LocalMux I__3961 (
            .O(N__27174),
            .I(N__27171));
    Odrv4 I__3960 (
            .O(N__27171),
            .I(\spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1 ));
    InMux I__3959 (
            .O(N__27168),
            .I(N__27165));
    LocalMux I__3958 (
            .O(N__27165),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_1 ));
    InMux I__3957 (
            .O(N__27162),
            .I(N__27159));
    LocalMux I__3956 (
            .O(N__27159),
            .I(N__27156));
    Odrv4 I__3955 (
            .O(N__27156),
            .I(\spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2 ));
    InMux I__3954 (
            .O(N__27153),
            .I(N__27150));
    LocalMux I__3953 (
            .O(N__27150),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_2 ));
    InMux I__3952 (
            .O(N__27147),
            .I(N__27144));
    LocalMux I__3951 (
            .O(N__27144),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_6 ));
    CascadeMux I__3950 (
            .O(N__27141),
            .I(N__27138));
    InMux I__3949 (
            .O(N__27138),
            .I(N__27135));
    LocalMux I__3948 (
            .O(N__27135),
            .I(N__27132));
    Odrv4 I__3947 (
            .O(N__27132),
            .I(N_206));
    CascadeMux I__3946 (
            .O(N__27129),
            .I(\spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3_cascade_ ));
    InMux I__3945 (
            .O(N__27126),
            .I(N__27123));
    LocalMux I__3944 (
            .O(N__27123),
            .I(\spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0 ));
    InMux I__3943 (
            .O(N__27120),
            .I(N__27117));
    LocalMux I__3942 (
            .O(N__27117),
            .I(\spi_slave_inst.N_1394 ));
    CascadeMux I__3941 (
            .O(N__27114),
            .I(\spi_slave_inst.N_1397_cascade_ ));
    InMux I__3940 (
            .O(N__27111),
            .I(N__27108));
    LocalMux I__3939 (
            .O(N__27108),
            .I(\spi_slave_inst.tx_done_reg1_iZ0 ));
    InMux I__3938 (
            .O(N__27105),
            .I(N__27101));
    InMux I__3937 (
            .O(N__27104),
            .I(N__27098));
    LocalMux I__3936 (
            .O(N__27101),
            .I(N__27095));
    LocalMux I__3935 (
            .O(N__27098),
            .I(\spi_slave_inst.tx_done_reg2_iZ0 ));
    Odrv4 I__3934 (
            .O(N__27095),
            .I(\spi_slave_inst.tx_done_reg2_iZ0 ));
    InMux I__3933 (
            .O(N__27090),
            .I(N__27087));
    LocalMux I__3932 (
            .O(N__27087),
            .I(N__27084));
    Span4Mux_v I__3931 (
            .O(N__27084),
            .I(N__27081));
    Odrv4 I__3930 (
            .O(N__27081),
            .I(\spi_slave_inst.tx_done_reg3_iZ0 ));
    InMux I__3929 (
            .O(N__27078),
            .I(N__27075));
    LocalMux I__3928 (
            .O(N__27075),
            .I(N__27072));
    Span4Mux_v I__3927 (
            .O(N__27072),
            .I(N__27069));
    Odrv4 I__3926 (
            .O(N__27069),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_0 ));
    InMux I__3925 (
            .O(N__27066),
            .I(N__27062));
    InMux I__3924 (
            .O(N__27065),
            .I(N__27059));
    LocalMux I__3923 (
            .O(N__27062),
            .I(\spi_slave_inst.rx_done_neg_sclk_iZ0 ));
    LocalMux I__3922 (
            .O(N__27059),
            .I(\spi_slave_inst.rx_done_neg_sclk_iZ0 ));
    InMux I__3921 (
            .O(N__27054),
            .I(N__27051));
    LocalMux I__3920 (
            .O(N__27051),
            .I(\spi_slave_inst.rx_done_pos_sclk_iZ0 ));
    InMux I__3919 (
            .O(N__27048),
            .I(N__27045));
    LocalMux I__3918 (
            .O(N__27045),
            .I(\spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0 ));
    InMux I__3917 (
            .O(N__27042),
            .I(N__27036));
    InMux I__3916 (
            .O(N__27041),
            .I(N__27036));
    LocalMux I__3915 (
            .O(N__27036),
            .I(\spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0 ));
    InMux I__3914 (
            .O(N__27033),
            .I(N__27030));
    LocalMux I__3913 (
            .O(N__27030),
            .I(N__27027));
    Span4Mux_v I__3912 (
            .O(N__27027),
            .I(N__27023));
    CascadeMux I__3911 (
            .O(N__27026),
            .I(N__27020));
    Sp12to4 I__3910 (
            .O(N__27023),
            .I(N__27017));
    InMux I__3909 (
            .O(N__27020),
            .I(N__27014));
    Odrv12 I__3908 (
            .O(N__27017),
            .I(\spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0 ));
    LocalMux I__3907 (
            .O(N__27014),
            .I(\spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0 ));
    InMux I__3906 (
            .O(N__27009),
            .I(N__27006));
    LocalMux I__3905 (
            .O(N__27006),
            .I(\spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0 ));
    InMux I__3904 (
            .O(N__27003),
            .I(N__26995));
    InMux I__3903 (
            .O(N__27002),
            .I(N__26995));
    InMux I__3902 (
            .O(N__27001),
            .I(N__26989));
    InMux I__3901 (
            .O(N__27000),
            .I(N__26989));
    LocalMux I__3900 (
            .O(N__26995),
            .I(N__26986));
    InMux I__3899 (
            .O(N__26994),
            .I(N__26983));
    LocalMux I__3898 (
            .O(N__26989),
            .I(N__26980));
    Span4Mux_v I__3897 (
            .O(N__26986),
            .I(N__26977));
    LocalMux I__3896 (
            .O(N__26983),
            .I(N__26974));
    Span4Mux_v I__3895 (
            .O(N__26980),
            .I(N__26971));
    Span4Mux_h I__3894 (
            .O(N__26977),
            .I(N__26966));
    Span4Mux_v I__3893 (
            .O(N__26974),
            .I(N__26966));
    Span4Mux_h I__3892 (
            .O(N__26971),
            .I(N__26963));
    Odrv4 I__3891 (
            .O(N__26966),
            .I(\spi_master_inst.sclk_gen_u0.spi_start_iZ0 ));
    Odrv4 I__3890 (
            .O(N__26963),
            .I(\spi_master_inst.sclk_gen_u0.spi_start_iZ0 ));
    InMux I__3889 (
            .O(N__26958),
            .I(N__26955));
    LocalMux I__3888 (
            .O(N__26955),
            .I(\spi_slave_inst.txdata_reg_iZ0Z_4 ));
    InMux I__3887 (
            .O(N__26952),
            .I(N__26949));
    LocalMux I__3886 (
            .O(N__26949),
            .I(sEEDelayACQZ0Z_9));
    CEMux I__3885 (
            .O(N__26946),
            .I(N__26943));
    LocalMux I__3884 (
            .O(N__26943),
            .I(N__26940));
    Span4Mux_v I__3883 (
            .O(N__26940),
            .I(N__26937));
    Odrv4 I__3882 (
            .O(N__26937),
            .I(sAddress_RNIA6242Z0Z_0));
    CascadeMux I__3881 (
            .O(N__26934),
            .I(N_99_cascade_));
    IoInMux I__3880 (
            .O(N__26931),
            .I(N__26928));
    LocalMux I__3879 (
            .O(N__26928),
            .I(N__26925));
    Span4Mux_s2_v I__3878 (
            .O(N__26925),
            .I(N__26922));
    Span4Mux_h I__3877 (
            .O(N__26922),
            .I(N__26919));
    Span4Mux_h I__3876 (
            .O(N__26919),
            .I(N__26916));
    Span4Mux_h I__3875 (
            .O(N__26916),
            .I(N__26913));
    Span4Mux_v I__3874 (
            .O(N__26913),
            .I(N__26909));
    InMux I__3873 (
            .O(N__26912),
            .I(N__26906));
    Odrv4 I__3872 (
            .O(N__26909),
            .I(RAM_DATA_cl_12Z0Z_15));
    LocalMux I__3871 (
            .O(N__26906),
            .I(RAM_DATA_cl_12Z0Z_15));
    CascadeMux I__3870 (
            .O(N__26901),
            .I(N_94_cascade_));
    IoInMux I__3869 (
            .O(N__26898),
            .I(N__26895));
    LocalMux I__3868 (
            .O(N__26895),
            .I(N__26892));
    IoSpan4Mux I__3867 (
            .O(N__26892),
            .I(N__26889));
    Span4Mux_s2_h I__3866 (
            .O(N__26889),
            .I(N__26886));
    Sp12to4 I__3865 (
            .O(N__26886),
            .I(N__26883));
    Span12Mux_v I__3864 (
            .O(N__26883),
            .I(N__26880));
    Span12Mux_h I__3863 (
            .O(N__26880),
            .I(N__26876));
    InMux I__3862 (
            .O(N__26879),
            .I(N__26873));
    Odrv12 I__3861 (
            .O(N__26876),
            .I(RAM_DATA_cl_11Z0Z_15));
    LocalMux I__3860 (
            .O(N__26873),
            .I(RAM_DATA_cl_11Z0Z_15));
    CascadeMux I__3859 (
            .O(N__26868),
            .I(N_104_cascade_));
    IoInMux I__3858 (
            .O(N__26865),
            .I(N__26862));
    LocalMux I__3857 (
            .O(N__26862),
            .I(N__26859));
    Span4Mux_s0_v I__3856 (
            .O(N__26859),
            .I(N__26856));
    Sp12to4 I__3855 (
            .O(N__26856),
            .I(N__26853));
    Span12Mux_h I__3854 (
            .O(N__26853),
            .I(N__26849));
    InMux I__3853 (
            .O(N__26852),
            .I(N__26846));
    Odrv12 I__3852 (
            .O(N__26849),
            .I(RAM_DATA_cl_14Z0Z_15));
    LocalMux I__3851 (
            .O(N__26846),
            .I(RAM_DATA_cl_14Z0Z_15));
    InMux I__3850 (
            .O(N__26841),
            .I(N__26838));
    LocalMux I__3849 (
            .O(N__26838),
            .I(N__26835));
    Span4Mux_v I__3848 (
            .O(N__26835),
            .I(N__26832));
    Odrv4 I__3847 (
            .O(N__26832),
            .I(sDAC_dataZ0Z_2));
    InMux I__3846 (
            .O(N__26829),
            .I(N__26823));
    InMux I__3845 (
            .O(N__26828),
            .I(N__26820));
    InMux I__3844 (
            .O(N__26827),
            .I(N__26815));
    InMux I__3843 (
            .O(N__26826),
            .I(N__26815));
    LocalMux I__3842 (
            .O(N__26823),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_i6 ));
    LocalMux I__3841 (
            .O(N__26820),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_i6 ));
    LocalMux I__3840 (
            .O(N__26815),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_i6 ));
    InMux I__3839 (
            .O(N__26808),
            .I(N__26805));
    LocalMux I__3838 (
            .O(N__26805),
            .I(sEEDelayACQZ0Z_6));
    InMux I__3837 (
            .O(N__26802),
            .I(N__26799));
    LocalMux I__3836 (
            .O(N__26799),
            .I(sEEDelayACQZ0Z_7));
    InMux I__3835 (
            .O(N__26796),
            .I(N__26793));
    LocalMux I__3834 (
            .O(N__26793),
            .I(sEEDelayACQZ0Z_10));
    InMux I__3833 (
            .O(N__26790),
            .I(N__26787));
    LocalMux I__3832 (
            .O(N__26787),
            .I(sEEDelayACQZ0Z_11));
    InMux I__3831 (
            .O(N__26784),
            .I(N__26781));
    LocalMux I__3830 (
            .O(N__26781),
            .I(sEEDelayACQZ0Z_12));
    InMux I__3829 (
            .O(N__26778),
            .I(N__26775));
    LocalMux I__3828 (
            .O(N__26775),
            .I(sEEDelayACQZ0Z_13));
    InMux I__3827 (
            .O(N__26772),
            .I(N__26769));
    LocalMux I__3826 (
            .O(N__26769),
            .I(sEEDelayACQZ0Z_14));
    InMux I__3825 (
            .O(N__26766),
            .I(N__26763));
    LocalMux I__3824 (
            .O(N__26763),
            .I(sEEDelayACQZ0Z_15));
    InMux I__3823 (
            .O(N__26760),
            .I(N__26757));
    LocalMux I__3822 (
            .O(N__26757),
            .I(sEEDelayACQZ0Z_8));
    CEMux I__3821 (
            .O(N__26754),
            .I(N__26751));
    LocalMux I__3820 (
            .O(N__26751),
            .I(N__26748));
    Span4Mux_v I__3819 (
            .O(N__26748),
            .I(N__26745));
    Odrv4 I__3818 (
            .O(N__26745),
            .I(N_76_i));
    CascadeMux I__3817 (
            .O(N__26742),
            .I(N_71_cascade_));
    InMux I__3816 (
            .O(N__26739),
            .I(N__26736));
    LocalMux I__3815 (
            .O(N__26736),
            .I(sEEDelayACQZ0Z_0));
    InMux I__3814 (
            .O(N__26733),
            .I(N__26730));
    LocalMux I__3813 (
            .O(N__26730),
            .I(sEEDelayACQZ0Z_1));
    InMux I__3812 (
            .O(N__26727),
            .I(N__26724));
    LocalMux I__3811 (
            .O(N__26724),
            .I(sEEDelayACQZ0Z_2));
    InMux I__3810 (
            .O(N__26721),
            .I(N__26718));
    LocalMux I__3809 (
            .O(N__26718),
            .I(sEEDelayACQZ0Z_3));
    InMux I__3808 (
            .O(N__26715),
            .I(N__26712));
    LocalMux I__3807 (
            .O(N__26712),
            .I(sEEDelayACQZ0Z_4));
    InMux I__3806 (
            .O(N__26709),
            .I(N__26706));
    LocalMux I__3805 (
            .O(N__26706),
            .I(sEEDelayACQZ0Z_5));
    CascadeMux I__3804 (
            .O(N__26703),
            .I(N__26700));
    InMux I__3803 (
            .O(N__26700),
            .I(N__26697));
    LocalMux I__3802 (
            .O(N__26697),
            .I(un1_sacqtime_cry_18_sf));
    CascadeMux I__3801 (
            .O(N__26694),
            .I(N__26691));
    InMux I__3800 (
            .O(N__26691),
            .I(N__26688));
    LocalMux I__3799 (
            .O(N__26688),
            .I(un1_sacqtime_cry_19_sf));
    CascadeMux I__3798 (
            .O(N__26685),
            .I(N__26682));
    InMux I__3797 (
            .O(N__26682),
            .I(N__26679));
    LocalMux I__3796 (
            .O(N__26679),
            .I(un1_sacqtime_cry_20_sf));
    CascadeMux I__3795 (
            .O(N__26676),
            .I(N__26673));
    InMux I__3794 (
            .O(N__26673),
            .I(N__26670));
    LocalMux I__3793 (
            .O(N__26670),
            .I(un1_sacqtime_cry_21_sf));
    CascadeMux I__3792 (
            .O(N__26667),
            .I(N__26664));
    InMux I__3791 (
            .O(N__26664),
            .I(N__26661));
    LocalMux I__3790 (
            .O(N__26661),
            .I(un1_sacqtime_cry_22_sf));
    CascadeMux I__3789 (
            .O(N__26658),
            .I(N__26655));
    InMux I__3788 (
            .O(N__26655),
            .I(N__26652));
    LocalMux I__3787 (
            .O(N__26652),
            .I(un1_sacqtime_cry_23_sf));
    InMux I__3786 (
            .O(N__26649),
            .I(bfn_10_17_0_));
    IoInMux I__3785 (
            .O(N__26646),
            .I(N__26643));
    LocalMux I__3784 (
            .O(N__26643),
            .I(N__26640));
    IoSpan4Mux I__3783 (
            .O(N__26640),
            .I(N__26637));
    Span4Mux_s2_h I__3782 (
            .O(N__26637),
            .I(N__26634));
    Sp12to4 I__3781 (
            .O(N__26634),
            .I(N__26631));
    Span12Mux_s9_h I__3780 (
            .O(N__26631),
            .I(N__26628));
    Span12Mux_h I__3779 (
            .O(N__26628),
            .I(N__26624));
    InMux I__3778 (
            .O(N__26627),
            .I(N__26621));
    Span12Mux_v I__3777 (
            .O(N__26624),
            .I(N__26618));
    LocalMux I__3776 (
            .O(N__26621),
            .I(N__26615));
    Odrv12 I__3775 (
            .O(N__26618),
            .I(RAM_DATA_cl_10Z0Z_15));
    Odrv4 I__3774 (
            .O(N__26615),
            .I(RAM_DATA_cl_10Z0Z_15));
    InMux I__3773 (
            .O(N__26610),
            .I(N__26607));
    LocalMux I__3772 (
            .O(N__26607),
            .I(N__26604));
    Odrv12 I__3771 (
            .O(N__26604),
            .I(N_106));
    IoInMux I__3770 (
            .O(N__26601),
            .I(N__26598));
    LocalMux I__3769 (
            .O(N__26598),
            .I(N__26595));
    IoSpan4Mux I__3768 (
            .O(N__26595),
            .I(N__26592));
    Span4Mux_s2_v I__3767 (
            .O(N__26592),
            .I(N__26589));
    Span4Mux_v I__3766 (
            .O(N__26589),
            .I(N__26586));
    Odrv4 I__3765 (
            .O(N__26586),
            .I(N_26));
    CascadeMux I__3764 (
            .O(N__26583),
            .I(N__26579));
    CascadeMux I__3763 (
            .O(N__26582),
            .I(N__26576));
    InMux I__3762 (
            .O(N__26579),
            .I(N__26573));
    InMux I__3761 (
            .O(N__26576),
            .I(N__26570));
    LocalMux I__3760 (
            .O(N__26573),
            .I(sCounter_i_10));
    LocalMux I__3759 (
            .O(N__26570),
            .I(sCounter_i_10));
    CascadeMux I__3758 (
            .O(N__26565),
            .I(N__26561));
    CascadeMux I__3757 (
            .O(N__26564),
            .I(N__26558));
    InMux I__3756 (
            .O(N__26561),
            .I(N__26555));
    InMux I__3755 (
            .O(N__26558),
            .I(N__26552));
    LocalMux I__3754 (
            .O(N__26555),
            .I(sCounter_i_11));
    LocalMux I__3753 (
            .O(N__26552),
            .I(sCounter_i_11));
    CascadeMux I__3752 (
            .O(N__26547),
            .I(N__26543));
    CascadeMux I__3751 (
            .O(N__26546),
            .I(N__26540));
    InMux I__3750 (
            .O(N__26543),
            .I(N__26537));
    InMux I__3749 (
            .O(N__26540),
            .I(N__26534));
    LocalMux I__3748 (
            .O(N__26537),
            .I(sCounter_i_12));
    LocalMux I__3747 (
            .O(N__26534),
            .I(sCounter_i_12));
    CascadeMux I__3746 (
            .O(N__26529),
            .I(N__26525));
    CascadeMux I__3745 (
            .O(N__26528),
            .I(N__26522));
    InMux I__3744 (
            .O(N__26525),
            .I(N__26519));
    InMux I__3743 (
            .O(N__26522),
            .I(N__26516));
    LocalMux I__3742 (
            .O(N__26519),
            .I(sCounter_i_13));
    LocalMux I__3741 (
            .O(N__26516),
            .I(sCounter_i_13));
    CascadeMux I__3740 (
            .O(N__26511),
            .I(N__26507));
    CascadeMux I__3739 (
            .O(N__26510),
            .I(N__26504));
    InMux I__3738 (
            .O(N__26507),
            .I(N__26501));
    InMux I__3737 (
            .O(N__26504),
            .I(N__26498));
    LocalMux I__3736 (
            .O(N__26501),
            .I(sCounter_i_14));
    LocalMux I__3735 (
            .O(N__26498),
            .I(sCounter_i_14));
    CascadeMux I__3734 (
            .O(N__26493),
            .I(N__26489));
    InMux I__3733 (
            .O(N__26492),
            .I(N__26486));
    InMux I__3732 (
            .O(N__26489),
            .I(N__26483));
    LocalMux I__3731 (
            .O(N__26486),
            .I(sCounter_i_15));
    LocalMux I__3730 (
            .O(N__26483),
            .I(sCounter_i_15));
    CascadeMux I__3729 (
            .O(N__26478),
            .I(N__26475));
    InMux I__3728 (
            .O(N__26475),
            .I(N__26472));
    LocalMux I__3727 (
            .O(N__26472),
            .I(un1_sacqtime_cry_16_sf));
    CascadeMux I__3726 (
            .O(N__26469),
            .I(N__26466));
    InMux I__3725 (
            .O(N__26466),
            .I(N__26463));
    LocalMux I__3724 (
            .O(N__26463),
            .I(un1_sacqtime_cry_17_sf));
    CascadeMux I__3723 (
            .O(N__26460),
            .I(N__26456));
    CascadeMux I__3722 (
            .O(N__26459),
            .I(N__26453));
    InMux I__3721 (
            .O(N__26456),
            .I(N__26450));
    InMux I__3720 (
            .O(N__26453),
            .I(N__26447));
    LocalMux I__3719 (
            .O(N__26450),
            .I(sCounter_i_2));
    LocalMux I__3718 (
            .O(N__26447),
            .I(sCounter_i_2));
    CascadeMux I__3717 (
            .O(N__26442),
            .I(N__26438));
    CascadeMux I__3716 (
            .O(N__26441),
            .I(N__26435));
    InMux I__3715 (
            .O(N__26438),
            .I(N__26432));
    InMux I__3714 (
            .O(N__26435),
            .I(N__26429));
    LocalMux I__3713 (
            .O(N__26432),
            .I(sCounter_i_3));
    LocalMux I__3712 (
            .O(N__26429),
            .I(sCounter_i_3));
    CascadeMux I__3711 (
            .O(N__26424),
            .I(N__26420));
    CascadeMux I__3710 (
            .O(N__26423),
            .I(N__26417));
    InMux I__3709 (
            .O(N__26420),
            .I(N__26414));
    InMux I__3708 (
            .O(N__26417),
            .I(N__26411));
    LocalMux I__3707 (
            .O(N__26414),
            .I(sCounter_i_4));
    LocalMux I__3706 (
            .O(N__26411),
            .I(sCounter_i_4));
    CascadeMux I__3705 (
            .O(N__26406),
            .I(N__26402));
    CascadeMux I__3704 (
            .O(N__26405),
            .I(N__26399));
    InMux I__3703 (
            .O(N__26402),
            .I(N__26396));
    InMux I__3702 (
            .O(N__26399),
            .I(N__26393));
    LocalMux I__3701 (
            .O(N__26396),
            .I(sCounter_i_5));
    LocalMux I__3700 (
            .O(N__26393),
            .I(sCounter_i_5));
    CascadeMux I__3699 (
            .O(N__26388),
            .I(N__26384));
    CascadeMux I__3698 (
            .O(N__26387),
            .I(N__26381));
    InMux I__3697 (
            .O(N__26384),
            .I(N__26378));
    InMux I__3696 (
            .O(N__26381),
            .I(N__26375));
    LocalMux I__3695 (
            .O(N__26378),
            .I(sCounter_i_6));
    LocalMux I__3694 (
            .O(N__26375),
            .I(sCounter_i_6));
    CascadeMux I__3693 (
            .O(N__26370),
            .I(N__26367));
    InMux I__3692 (
            .O(N__26367),
            .I(N__26363));
    CascadeMux I__3691 (
            .O(N__26366),
            .I(N__26360));
    LocalMux I__3690 (
            .O(N__26363),
            .I(N__26357));
    InMux I__3689 (
            .O(N__26360),
            .I(N__26354));
    Odrv4 I__3688 (
            .O(N__26357),
            .I(sCounter_i_7));
    LocalMux I__3687 (
            .O(N__26354),
            .I(sCounter_i_7));
    CascadeMux I__3686 (
            .O(N__26349),
            .I(N__26345));
    CascadeMux I__3685 (
            .O(N__26348),
            .I(N__26342));
    InMux I__3684 (
            .O(N__26345),
            .I(N__26339));
    InMux I__3683 (
            .O(N__26342),
            .I(N__26336));
    LocalMux I__3682 (
            .O(N__26339),
            .I(sCounter_i_8));
    LocalMux I__3681 (
            .O(N__26336),
            .I(sCounter_i_8));
    CascadeMux I__3680 (
            .O(N__26331),
            .I(N__26327));
    CascadeMux I__3679 (
            .O(N__26330),
            .I(N__26324));
    InMux I__3678 (
            .O(N__26327),
            .I(N__26321));
    InMux I__3677 (
            .O(N__26324),
            .I(N__26318));
    LocalMux I__3676 (
            .O(N__26321),
            .I(sCounter_i_9));
    LocalMux I__3675 (
            .O(N__26318),
            .I(sCounter_i_9));
    CascadeMux I__3674 (
            .O(N__26313),
            .I(N__26310));
    InMux I__3673 (
            .O(N__26310),
            .I(N__26306));
    InMux I__3672 (
            .O(N__26309),
            .I(N__26303));
    LocalMux I__3671 (
            .O(N__26306),
            .I(N__26300));
    LocalMux I__3670 (
            .O(N__26303),
            .I(N__26295));
    Span4Mux_h I__3669 (
            .O(N__26300),
            .I(N__26292));
    InMux I__3668 (
            .O(N__26299),
            .I(N__26287));
    InMux I__3667 (
            .O(N__26298),
            .I(N__26287));
    Sp12to4 I__3666 (
            .O(N__26295),
            .I(N__26284));
    Span4Mux_v I__3665 (
            .O(N__26292),
            .I(N__26281));
    LocalMux I__3664 (
            .O(N__26287),
            .I(button_debounce_counterZ0Z_0));
    Odrv12 I__3663 (
            .O(N__26284),
            .I(button_debounce_counterZ0Z_0));
    Odrv4 I__3662 (
            .O(N__26281),
            .I(button_debounce_counterZ0Z_0));
    InMux I__3661 (
            .O(N__26274),
            .I(N__26271));
    LocalMux I__3660 (
            .O(N__26271),
            .I(N__26268));
    Span4Mux_v I__3659 (
            .O(N__26268),
            .I(N__26264));
    InMux I__3658 (
            .O(N__26267),
            .I(N__26261));
    Span4Mux_v I__3657 (
            .O(N__26264),
            .I(N__26258));
    LocalMux I__3656 (
            .O(N__26261),
            .I(N__26253));
    Span4Mux_h I__3655 (
            .O(N__26258),
            .I(N__26253));
    Odrv4 I__3654 (
            .O(N__26253),
            .I(button_debounce_counterZ0Z_1));
    InMux I__3653 (
            .O(N__26250),
            .I(N__26247));
    LocalMux I__3652 (
            .O(N__26247),
            .I(N__26244));
    Glb2LocalMux I__3651 (
            .O(N__26244),
            .I(N__26226));
    SRMux I__3650 (
            .O(N__26243),
            .I(N__26226));
    SRMux I__3649 (
            .O(N__26242),
            .I(N__26226));
    SRMux I__3648 (
            .O(N__26241),
            .I(N__26226));
    SRMux I__3647 (
            .O(N__26240),
            .I(N__26226));
    SRMux I__3646 (
            .O(N__26239),
            .I(N__26226));
    GlobalMux I__3645 (
            .O(N__26226),
            .I(N__26223));
    gio2CtrlBuf I__3644 (
            .O(N__26223),
            .I(N_3089_g));
    InMux I__3643 (
            .O(N__26220),
            .I(N__26216));
    InMux I__3642 (
            .O(N__26219),
            .I(N__26213));
    LocalMux I__3641 (
            .O(N__26216),
            .I(spi_mosi_ready_prevZ0Z2));
    LocalMux I__3640 (
            .O(N__26213),
            .I(spi_mosi_ready_prevZ0Z2));
    InMux I__3639 (
            .O(N__26208),
            .I(N__26204));
    InMux I__3638 (
            .O(N__26207),
            .I(N__26201));
    LocalMux I__3637 (
            .O(N__26204),
            .I(spi_mosi_ready_prevZ0));
    LocalMux I__3636 (
            .O(N__26201),
            .I(spi_mosi_ready_prevZ0));
    CascadeMux I__3635 (
            .O(N__26196),
            .I(N__26193));
    InMux I__3634 (
            .O(N__26193),
            .I(N__26190));
    LocalMux I__3633 (
            .O(N__26190),
            .I(spi_mosi_ready_prevZ0Z3));
    CascadeMux I__3632 (
            .O(N__26187),
            .I(spi_mosi_ready_prev3_RNILKERZ0_cascade_));
    InMux I__3631 (
            .O(N__26184),
            .I(N__26180));
    InMux I__3630 (
            .O(N__26183),
            .I(N__26177));
    LocalMux I__3629 (
            .O(N__26180),
            .I(N__26174));
    LocalMux I__3628 (
            .O(N__26177),
            .I(\spi_slave_inst.tx_ready_iZ0 ));
    Odrv4 I__3627 (
            .O(N__26174),
            .I(\spi_slave_inst.tx_ready_iZ0 ));
    CascadeMux I__3626 (
            .O(N__26169),
            .I(N__26165));
    CascadeMux I__3625 (
            .O(N__26168),
            .I(N__26162));
    InMux I__3624 (
            .O(N__26165),
            .I(N__26159));
    InMux I__3623 (
            .O(N__26162),
            .I(N__26156));
    LocalMux I__3622 (
            .O(N__26159),
            .I(sCounter_i_0));
    LocalMux I__3621 (
            .O(N__26156),
            .I(sCounter_i_0));
    InMux I__3620 (
            .O(N__26151),
            .I(N__26147));
    CascadeMux I__3619 (
            .O(N__26150),
            .I(N__26144));
    LocalMux I__3618 (
            .O(N__26147),
            .I(N__26141));
    InMux I__3617 (
            .O(N__26144),
            .I(N__26138));
    Odrv4 I__3616 (
            .O(N__26141),
            .I(sCounter_i_1));
    LocalMux I__3615 (
            .O(N__26138),
            .I(sCounter_i_1));
    InMux I__3614 (
            .O(N__26133),
            .I(N__26130));
    LocalMux I__3613 (
            .O(N__26130),
            .I(\spi_slave_inst.rx_done_reg3_iZ0 ));
    CascadeMux I__3612 (
            .O(N__26127),
            .I(\spi_slave_inst.rx_ready_i_RNOZ0Z_0_cascade_ ));
    CascadeMux I__3611 (
            .O(N__26124),
            .I(\spi_slave_inst.un4_tx_done_reg2_i_cascade_ ));
    CascadeMux I__3610 (
            .O(N__26121),
            .I(N__26117));
    CascadeMux I__3609 (
            .O(N__26120),
            .I(N__26112));
    InMux I__3608 (
            .O(N__26117),
            .I(N__26108));
    InMux I__3607 (
            .O(N__26116),
            .I(N__26099));
    InMux I__3606 (
            .O(N__26115),
            .I(N__26099));
    InMux I__3605 (
            .O(N__26112),
            .I(N__26099));
    InMux I__3604 (
            .O(N__26111),
            .I(N__26099));
    LocalMux I__3603 (
            .O(N__26108),
            .I(sEETrigCounterZ0Z_3));
    LocalMux I__3602 (
            .O(N__26099),
            .I(sEETrigCounterZ0Z_3));
    CascadeMux I__3601 (
            .O(N__26094),
            .I(N__26091));
    InMux I__3600 (
            .O(N__26091),
            .I(N__26088));
    LocalMux I__3599 (
            .O(N__26088),
            .I(N__26085));
    Odrv4 I__3598 (
            .O(N__26085),
            .I(un10_trig_prev_3));
    CascadeMux I__3597 (
            .O(N__26082),
            .I(N__26077));
    InMux I__3596 (
            .O(N__26081),
            .I(N__26071));
    InMux I__3595 (
            .O(N__26080),
            .I(N__26071));
    InMux I__3594 (
            .O(N__26077),
            .I(N__26066));
    InMux I__3593 (
            .O(N__26076),
            .I(N__26066));
    LocalMux I__3592 (
            .O(N__26071),
            .I(sEETrigCounterZ0Z_2));
    LocalMux I__3591 (
            .O(N__26066),
            .I(sEETrigCounterZ0Z_2));
    InMux I__3590 (
            .O(N__26061),
            .I(N__26058));
    LocalMux I__3589 (
            .O(N__26058),
            .I(un10_trig_prev_2));
    CascadeMux I__3588 (
            .O(N__26055),
            .I(N__26052));
    InMux I__3587 (
            .O(N__26052),
            .I(N__26049));
    LocalMux I__3586 (
            .O(N__26049),
            .I(N__26046));
    Odrv4 I__3585 (
            .O(N__26046),
            .I(un10_trig_prev_0));
    CascadeMux I__3584 (
            .O(N__26043),
            .I(N__26039));
    InMux I__3583 (
            .O(N__26042),
            .I(N__26026));
    InMux I__3582 (
            .O(N__26039),
            .I(N__26026));
    InMux I__3581 (
            .O(N__26038),
            .I(N__26026));
    InMux I__3580 (
            .O(N__26037),
            .I(N__26026));
    InMux I__3579 (
            .O(N__26036),
            .I(N__26021));
    InMux I__3578 (
            .O(N__26035),
            .I(N__26021));
    LocalMux I__3577 (
            .O(N__26026),
            .I(sEETrigCounterZ0Z_0));
    LocalMux I__3576 (
            .O(N__26021),
            .I(sEETrigCounterZ0Z_0));
    InMux I__3575 (
            .O(N__26016),
            .I(N__26005));
    InMux I__3574 (
            .O(N__26015),
            .I(N__26005));
    InMux I__3573 (
            .O(N__26014),
            .I(N__26005));
    InMux I__3572 (
            .O(N__26013),
            .I(N__26000));
    InMux I__3571 (
            .O(N__26012),
            .I(N__26000));
    LocalMux I__3570 (
            .O(N__26005),
            .I(sEETrigCounterZ0Z_1));
    LocalMux I__3569 (
            .O(N__26000),
            .I(sEETrigCounterZ0Z_1));
    CascadeMux I__3568 (
            .O(N__25995),
            .I(N__25992));
    InMux I__3567 (
            .O(N__25992),
            .I(N__25989));
    LocalMux I__3566 (
            .O(N__25989),
            .I(un10_trig_prev_1));
    InMux I__3565 (
            .O(N__25986),
            .I(N__25983));
    LocalMux I__3564 (
            .O(N__25983),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_15 ));
    InMux I__3563 (
            .O(N__25980),
            .I(N__25976));
    InMux I__3562 (
            .O(N__25979),
            .I(N__25973));
    LocalMux I__3561 (
            .O(N__25976),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0 ));
    LocalMux I__3560 (
            .O(N__25973),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0 ));
    InMux I__3559 (
            .O(N__25968),
            .I(bfn_10_6_0_));
    InMux I__3558 (
            .O(N__25965),
            .I(N__25961));
    InMux I__3557 (
            .O(N__25964),
            .I(N__25958));
    LocalMux I__3556 (
            .O(N__25961),
            .I(N__25953));
    LocalMux I__3555 (
            .O(N__25958),
            .I(N__25953));
    Odrv4 I__3554 (
            .O(N__25953),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1 ));
    InMux I__3553 (
            .O(N__25950),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0 ));
    CascadeMux I__3552 (
            .O(N__25947),
            .I(N__25943));
    InMux I__3551 (
            .O(N__25946),
            .I(N__25940));
    InMux I__3550 (
            .O(N__25943),
            .I(N__25937));
    LocalMux I__3549 (
            .O(N__25940),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2 ));
    LocalMux I__3548 (
            .O(N__25937),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2 ));
    InMux I__3547 (
            .O(N__25932),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1 ));
    InMux I__3546 (
            .O(N__25929),
            .I(N__25925));
    InMux I__3545 (
            .O(N__25928),
            .I(N__25922));
    LocalMux I__3544 (
            .O(N__25925),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3 ));
    LocalMux I__3543 (
            .O(N__25922),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3 ));
    InMux I__3542 (
            .O(N__25917),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2 ));
    InMux I__3541 (
            .O(N__25914),
            .I(N__25910));
    InMux I__3540 (
            .O(N__25913),
            .I(N__25907));
    LocalMux I__3539 (
            .O(N__25910),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4 ));
    LocalMux I__3538 (
            .O(N__25907),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4 ));
    InMux I__3537 (
            .O(N__25902),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3 ));
    InMux I__3536 (
            .O(N__25899),
            .I(N__25895));
    InMux I__3535 (
            .O(N__25898),
            .I(N__25892));
    LocalMux I__3534 (
            .O(N__25895),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5 ));
    LocalMux I__3533 (
            .O(N__25892),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5 ));
    InMux I__3532 (
            .O(N__25887),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4 ));
    CascadeMux I__3531 (
            .O(N__25884),
            .I(N__25880));
    InMux I__3530 (
            .O(N__25883),
            .I(N__25877));
    InMux I__3529 (
            .O(N__25880),
            .I(N__25874));
    LocalMux I__3528 (
            .O(N__25877),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6 ));
    LocalMux I__3527 (
            .O(N__25874),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6 ));
    InMux I__3526 (
            .O(N__25869),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5 ));
    InMux I__3525 (
            .O(N__25866),
            .I(N__25848));
    InMux I__3524 (
            .O(N__25865),
            .I(N__25848));
    InMux I__3523 (
            .O(N__25864),
            .I(N__25848));
    InMux I__3522 (
            .O(N__25863),
            .I(N__25848));
    InMux I__3521 (
            .O(N__25862),
            .I(N__25848));
    InMux I__3520 (
            .O(N__25861),
            .I(N__25841));
    InMux I__3519 (
            .O(N__25860),
            .I(N__25841));
    InMux I__3518 (
            .O(N__25859),
            .I(N__25841));
    LocalMux I__3517 (
            .O(N__25848),
            .I(N__25836));
    LocalMux I__3516 (
            .O(N__25841),
            .I(N__25836));
    Odrv4 I__3515 (
            .O(N__25836),
            .I(\spi_master_inst.sclk_gen_u0.falling_count_start_i_i ));
    InMux I__3514 (
            .O(N__25833),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6 ));
    InMux I__3513 (
            .O(N__25830),
            .I(N__25826));
    InMux I__3512 (
            .O(N__25829),
            .I(N__25823));
    LocalMux I__3511 (
            .O(N__25826),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7 ));
    LocalMux I__3510 (
            .O(N__25823),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7 ));
    CEMux I__3509 (
            .O(N__25818),
            .I(N__25815));
    LocalMux I__3508 (
            .O(N__25815),
            .I(N__25812));
    Span4Mux_h I__3507 (
            .O(N__25812),
            .I(N__25809));
    Sp12to4 I__3506 (
            .O(N__25809),
            .I(N__25806));
    Odrv12 I__3505 (
            .O(N__25806),
            .I(\spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i ));
    InMux I__3504 (
            .O(N__25803),
            .I(N__25800));
    LocalMux I__3503 (
            .O(N__25800),
            .I(\spi_slave_inst.un23_i_ssn_3 ));
    InMux I__3502 (
            .O(N__25797),
            .I(N__25792));
    InMux I__3501 (
            .O(N__25796),
            .I(N__25789));
    InMux I__3500 (
            .O(N__25795),
            .I(N__25786));
    LocalMux I__3499 (
            .O(N__25792),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5 ));
    LocalMux I__3498 (
            .O(N__25789),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5 ));
    LocalMux I__3497 (
            .O(N__25786),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5 ));
    CascadeMux I__3496 (
            .O(N__25779),
            .I(N__25775));
    InMux I__3495 (
            .O(N__25778),
            .I(N__25770));
    InMux I__3494 (
            .O(N__25775),
            .I(N__25767));
    InMux I__3493 (
            .O(N__25774),
            .I(N__25764));
    InMux I__3492 (
            .O(N__25773),
            .I(N__25761));
    LocalMux I__3491 (
            .O(N__25770),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2 ));
    LocalMux I__3490 (
            .O(N__25767),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2 ));
    LocalMux I__3489 (
            .O(N__25764),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2 ));
    LocalMux I__3488 (
            .O(N__25761),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2 ));
    InMux I__3487 (
            .O(N__25752),
            .I(N__25749));
    LocalMux I__3486 (
            .O(N__25749),
            .I(N__25746));
    Span12Mux_s9_h I__3485 (
            .O(N__25746),
            .I(N__25743));
    Odrv12 I__3484 (
            .O(N__25743),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_6 ));
    InMux I__3483 (
            .O(N__25740),
            .I(N__25737));
    LocalMux I__3482 (
            .O(N__25737),
            .I(N__25734));
    Span4Mux_v I__3481 (
            .O(N__25734),
            .I(N__25731));
    Odrv4 I__3480 (
            .O(N__25731),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_1 ));
    InMux I__3479 (
            .O(N__25728),
            .I(N__25725));
    LocalMux I__3478 (
            .O(N__25725),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_2 ));
    InMux I__3477 (
            .O(N__25722),
            .I(N__25719));
    LocalMux I__3476 (
            .O(N__25719),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_11 ));
    InMux I__3475 (
            .O(N__25716),
            .I(N__25713));
    LocalMux I__3474 (
            .O(N__25713),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_12 ));
    InMux I__3473 (
            .O(N__25710),
            .I(N__25707));
    LocalMux I__3472 (
            .O(N__25707),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_3 ));
    InMux I__3471 (
            .O(N__25704),
            .I(N__25701));
    LocalMux I__3470 (
            .O(N__25701),
            .I(N__25698));
    Span4Mux_h I__3469 (
            .O(N__25698),
            .I(N__25695));
    Odrv4 I__3468 (
            .O(N__25695),
            .I(\spi_master_inst.spi_data_path_u1.data_inZ0Z_14 ));
    InMux I__3467 (
            .O(N__25692),
            .I(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3 ));
    InMux I__3466 (
            .O(N__25689),
            .I(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4 ));
    InMux I__3465 (
            .O(N__25686),
            .I(N__25682));
    InMux I__3464 (
            .O(N__25685),
            .I(N__25679));
    LocalMux I__3463 (
            .O(N__25682),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4 ));
    LocalMux I__3462 (
            .O(N__25679),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4 ));
    InMux I__3461 (
            .O(N__25674),
            .I(N__25670));
    InMux I__3460 (
            .O(N__25673),
            .I(N__25667));
    LocalMux I__3459 (
            .O(N__25670),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1 ));
    LocalMux I__3458 (
            .O(N__25667),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1 ));
    CascadeMux I__3457 (
            .O(N__25662),
            .I(N__25658));
    InMux I__3456 (
            .O(N__25661),
            .I(N__25655));
    InMux I__3455 (
            .O(N__25658),
            .I(N__25652));
    LocalMux I__3454 (
            .O(N__25655),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0 ));
    LocalMux I__3453 (
            .O(N__25652),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0 ));
    InMux I__3452 (
            .O(N__25647),
            .I(N__25643));
    InMux I__3451 (
            .O(N__25646),
            .I(N__25640));
    LocalMux I__3450 (
            .O(N__25643),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3 ));
    LocalMux I__3449 (
            .O(N__25640),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3 ));
    InMux I__3448 (
            .O(N__25635),
            .I(N__25631));
    InMux I__3447 (
            .O(N__25634),
            .I(N__25628));
    LocalMux I__3446 (
            .O(N__25631),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5 ));
    LocalMux I__3445 (
            .O(N__25628),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5 ));
    CascadeMux I__3444 (
            .O(N__25623),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_i6_3_cascade_ ));
    InMux I__3443 (
            .O(N__25620),
            .I(N__25616));
    InMux I__3442 (
            .O(N__25619),
            .I(N__25613));
    LocalMux I__3441 (
            .O(N__25616),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2 ));
    LocalMux I__3440 (
            .O(N__25613),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2 ));
    CascadeMux I__3439 (
            .O(N__25608),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_ ));
    CascadeMux I__3438 (
            .O(N__25605),
            .I(N__25601));
    InMux I__3437 (
            .O(N__25604),
            .I(N__25598));
    InMux I__3436 (
            .O(N__25601),
            .I(N__25595));
    LocalMux I__3435 (
            .O(N__25598),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_5 ));
    LocalMux I__3434 (
            .O(N__25595),
            .I(\spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_5 ));
    InMux I__3433 (
            .O(N__25590),
            .I(N__25586));
    InMux I__3432 (
            .O(N__25589),
            .I(N__25583));
    LocalMux I__3431 (
            .O(N__25586),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3 ));
    LocalMux I__3430 (
            .O(N__25583),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3 ));
    CascadeMux I__3429 (
            .O(N__25578),
            .I(N__25575));
    InMux I__3428 (
            .O(N__25575),
            .I(N__25570));
    InMux I__3427 (
            .O(N__25574),
            .I(N__25567));
    InMux I__3426 (
            .O(N__25573),
            .I(N__25564));
    LocalMux I__3425 (
            .O(N__25570),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1 ));
    LocalMux I__3424 (
            .O(N__25567),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1 ));
    LocalMux I__3423 (
            .O(N__25564),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1 ));
    CascadeMux I__3422 (
            .O(N__25557),
            .I(N__25553));
    CascadeMux I__3421 (
            .O(N__25556),
            .I(N__25549));
    InMux I__3420 (
            .O(N__25553),
            .I(N__25546));
    InMux I__3419 (
            .O(N__25552),
            .I(N__25543));
    InMux I__3418 (
            .O(N__25549),
            .I(N__25540));
    LocalMux I__3417 (
            .O(N__25546),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0 ));
    LocalMux I__3416 (
            .O(N__25543),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0 ));
    LocalMux I__3415 (
            .O(N__25540),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0 ));
    InMux I__3414 (
            .O(N__25533),
            .I(N__25529));
    InMux I__3413 (
            .O(N__25532),
            .I(N__25526));
    LocalMux I__3412 (
            .O(N__25529),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4 ));
    LocalMux I__3411 (
            .O(N__25526),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4 ));
    CascadeMux I__3410 (
            .O(N__25521),
            .I(\spi_slave_inst.un23_i_ssn_3_cascade_ ));
    InMux I__3409 (
            .O(N__25518),
            .I(N__25509));
    InMux I__3408 (
            .O(N__25517),
            .I(N__25509));
    InMux I__3407 (
            .O(N__25516),
            .I(N__25509));
    LocalMux I__3406 (
            .O(N__25509),
            .I(\spi_slave_inst.un23_i_ssn ));
    CascadeMux I__3405 (
            .O(N__25506),
            .I(\spi_slave_inst.un23_i_ssn_cascade_ ));
    CascadeMux I__3404 (
            .O(N__25503),
            .I(N__25499));
    InMux I__3403 (
            .O(N__25502),
            .I(N__25496));
    InMux I__3402 (
            .O(N__25499),
            .I(N__25493));
    LocalMux I__3401 (
            .O(N__25496),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa ));
    LocalMux I__3400 (
            .O(N__25493),
            .I(\spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa ));
    InMux I__3399 (
            .O(N__25488),
            .I(N__25485));
    LocalMux I__3398 (
            .O(N__25485),
            .I(N__25482));
    Span4Mux_h I__3397 (
            .O(N__25482),
            .I(N__25479));
    Span4Mux_h I__3396 (
            .O(N__25479),
            .I(N__25476));
    Odrv4 I__3395 (
            .O(N__25476),
            .I(op_gt_op_gt_un13_striginternallto23_8));
    InMux I__3394 (
            .O(N__25473),
            .I(bfn_9_20_0_));
    CEMux I__3393 (
            .O(N__25470),
            .I(N__25467));
    LocalMux I__3392 (
            .O(N__25467),
            .I(N__25464));
    Odrv4 I__3391 (
            .O(N__25464),
            .I(LED3_c_0));
    InMux I__3390 (
            .O(N__25461),
            .I(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0 ));
    InMux I__3389 (
            .O(N__25458),
            .I(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1 ));
    InMux I__3388 (
            .O(N__25455),
            .I(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2 ));
    CascadeMux I__3387 (
            .O(N__25452),
            .I(N__25449));
    InMux I__3386 (
            .O(N__25449),
            .I(N__25446));
    LocalMux I__3385 (
            .O(N__25446),
            .I(sEEDelayACQ_i_12));
    CascadeMux I__3384 (
            .O(N__25443),
            .I(N__25440));
    InMux I__3383 (
            .O(N__25440),
            .I(N__25437));
    LocalMux I__3382 (
            .O(N__25437),
            .I(sEEDelayACQ_i_13));
    CascadeMux I__3381 (
            .O(N__25434),
            .I(N__25431));
    InMux I__3380 (
            .O(N__25431),
            .I(N__25428));
    LocalMux I__3379 (
            .O(N__25428),
            .I(sEEDelayACQ_i_14));
    InMux I__3378 (
            .O(N__25425),
            .I(N__25422));
    LocalMux I__3377 (
            .O(N__25422),
            .I(sEEDelayACQ_i_15));
    CascadeMux I__3376 (
            .O(N__25419),
            .I(N__25416));
    InMux I__3375 (
            .O(N__25416),
            .I(N__25413));
    LocalMux I__3374 (
            .O(N__25413),
            .I(sEEDelayACQ_i_4));
    CascadeMux I__3373 (
            .O(N__25410),
            .I(N__25407));
    InMux I__3372 (
            .O(N__25407),
            .I(N__25404));
    LocalMux I__3371 (
            .O(N__25404),
            .I(sEEDelayACQ_i_5));
    CascadeMux I__3370 (
            .O(N__25401),
            .I(N__25398));
    InMux I__3369 (
            .O(N__25398),
            .I(N__25395));
    LocalMux I__3368 (
            .O(N__25395),
            .I(sEEDelayACQ_i_6));
    InMux I__3367 (
            .O(N__25392),
            .I(N__25389));
    LocalMux I__3366 (
            .O(N__25389),
            .I(sEEDelayACQ_i_7));
    CascadeMux I__3365 (
            .O(N__25386),
            .I(N__25383));
    InMux I__3364 (
            .O(N__25383),
            .I(N__25380));
    LocalMux I__3363 (
            .O(N__25380),
            .I(sEEDelayACQ_i_8));
    CascadeMux I__3362 (
            .O(N__25377),
            .I(N__25374));
    InMux I__3361 (
            .O(N__25374),
            .I(N__25371));
    LocalMux I__3360 (
            .O(N__25371),
            .I(sEEDelayACQ_i_9));
    CascadeMux I__3359 (
            .O(N__25368),
            .I(N__25365));
    InMux I__3358 (
            .O(N__25365),
            .I(N__25362));
    LocalMux I__3357 (
            .O(N__25362),
            .I(sEEDelayACQ_i_10));
    CascadeMux I__3356 (
            .O(N__25359),
            .I(N__25356));
    InMux I__3355 (
            .O(N__25356),
            .I(N__25353));
    LocalMux I__3354 (
            .O(N__25353),
            .I(sEEDelayACQ_i_11));
    InMux I__3353 (
            .O(N__25350),
            .I(N__25347));
    LocalMux I__3352 (
            .O(N__25347),
            .I(N__25344));
    Span4Mux_v I__3351 (
            .O(N__25344),
            .I(N__25341));
    Odrv4 I__3350 (
            .O(N__25341),
            .I(un4_spoff_cry_23_THRU_CO));
    InMux I__3349 (
            .O(N__25338),
            .I(bfn_9_16_0_));
    IoInMux I__3348 (
            .O(N__25335),
            .I(N__25332));
    LocalMux I__3347 (
            .O(N__25332),
            .I(N__25329));
    Span12Mux_s8_h I__3346 (
            .O(N__25329),
            .I(N__25326));
    Odrv12 I__3345 (
            .O(N__25326),
            .I(N_1612_i));
    InMux I__3344 (
            .O(N__25323),
            .I(N__25319));
    InMux I__3343 (
            .O(N__25322),
            .I(N__25316));
    LocalMux I__3342 (
            .O(N__25319),
            .I(N__25311));
    LocalMux I__3341 (
            .O(N__25316),
            .I(N__25311));
    Odrv4 I__3340 (
            .O(N__25311),
            .I(sCounterRAMZ0Z_6));
    InMux I__3339 (
            .O(N__25308),
            .I(N__25304));
    InMux I__3338 (
            .O(N__25307),
            .I(N__25301));
    LocalMux I__3337 (
            .O(N__25304),
            .I(N__25298));
    LocalMux I__3336 (
            .O(N__25301),
            .I(sCounterRAMZ0Z_3));
    Odrv4 I__3335 (
            .O(N__25298),
            .I(sCounterRAMZ0Z_3));
    InMux I__3334 (
            .O(N__25293),
            .I(N__25290));
    LocalMux I__3333 (
            .O(N__25290),
            .I(N__25287));
    Span4Mux_v I__3332 (
            .O(N__25287),
            .I(N__25283));
    InMux I__3331 (
            .O(N__25286),
            .I(N__25280));
    Odrv4 I__3330 (
            .O(N__25283),
            .I(button_debounce_counterZ0Z_21));
    LocalMux I__3329 (
            .O(N__25280),
            .I(button_debounce_counterZ0Z_21));
    CascadeMux I__3328 (
            .O(N__25275),
            .I(N__25272));
    InMux I__3327 (
            .O(N__25272),
            .I(N__25269));
    LocalMux I__3326 (
            .O(N__25269),
            .I(N__25266));
    Span4Mux_v I__3325 (
            .O(N__25266),
            .I(N__25262));
    InMux I__3324 (
            .O(N__25265),
            .I(N__25259));
    Odrv4 I__3323 (
            .O(N__25262),
            .I(button_debounce_counterZ0Z_22));
    LocalMux I__3322 (
            .O(N__25259),
            .I(button_debounce_counterZ0Z_22));
    InMux I__3321 (
            .O(N__25254),
            .I(N__25251));
    LocalMux I__3320 (
            .O(N__25251),
            .I(sbuttonModeStatus_0_sqmuxa_0));
    InMux I__3319 (
            .O(N__25248),
            .I(N__25245));
    LocalMux I__3318 (
            .O(N__25245),
            .I(N__25242));
    Span4Mux_h I__3317 (
            .O(N__25242),
            .I(N__25239));
    Odrv4 I__3316 (
            .O(N__25239),
            .I(sbuttonModeStatus_0_sqmuxa_18));
    InMux I__3315 (
            .O(N__25236),
            .I(N__25232));
    InMux I__3314 (
            .O(N__25235),
            .I(N__25229));
    LocalMux I__3313 (
            .O(N__25232),
            .I(button_debounce_counterZ0Z_4));
    LocalMux I__3312 (
            .O(N__25229),
            .I(button_debounce_counterZ0Z_4));
    InMux I__3311 (
            .O(N__25224),
            .I(N__25220));
    InMux I__3310 (
            .O(N__25223),
            .I(N__25217));
    LocalMux I__3309 (
            .O(N__25220),
            .I(button_debounce_counterZ0Z_3));
    LocalMux I__3308 (
            .O(N__25217),
            .I(button_debounce_counterZ0Z_3));
    CascadeMux I__3307 (
            .O(N__25212),
            .I(N__25208));
    InMux I__3306 (
            .O(N__25211),
            .I(N__25205));
    InMux I__3305 (
            .O(N__25208),
            .I(N__25202));
    LocalMux I__3304 (
            .O(N__25205),
            .I(button_debounce_counterZ0Z_5));
    LocalMux I__3303 (
            .O(N__25202),
            .I(button_debounce_counterZ0Z_5));
    InMux I__3302 (
            .O(N__25197),
            .I(N__25193));
    InMux I__3301 (
            .O(N__25196),
            .I(N__25190));
    LocalMux I__3300 (
            .O(N__25193),
            .I(button_debounce_counterZ0Z_2));
    LocalMux I__3299 (
            .O(N__25190),
            .I(button_debounce_counterZ0Z_2));
    InMux I__3298 (
            .O(N__25185),
            .I(N__25182));
    LocalMux I__3297 (
            .O(N__25182),
            .I(N__25179));
    Span4Mux_h I__3296 (
            .O(N__25179),
            .I(N__25176));
    Odrv4 I__3295 (
            .O(N__25176),
            .I(sbuttonModeStatus_0_sqmuxa_13));
    CascadeMux I__3294 (
            .O(N__25173),
            .I(N__25170));
    InMux I__3293 (
            .O(N__25170),
            .I(N__25167));
    LocalMux I__3292 (
            .O(N__25167),
            .I(sEEDelayACQ_i_0));
    CascadeMux I__3291 (
            .O(N__25164),
            .I(N__25161));
    InMux I__3290 (
            .O(N__25161),
            .I(N__25158));
    LocalMux I__3289 (
            .O(N__25158),
            .I(sEEDelayACQ_i_1));
    CascadeMux I__3288 (
            .O(N__25155),
            .I(N__25152));
    InMux I__3287 (
            .O(N__25152),
            .I(N__25149));
    LocalMux I__3286 (
            .O(N__25149),
            .I(sEEDelayACQ_i_2));
    CascadeMux I__3285 (
            .O(N__25146),
            .I(N__25143));
    InMux I__3284 (
            .O(N__25143),
            .I(N__25140));
    LocalMux I__3283 (
            .O(N__25140),
            .I(sEEDelayACQ_i_3));
    InMux I__3282 (
            .O(N__25137),
            .I(N__25134));
    LocalMux I__3281 (
            .O(N__25134),
            .I(sCounter_i_16));
    InMux I__3280 (
            .O(N__25131),
            .I(N__25128));
    LocalMux I__3279 (
            .O(N__25128),
            .I(sCounter_i_17));
    InMux I__3278 (
            .O(N__25125),
            .I(N__25122));
    LocalMux I__3277 (
            .O(N__25122),
            .I(sCounter_i_18));
    InMux I__3276 (
            .O(N__25119),
            .I(N__25116));
    LocalMux I__3275 (
            .O(N__25116),
            .I(sCounter_i_19));
    InMux I__3274 (
            .O(N__25113),
            .I(N__25110));
    LocalMux I__3273 (
            .O(N__25110),
            .I(sCounter_i_20));
    InMux I__3272 (
            .O(N__25107),
            .I(N__25104));
    LocalMux I__3271 (
            .O(N__25104),
            .I(sCounter_i_21));
    InMux I__3270 (
            .O(N__25101),
            .I(N__25098));
    LocalMux I__3269 (
            .O(N__25098),
            .I(sCounter_i_22));
    InMux I__3268 (
            .O(N__25095),
            .I(N__25092));
    LocalMux I__3267 (
            .O(N__25092),
            .I(sCounter_i_23));
    CascadeMux I__3266 (
            .O(N__25089),
            .I(un1_reset_rpi_inv_2_i_1_cascade_));
    InMux I__3265 (
            .O(N__25086),
            .I(N__25083));
    LocalMux I__3264 (
            .O(N__25083),
            .I(N__25080));
    Odrv4 I__3263 (
            .O(N__25080),
            .I(un1_sTrigCounter_ac0_0_4));
    InMux I__3262 (
            .O(N__25077),
            .I(N__25072));
    InMux I__3261 (
            .O(N__25076),
            .I(N__25069));
    InMux I__3260 (
            .O(N__25075),
            .I(N__25066));
    LocalMux I__3259 (
            .O(N__25072),
            .I(N__25061));
    LocalMux I__3258 (
            .O(N__25069),
            .I(N__25061));
    LocalMux I__3257 (
            .O(N__25066),
            .I(sTrigCounterZ0Z_6));
    Odrv12 I__3256 (
            .O(N__25061),
            .I(sTrigCounterZ0Z_6));
    InMux I__3255 (
            .O(N__25056),
            .I(N__25053));
    LocalMux I__3254 (
            .O(N__25053),
            .I(N__25050));
    Odrv4 I__3253 (
            .O(N__25050),
            .I(un1_sTrigCounter_axbxc7_m7_0_a2_2));
    InMux I__3252 (
            .O(N__25047),
            .I(N__25044));
    LocalMux I__3251 (
            .O(N__25044),
            .I(un1_reset_rpi_inv_2_i_1));
    InMux I__3250 (
            .O(N__25041),
            .I(N__25038));
    LocalMux I__3249 (
            .O(N__25038),
            .I(N__25035));
    Odrv4 I__3248 (
            .O(N__25035),
            .I(N_123));
    InMux I__3247 (
            .O(N__25032),
            .I(N__25028));
    CascadeMux I__3246 (
            .O(N__25031),
            .I(N__25025));
    LocalMux I__3245 (
            .O(N__25028),
            .I(N__25022));
    InMux I__3244 (
            .O(N__25025),
            .I(N__25019));
    Span4Mux_v I__3243 (
            .O(N__25022),
            .I(N__25016));
    LocalMux I__3242 (
            .O(N__25019),
            .I(sTrigCounterZ0Z_7));
    Odrv4 I__3241 (
            .O(N__25016),
            .I(sTrigCounterZ0Z_7));
    InMux I__3240 (
            .O(N__25011),
            .I(N__25008));
    LocalMux I__3239 (
            .O(N__25008),
            .I(sEEPeriodZ0Z_14));
    InMux I__3238 (
            .O(N__25005),
            .I(N__25002));
    LocalMux I__3237 (
            .O(N__25002),
            .I(sEEPeriodZ0Z_15));
    InMux I__3236 (
            .O(N__24999),
            .I(N__24996));
    LocalMux I__3235 (
            .O(N__24996),
            .I(sEEPeriodZ0Z_8));
    InMux I__3234 (
            .O(N__24993),
            .I(N__24990));
    LocalMux I__3233 (
            .O(N__24990),
            .I(sEEPeriodZ0Z_9));
    InMux I__3232 (
            .O(N__24987),
            .I(N__24984));
    LocalMux I__3231 (
            .O(N__24984),
            .I(N__24981));
    Span4Mux_v I__3230 (
            .O(N__24981),
            .I(N__24978));
    Span4Mux_h I__3229 (
            .O(N__24978),
            .I(N__24975));
    Odrv4 I__3228 (
            .O(N__24975),
            .I(op_gt_op_gt_un13_striginternallto23_12));
    InMux I__3227 (
            .O(N__24972),
            .I(N__24969));
    LocalMux I__3226 (
            .O(N__24969),
            .I(N__24966));
    Span4Mux_h I__3225 (
            .O(N__24966),
            .I(N__24963));
    Odrv4 I__3224 (
            .O(N__24963),
            .I(un1_reset_rpi_inv_2_i_o3_12));
    CascadeMux I__3223 (
            .O(N__24960),
            .I(N__24957));
    InMux I__3222 (
            .O(N__24957),
            .I(N__24954));
    LocalMux I__3221 (
            .O(N__24954),
            .I(N__24951));
    Span4Mux_h I__3220 (
            .O(N__24951),
            .I(N__24948));
    Odrv4 I__3219 (
            .O(N__24948),
            .I(op_gt_op_gt_un13_striginternallto23_15));
    CascadeMux I__3218 (
            .O(N__24945),
            .I(N__24935));
    InMux I__3217 (
            .O(N__24944),
            .I(N__24931));
    InMux I__3216 (
            .O(N__24943),
            .I(N__24928));
    InMux I__3215 (
            .O(N__24942),
            .I(N__24924));
    InMux I__3214 (
            .O(N__24941),
            .I(N__24921));
    CascadeMux I__3213 (
            .O(N__24940),
            .I(N__24918));
    CascadeMux I__3212 (
            .O(N__24939),
            .I(N__24915));
    CascadeMux I__3211 (
            .O(N__24938),
            .I(N__24912));
    InMux I__3210 (
            .O(N__24935),
            .I(N__24904));
    InMux I__3209 (
            .O(N__24934),
            .I(N__24904));
    LocalMux I__3208 (
            .O(N__24931),
            .I(N__24901));
    LocalMux I__3207 (
            .O(N__24928),
            .I(N__24898));
    InMux I__3206 (
            .O(N__24927),
            .I(N__24895));
    LocalMux I__3205 (
            .O(N__24924),
            .I(N__24890));
    LocalMux I__3204 (
            .O(N__24921),
            .I(N__24890));
    InMux I__3203 (
            .O(N__24918),
            .I(N__24879));
    InMux I__3202 (
            .O(N__24915),
            .I(N__24879));
    InMux I__3201 (
            .O(N__24912),
            .I(N__24879));
    InMux I__3200 (
            .O(N__24911),
            .I(N__24879));
    InMux I__3199 (
            .O(N__24910),
            .I(N__24879));
    CascadeMux I__3198 (
            .O(N__24909),
            .I(N__24875));
    LocalMux I__3197 (
            .O(N__24904),
            .I(N__24871));
    Span4Mux_v I__3196 (
            .O(N__24901),
            .I(N__24866));
    Span4Mux_v I__3195 (
            .O(N__24898),
            .I(N__24866));
    LocalMux I__3194 (
            .O(N__24895),
            .I(N__24859));
    Span4Mux_h I__3193 (
            .O(N__24890),
            .I(N__24859));
    LocalMux I__3192 (
            .O(N__24879),
            .I(N__24859));
    InMux I__3191 (
            .O(N__24878),
            .I(N__24852));
    InMux I__3190 (
            .O(N__24875),
            .I(N__24852));
    InMux I__3189 (
            .O(N__24874),
            .I(N__24852));
    Odrv4 I__3188 (
            .O(N__24871),
            .I(sEETrigInternal_prevZ0));
    Odrv4 I__3187 (
            .O(N__24866),
            .I(sEETrigInternal_prevZ0));
    Odrv4 I__3186 (
            .O(N__24859),
            .I(sEETrigInternal_prevZ0));
    LocalMux I__3185 (
            .O(N__24852),
            .I(sEETrigInternal_prevZ0));
    CascadeMux I__3184 (
            .O(N__24843),
            .I(N__24840));
    InMux I__3183 (
            .O(N__24840),
            .I(N__24837));
    LocalMux I__3182 (
            .O(N__24837),
            .I(N__24834));
    Span4Mux_h I__3181 (
            .O(N__24834),
            .I(N__24831));
    Span4Mux_v I__3180 (
            .O(N__24831),
            .I(N__24828));
    Odrv4 I__3179 (
            .O(N__24828),
            .I(N_5_0));
    InMux I__3178 (
            .O(N__24825),
            .I(N__24819));
    InMux I__3177 (
            .O(N__24824),
            .I(N__24811));
    InMux I__3176 (
            .O(N__24823),
            .I(N__24811));
    InMux I__3175 (
            .O(N__24822),
            .I(N__24808));
    LocalMux I__3174 (
            .O(N__24819),
            .I(N__24805));
    InMux I__3173 (
            .O(N__24818),
            .I(N__24800));
    InMux I__3172 (
            .O(N__24817),
            .I(N__24800));
    InMux I__3171 (
            .O(N__24816),
            .I(N__24794));
    LocalMux I__3170 (
            .O(N__24811),
            .I(N__24791));
    LocalMux I__3169 (
            .O(N__24808),
            .I(N__24787));
    Span4Mux_v I__3168 (
            .O(N__24805),
            .I(N__24782));
    LocalMux I__3167 (
            .O(N__24800),
            .I(N__24782));
    InMux I__3166 (
            .O(N__24799),
            .I(N__24779));
    InMux I__3165 (
            .O(N__24798),
            .I(N__24776));
    InMux I__3164 (
            .O(N__24797),
            .I(N__24773));
    LocalMux I__3163 (
            .O(N__24794),
            .I(N__24768));
    Span4Mux_v I__3162 (
            .O(N__24791),
            .I(N__24768));
    InMux I__3161 (
            .O(N__24790),
            .I(N__24765));
    Span4Mux_h I__3160 (
            .O(N__24787),
            .I(N__24758));
    Span4Mux_v I__3159 (
            .O(N__24782),
            .I(N__24758));
    LocalMux I__3158 (
            .O(N__24779),
            .I(N__24758));
    LocalMux I__3157 (
            .O(N__24776),
            .I(un4_speriod_cry_23_THRU_CO));
    LocalMux I__3156 (
            .O(N__24773),
            .I(un4_speriod_cry_23_THRU_CO));
    Odrv4 I__3155 (
            .O(N__24768),
            .I(un4_speriod_cry_23_THRU_CO));
    LocalMux I__3154 (
            .O(N__24765),
            .I(un4_speriod_cry_23_THRU_CO));
    Odrv4 I__3153 (
            .O(N__24758),
            .I(un4_speriod_cry_23_THRU_CO));
    CascadeMux I__3152 (
            .O(N__24747),
            .I(un1_reset_rpi_inv_2_i_1_1_0_cascade_));
    CascadeMux I__3151 (
            .O(N__24744),
            .I(un1_sTrigCounter_ac0_0_0_cascade_));
    InMux I__3150 (
            .O(N__24741),
            .I(N__24737));
    InMux I__3149 (
            .O(N__24740),
            .I(N__24734));
    LocalMux I__3148 (
            .O(N__24737),
            .I(N__24731));
    LocalMux I__3147 (
            .O(N__24734),
            .I(N__24726));
    Span4Mux_h I__3146 (
            .O(N__24731),
            .I(N__24726));
    Odrv4 I__3145 (
            .O(N__24726),
            .I(un1_reset_rpi_inv_2_i_o3_0_0));
    CascadeMux I__3144 (
            .O(N__24723),
            .I(un1_sTrigCounter_ac0_0_2_0_cascade_));
    InMux I__3143 (
            .O(N__24720),
            .I(N__24715));
    InMux I__3142 (
            .O(N__24719),
            .I(N__24710));
    InMux I__3141 (
            .O(N__24718),
            .I(N__24707));
    LocalMux I__3140 (
            .O(N__24715),
            .I(N__24704));
    CascadeMux I__3139 (
            .O(N__24714),
            .I(N__24700));
    CascadeMux I__3138 (
            .O(N__24713),
            .I(N__24695));
    LocalMux I__3137 (
            .O(N__24710),
            .I(N__24691));
    LocalMux I__3136 (
            .O(N__24707),
            .I(N__24686));
    Span4Mux_v I__3135 (
            .O(N__24704),
            .I(N__24686));
    InMux I__3134 (
            .O(N__24703),
            .I(N__24683));
    InMux I__3133 (
            .O(N__24700),
            .I(N__24680));
    InMux I__3132 (
            .O(N__24699),
            .I(N__24677));
    InMux I__3131 (
            .O(N__24698),
            .I(N__24674));
    InMux I__3130 (
            .O(N__24695),
            .I(N__24669));
    InMux I__3129 (
            .O(N__24694),
            .I(N__24669));
    Span4Mux_v I__3128 (
            .O(N__24691),
            .I(N__24664));
    Span4Mux_v I__3127 (
            .O(N__24686),
            .I(N__24664));
    LocalMux I__3126 (
            .O(N__24683),
            .I(un10_trig_prev_cry_7_THRU_CO));
    LocalMux I__3125 (
            .O(N__24680),
            .I(un10_trig_prev_cry_7_THRU_CO));
    LocalMux I__3124 (
            .O(N__24677),
            .I(un10_trig_prev_cry_7_THRU_CO));
    LocalMux I__3123 (
            .O(N__24674),
            .I(un10_trig_prev_cry_7_THRU_CO));
    LocalMux I__3122 (
            .O(N__24669),
            .I(un10_trig_prev_cry_7_THRU_CO));
    Odrv4 I__3121 (
            .O(N__24664),
            .I(un10_trig_prev_cry_7_THRU_CO));
    InMux I__3120 (
            .O(N__24651),
            .I(N__24648));
    LocalMux I__3119 (
            .O(N__24648),
            .I(N__24642));
    InMux I__3118 (
            .O(N__24647),
            .I(N__24637));
    InMux I__3117 (
            .O(N__24646),
            .I(N__24637));
    InMux I__3116 (
            .O(N__24645),
            .I(N__24634));
    Odrv4 I__3115 (
            .O(N__24642),
            .I(sTrigCounterZ0Z_5));
    LocalMux I__3114 (
            .O(N__24637),
            .I(sTrigCounterZ0Z_5));
    LocalMux I__3113 (
            .O(N__24634),
            .I(sTrigCounterZ0Z_5));
    InMux I__3112 (
            .O(N__24627),
            .I(N__24621));
    InMux I__3111 (
            .O(N__24626),
            .I(N__24621));
    LocalMux I__3110 (
            .O(N__24621),
            .I(un1_sTrigCounter_ac0_0_2));
    CascadeMux I__3109 (
            .O(N__24618),
            .I(un1_sTrigCounter_ac0_3_out_cascade_));
    InMux I__3108 (
            .O(N__24615),
            .I(N__24603));
    InMux I__3107 (
            .O(N__24614),
            .I(N__24603));
    InMux I__3106 (
            .O(N__24613),
            .I(N__24603));
    InMux I__3105 (
            .O(N__24612),
            .I(N__24599));
    InMux I__3104 (
            .O(N__24611),
            .I(N__24594));
    InMux I__3103 (
            .O(N__24610),
            .I(N__24594));
    LocalMux I__3102 (
            .O(N__24603),
            .I(N__24591));
    InMux I__3101 (
            .O(N__24602),
            .I(N__24588));
    LocalMux I__3100 (
            .O(N__24599),
            .I(N__24585));
    LocalMux I__3099 (
            .O(N__24594),
            .I(sTrigCounterZ0Z_2));
    Odrv4 I__3098 (
            .O(N__24591),
            .I(sTrigCounterZ0Z_2));
    LocalMux I__3097 (
            .O(N__24588),
            .I(sTrigCounterZ0Z_2));
    Odrv4 I__3096 (
            .O(N__24585),
            .I(sTrigCounterZ0Z_2));
    CascadeMux I__3095 (
            .O(N__24576),
            .I(N__24573));
    InMux I__3094 (
            .O(N__24573),
            .I(N__24570));
    LocalMux I__3093 (
            .O(N__24570),
            .I(g1_0_1_0));
    InMux I__3092 (
            .O(N__24567),
            .I(N__24564));
    LocalMux I__3091 (
            .O(N__24564),
            .I(g1_3_0));
    InMux I__3090 (
            .O(N__24561),
            .I(N__24558));
    LocalMux I__3089 (
            .O(N__24558),
            .I(sEEPeriodZ0Z_10));
    InMux I__3088 (
            .O(N__24555),
            .I(N__24552));
    LocalMux I__3087 (
            .O(N__24552),
            .I(sEEPeriodZ0Z_11));
    InMux I__3086 (
            .O(N__24549),
            .I(N__24546));
    LocalMux I__3085 (
            .O(N__24546),
            .I(sEEPeriodZ0Z_12));
    InMux I__3084 (
            .O(N__24543),
            .I(N__24540));
    LocalMux I__3083 (
            .O(N__24540),
            .I(sEEPeriodZ0Z_13));
    CascadeMux I__3082 (
            .O(N__24537),
            .I(N__24534));
    InMux I__3081 (
            .O(N__24534),
            .I(N__24531));
    LocalMux I__3080 (
            .O(N__24531),
            .I(un10_trig_prev_7));
    InMux I__3079 (
            .O(N__24528),
            .I(N__24525));
    LocalMux I__3078 (
            .O(N__24525),
            .I(sTrigCounter_i_7));
    InMux I__3077 (
            .O(N__24522),
            .I(bfn_9_9_0_));
    CEMux I__3076 (
            .O(N__24519),
            .I(N__24516));
    LocalMux I__3075 (
            .O(N__24516),
            .I(N__24513));
    Odrv4 I__3074 (
            .O(N__24513),
            .I(sAddress_RNI9IH12_1Z0Z_1));
    InMux I__3073 (
            .O(N__24510),
            .I(N__24503));
    InMux I__3072 (
            .O(N__24509),
            .I(N__24498));
    InMux I__3071 (
            .O(N__24508),
            .I(N__24498));
    InMux I__3070 (
            .O(N__24507),
            .I(N__24495));
    InMux I__3069 (
            .O(N__24506),
            .I(N__24492));
    LocalMux I__3068 (
            .O(N__24503),
            .I(N__24485));
    LocalMux I__3067 (
            .O(N__24498),
            .I(N__24482));
    LocalMux I__3066 (
            .O(N__24495),
            .I(N__24477));
    LocalMux I__3065 (
            .O(N__24492),
            .I(N__24477));
    InMux I__3064 (
            .O(N__24491),
            .I(N__24470));
    InMux I__3063 (
            .O(N__24490),
            .I(N__24470));
    InMux I__3062 (
            .O(N__24489),
            .I(N__24470));
    InMux I__3061 (
            .O(N__24488),
            .I(N__24461));
    Span4Mux_v I__3060 (
            .O(N__24485),
            .I(N__24458));
    Span4Mux_v I__3059 (
            .O(N__24482),
            .I(N__24451));
    Span4Mux_h I__3058 (
            .O(N__24477),
            .I(N__24451));
    LocalMux I__3057 (
            .O(N__24470),
            .I(N__24451));
    InMux I__3056 (
            .O(N__24469),
            .I(N__24438));
    InMux I__3055 (
            .O(N__24468),
            .I(N__24438));
    InMux I__3054 (
            .O(N__24467),
            .I(N__24438));
    InMux I__3053 (
            .O(N__24466),
            .I(N__24438));
    InMux I__3052 (
            .O(N__24465),
            .I(N__24438));
    InMux I__3051 (
            .O(N__24464),
            .I(N__24438));
    LocalMux I__3050 (
            .O(N__24461),
            .I(trig_prevZ0));
    Odrv4 I__3049 (
            .O(N__24458),
            .I(trig_prevZ0));
    Odrv4 I__3048 (
            .O(N__24451),
            .I(trig_prevZ0));
    LocalMux I__3047 (
            .O(N__24438),
            .I(trig_prevZ0));
    InMux I__3046 (
            .O(N__24429),
            .I(N__24425));
    CascadeMux I__3045 (
            .O(N__24428),
            .I(N__24422));
    LocalMux I__3044 (
            .O(N__24425),
            .I(N__24419));
    InMux I__3043 (
            .O(N__24422),
            .I(N__24416));
    Span4Mux_v I__3042 (
            .O(N__24419),
            .I(N__24413));
    LocalMux I__3041 (
            .O(N__24416),
            .I(N__24410));
    Odrv4 I__3040 (
            .O(N__24413),
            .I(un3_trig_0_3));
    Odrv4 I__3039 (
            .O(N__24410),
            .I(un3_trig_0_3));
    InMux I__3038 (
            .O(N__24405),
            .I(N__24402));
    LocalMux I__3037 (
            .O(N__24402),
            .I(g1_0_0_2));
    InMux I__3036 (
            .O(N__24399),
            .I(N__24396));
    LocalMux I__3035 (
            .O(N__24396),
            .I(N__24393));
    Odrv4 I__3034 (
            .O(N__24393),
            .I(g1_0_0));
    InMux I__3033 (
            .O(N__24390),
            .I(N__24387));
    LocalMux I__3032 (
            .O(N__24387),
            .I(g1_0));
    InMux I__3031 (
            .O(N__24384),
            .I(N__24381));
    LocalMux I__3030 (
            .O(N__24381),
            .I(N__24373));
    InMux I__3029 (
            .O(N__24380),
            .I(N__24370));
    InMux I__3028 (
            .O(N__24379),
            .I(N__24365));
    InMux I__3027 (
            .O(N__24378),
            .I(N__24365));
    InMux I__3026 (
            .O(N__24377),
            .I(N__24362));
    CascadeMux I__3025 (
            .O(N__24376),
            .I(N__24358));
    Span4Mux_v I__3024 (
            .O(N__24373),
            .I(N__24352));
    LocalMux I__3023 (
            .O(N__24370),
            .I(N__24352));
    LocalMux I__3022 (
            .O(N__24365),
            .I(N__24347));
    LocalMux I__3021 (
            .O(N__24362),
            .I(N__24347));
    InMux I__3020 (
            .O(N__24361),
            .I(N__24344));
    InMux I__3019 (
            .O(N__24358),
            .I(N__24339));
    InMux I__3018 (
            .O(N__24357),
            .I(N__24339));
    Span4Mux_v I__3017 (
            .O(N__24352),
            .I(N__24332));
    Span4Mux_h I__3016 (
            .O(N__24347),
            .I(N__24332));
    LocalMux I__3015 (
            .O(N__24344),
            .I(N__24332));
    LocalMux I__3014 (
            .O(N__24339),
            .I(N__24329));
    Span4Mux_v I__3013 (
            .O(N__24332),
            .I(N__24326));
    Odrv12 I__3012 (
            .O(N__24329),
            .I(sPeriod_prevZ0));
    Odrv4 I__3011 (
            .O(N__24326),
            .I(sPeriod_prevZ0));
    IoInMux I__3010 (
            .O(N__24321),
            .I(N__24318));
    LocalMux I__3009 (
            .O(N__24318),
            .I(N__24315));
    Span4Mux_s1_h I__3008 (
            .O(N__24315),
            .I(N__24311));
    CascadeMux I__3007 (
            .O(N__24314),
            .I(N__24306));
    Span4Mux_h I__3006 (
            .O(N__24311),
            .I(N__24303));
    CascadeMux I__3005 (
            .O(N__24310),
            .I(N__24300));
    CascadeMux I__3004 (
            .O(N__24309),
            .I(N__24297));
    InMux I__3003 (
            .O(N__24306),
            .I(N__24294));
    Span4Mux_h I__3002 (
            .O(N__24303),
            .I(N__24291));
    InMux I__3001 (
            .O(N__24300),
            .I(N__24288));
    InMux I__3000 (
            .O(N__24297),
            .I(N__24285));
    LocalMux I__2999 (
            .O(N__24294),
            .I(N__24282));
    Span4Mux_v I__2998 (
            .O(N__24291),
            .I(N__24277));
    LocalMux I__2997 (
            .O(N__24288),
            .I(N__24277));
    LocalMux I__2996 (
            .O(N__24285),
            .I(N__24274));
    Span4Mux_h I__2995 (
            .O(N__24282),
            .I(N__24265));
    Span4Mux_v I__2994 (
            .O(N__24277),
            .I(N__24265));
    Span4Mux_h I__2993 (
            .O(N__24274),
            .I(N__24265));
    InMux I__2992 (
            .O(N__24273),
            .I(N__24260));
    InMux I__2991 (
            .O(N__24272),
            .I(N__24260));
    Span4Mux_v I__2990 (
            .O(N__24265),
            .I(N__24252));
    LocalMux I__2989 (
            .O(N__24260),
            .I(N__24252));
    InMux I__2988 (
            .O(N__24259),
            .I(N__24247));
    InMux I__2987 (
            .O(N__24258),
            .I(N__24247));
    InMux I__2986 (
            .O(N__24257),
            .I(N__24244));
    Span4Mux_h I__2985 (
            .O(N__24252),
            .I(N__24241));
    LocalMux I__2984 (
            .O(N__24247),
            .I(N__24236));
    LocalMux I__2983 (
            .O(N__24244),
            .I(N__24236));
    Odrv4 I__2982 (
            .O(N__24241),
            .I(LED_MODE_c));
    Odrv12 I__2981 (
            .O(N__24236),
            .I(LED_MODE_c));
    InMux I__2980 (
            .O(N__24231),
            .I(N__24225));
    InMux I__2979 (
            .O(N__24230),
            .I(N__24222));
    InMux I__2978 (
            .O(N__24229),
            .I(N__24219));
    InMux I__2977 (
            .O(N__24228),
            .I(N__24216));
    LocalMux I__2976 (
            .O(N__24225),
            .I(N__24213));
    LocalMux I__2975 (
            .O(N__24222),
            .I(sTrigCounterZ0Z_4));
    LocalMux I__2974 (
            .O(N__24219),
            .I(sTrigCounterZ0Z_4));
    LocalMux I__2973 (
            .O(N__24216),
            .I(sTrigCounterZ0Z_4));
    Odrv4 I__2972 (
            .O(N__24213),
            .I(sTrigCounterZ0Z_4));
    InMux I__2971 (
            .O(N__24204),
            .I(N__24197));
    InMux I__2970 (
            .O(N__24203),
            .I(N__24194));
    InMux I__2969 (
            .O(N__24202),
            .I(N__24189));
    InMux I__2968 (
            .O(N__24201),
            .I(N__24189));
    InMux I__2967 (
            .O(N__24200),
            .I(N__24186));
    LocalMux I__2966 (
            .O(N__24197),
            .I(sTrigCounterZ0Z_3));
    LocalMux I__2965 (
            .O(N__24194),
            .I(sTrigCounterZ0Z_3));
    LocalMux I__2964 (
            .O(N__24189),
            .I(sTrigCounterZ0Z_3));
    LocalMux I__2963 (
            .O(N__24186),
            .I(sTrigCounterZ0Z_3));
    CascadeMux I__2962 (
            .O(N__24177),
            .I(N__24173));
    InMux I__2961 (
            .O(N__24176),
            .I(N__24168));
    InMux I__2960 (
            .O(N__24173),
            .I(N__24168));
    LocalMux I__2959 (
            .O(N__24168),
            .I(sEETrigCounterZ0Z_4));
    CascadeMux I__2958 (
            .O(N__24165),
            .I(N__24160));
    InMux I__2957 (
            .O(N__24164),
            .I(N__24155));
    InMux I__2956 (
            .O(N__24163),
            .I(N__24155));
    InMux I__2955 (
            .O(N__24160),
            .I(N__24152));
    LocalMux I__2954 (
            .O(N__24155),
            .I(un8_trig_prev_0_c5_a0_0));
    LocalMux I__2953 (
            .O(N__24152),
            .I(un8_trig_prev_0_c5_a0_0));
    InMux I__2952 (
            .O(N__24147),
            .I(N__24144));
    LocalMux I__2951 (
            .O(N__24144),
            .I(sTrigCounter_i_0));
    InMux I__2950 (
            .O(N__24141),
            .I(N__24138));
    LocalMux I__2949 (
            .O(N__24138),
            .I(sTrigCounter_i_1));
    CascadeMux I__2948 (
            .O(N__24135),
            .I(N__24132));
    InMux I__2947 (
            .O(N__24132),
            .I(N__24129));
    LocalMux I__2946 (
            .O(N__24129),
            .I(sTrigCounter_i_2));
    InMux I__2945 (
            .O(N__24126),
            .I(N__24123));
    LocalMux I__2944 (
            .O(N__24123),
            .I(sTrigCounter_i_3));
    CascadeMux I__2943 (
            .O(N__24120),
            .I(N__24117));
    InMux I__2942 (
            .O(N__24117),
            .I(N__24114));
    LocalMux I__2941 (
            .O(N__24114),
            .I(un10_trig_prev_4));
    InMux I__2940 (
            .O(N__24111),
            .I(N__24108));
    LocalMux I__2939 (
            .O(N__24108),
            .I(sTrigCounter_i_4));
    CascadeMux I__2938 (
            .O(N__24105),
            .I(N__24102));
    InMux I__2937 (
            .O(N__24102),
            .I(N__24099));
    LocalMux I__2936 (
            .O(N__24099),
            .I(un10_trig_prev_5));
    InMux I__2935 (
            .O(N__24096),
            .I(N__24093));
    LocalMux I__2934 (
            .O(N__24093),
            .I(sTrigCounter_i_5));
    CascadeMux I__2933 (
            .O(N__24090),
            .I(N__24087));
    InMux I__2932 (
            .O(N__24087),
            .I(N__24084));
    LocalMux I__2931 (
            .O(N__24084),
            .I(un10_trig_prev_6));
    InMux I__2930 (
            .O(N__24081),
            .I(N__24078));
    LocalMux I__2929 (
            .O(N__24078),
            .I(N__24075));
    Odrv4 I__2928 (
            .O(N__24075),
            .I(sTrigCounter_i_6));
    InMux I__2927 (
            .O(N__24072),
            .I(N__24069));
    LocalMux I__2926 (
            .O(N__24069),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2 ));
    InMux I__2925 (
            .O(N__24066),
            .I(N__24060));
    InMux I__2924 (
            .O(N__24065),
            .I(N__24060));
    LocalMux I__2923 (
            .O(N__24060),
            .I(N__24053));
    InMux I__2922 (
            .O(N__24059),
            .I(N__24048));
    InMux I__2921 (
            .O(N__24058),
            .I(N__24048));
    InMux I__2920 (
            .O(N__24057),
            .I(N__24045));
    CascadeMux I__2919 (
            .O(N__24056),
            .I(N__24042));
    Span4Mux_h I__2918 (
            .O(N__24053),
            .I(N__24033));
    LocalMux I__2917 (
            .O(N__24048),
            .I(N__24033));
    LocalMux I__2916 (
            .O(N__24045),
            .I(N__24033));
    InMux I__2915 (
            .O(N__24042),
            .I(N__24028));
    InMux I__2914 (
            .O(N__24041),
            .I(N__24028));
    InMux I__2913 (
            .O(N__24040),
            .I(N__24025));
    Span4Mux_v I__2912 (
            .O(N__24033),
            .I(N__24021));
    LocalMux I__2911 (
            .O(N__24028),
            .I(N__24018));
    LocalMux I__2910 (
            .O(N__24025),
            .I(N__24015));
    InMux I__2909 (
            .O(N__24024),
            .I(N__24012));
    Span4Mux_v I__2908 (
            .O(N__24021),
            .I(N__24009));
    Span4Mux_v I__2907 (
            .O(N__24018),
            .I(N__24006));
    Span4Mux_v I__2906 (
            .O(N__24015),
            .I(N__24001));
    LocalMux I__2905 (
            .O(N__24012),
            .I(N__24001));
    Span4Mux_h I__2904 (
            .O(N__24009),
            .I(N__23998));
    Span4Mux_v I__2903 (
            .O(N__24006),
            .I(N__23995));
    Span4Mux_h I__2902 (
            .O(N__24001),
            .I(N__23992));
    Sp12to4 I__2901 (
            .O(N__23998),
            .I(N__23987));
    Sp12to4 I__2900 (
            .O(N__23995),
            .I(N__23987));
    Span4Mux_v I__2899 (
            .O(N__23992),
            .I(N__23984));
    Odrv12 I__2898 (
            .O(N__23987),
            .I(trig_ext_c));
    Odrv4 I__2897 (
            .O(N__23984),
            .I(trig_ext_c));
    InMux I__2896 (
            .O(N__23979),
            .I(N__23973));
    InMux I__2895 (
            .O(N__23978),
            .I(N__23973));
    LocalMux I__2894 (
            .O(N__23973),
            .I(N__23967));
    InMux I__2893 (
            .O(N__23972),
            .I(N__23959));
    InMux I__2892 (
            .O(N__23971),
            .I(N__23959));
    InMux I__2891 (
            .O(N__23970),
            .I(N__23956));
    Span4Mux_h I__2890 (
            .O(N__23967),
            .I(N__23953));
    InMux I__2889 (
            .O(N__23966),
            .I(N__23948));
    InMux I__2888 (
            .O(N__23965),
            .I(N__23948));
    InMux I__2887 (
            .O(N__23964),
            .I(N__23945));
    LocalMux I__2886 (
            .O(N__23959),
            .I(N__23940));
    LocalMux I__2885 (
            .O(N__23956),
            .I(N__23940));
    Span4Mux_h I__2884 (
            .O(N__23953),
            .I(N__23935));
    LocalMux I__2883 (
            .O(N__23948),
            .I(N__23935));
    LocalMux I__2882 (
            .O(N__23945),
            .I(N__23932));
    Span4Mux_v I__2881 (
            .O(N__23940),
            .I(N__23928));
    Span4Mux_v I__2880 (
            .O(N__23935),
            .I(N__23925));
    Span4Mux_v I__2879 (
            .O(N__23932),
            .I(N__23922));
    InMux I__2878 (
            .O(N__23931),
            .I(N__23919));
    Sp12to4 I__2877 (
            .O(N__23928),
            .I(N__23910));
    Sp12to4 I__2876 (
            .O(N__23925),
            .I(N__23910));
    Sp12to4 I__2875 (
            .O(N__23922),
            .I(N__23910));
    LocalMux I__2874 (
            .O(N__23919),
            .I(N__23910));
    Odrv12 I__2873 (
            .O(N__23910),
            .I(trig_rpi_c));
    InMux I__2872 (
            .O(N__23907),
            .I(N__23903));
    CascadeMux I__2871 (
            .O(N__23906),
            .I(N__23896));
    LocalMux I__2870 (
            .O(N__23903),
            .I(N__23893));
    InMux I__2869 (
            .O(N__23902),
            .I(N__23887));
    InMux I__2868 (
            .O(N__23901),
            .I(N__23887));
    InMux I__2867 (
            .O(N__23900),
            .I(N__23884));
    InMux I__2866 (
            .O(N__23899),
            .I(N__23879));
    InMux I__2865 (
            .O(N__23896),
            .I(N__23879));
    Span4Mux_v I__2864 (
            .O(N__23893),
            .I(N__23874));
    InMux I__2863 (
            .O(N__23892),
            .I(N__23871));
    LocalMux I__2862 (
            .O(N__23887),
            .I(N__23864));
    LocalMux I__2861 (
            .O(N__23884),
            .I(N__23864));
    LocalMux I__2860 (
            .O(N__23879),
            .I(N__23864));
    InMux I__2859 (
            .O(N__23878),
            .I(N__23859));
    InMux I__2858 (
            .O(N__23877),
            .I(N__23859));
    Span4Mux_h I__2857 (
            .O(N__23874),
            .I(N__23856));
    LocalMux I__2856 (
            .O(N__23871),
            .I(N__23853));
    Span4Mux_h I__2855 (
            .O(N__23864),
            .I(N__23848));
    LocalMux I__2854 (
            .O(N__23859),
            .I(N__23848));
    Sp12to4 I__2853 (
            .O(N__23856),
            .I(N__23845));
    Span12Mux_h I__2852 (
            .O(N__23853),
            .I(N__23840));
    Sp12to4 I__2851 (
            .O(N__23848),
            .I(N__23840));
    Span12Mux_h I__2850 (
            .O(N__23845),
            .I(N__23837));
    Span12Mux_v I__2849 (
            .O(N__23840),
            .I(N__23834));
    Span12Mux_v I__2848 (
            .O(N__23837),
            .I(N__23829));
    Span12Mux_h I__2847 (
            .O(N__23834),
            .I(N__23829));
    Odrv12 I__2846 (
            .O(N__23829),
            .I(trig_ft_c));
    CascadeMux I__2845 (
            .O(N__23826),
            .I(un8_trig_prev_0_c5_a0_0_0_cascade_));
    CascadeMux I__2844 (
            .O(N__23823),
            .I(un8_trig_prev_0_c4_a0_1_cascade_));
    InMux I__2843 (
            .O(N__23820),
            .I(N__23811));
    InMux I__2842 (
            .O(N__23819),
            .I(N__23811));
    InMux I__2841 (
            .O(N__23818),
            .I(N__23811));
    LocalMux I__2840 (
            .O(N__23811),
            .I(sEETrigCounterZ0Z_5));
    InMux I__2839 (
            .O(N__23808),
            .I(N__23802));
    InMux I__2838 (
            .O(N__23807),
            .I(N__23802));
    LocalMux I__2837 (
            .O(N__23802),
            .I(sEETrigCounterZ0Z_6));
    InMux I__2836 (
            .O(N__23799),
            .I(N__23796));
    LocalMux I__2835 (
            .O(N__23796),
            .I(sEETrigCounterZ0Z_7));
    CascadeMux I__2834 (
            .O(N__23793),
            .I(un8_trig_prev_0_c7_a0_1_cascade_));
    InMux I__2833 (
            .O(N__23790),
            .I(N__23784));
    InMux I__2832 (
            .O(N__23789),
            .I(N__23784));
    LocalMux I__2831 (
            .O(N__23784),
            .I(un8_trig_prev_0_c4_a0_1));
    InMux I__2830 (
            .O(N__23781),
            .I(N__23778));
    LocalMux I__2829 (
            .O(N__23778),
            .I(N__23775));
    Odrv4 I__2828 (
            .O(N__23775),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15 ));
    InMux I__2827 (
            .O(N__23772),
            .I(N__23769));
    LocalMux I__2826 (
            .O(N__23769),
            .I(N__23766));
    Odrv4 I__2825 (
            .O(N__23766),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11 ));
    InMux I__2824 (
            .O(N__23763),
            .I(N__23760));
    LocalMux I__2823 (
            .O(N__23760),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10 ));
    InMux I__2822 (
            .O(N__23757),
            .I(N__23751));
    InMux I__2821 (
            .O(N__23756),
            .I(N__23751));
    LocalMux I__2820 (
            .O(N__23751),
            .I(N__23747));
    InMux I__2819 (
            .O(N__23750),
            .I(N__23744));
    Odrv12 I__2818 (
            .O(N__23747),
            .I(\spi_master_inst.sclk_gen_u0.N_158_7 ));
    LocalMux I__2817 (
            .O(N__23744),
            .I(\spi_master_inst.sclk_gen_u0.N_158_7 ));
    CascadeMux I__2816 (
            .O(N__23739),
            .I(N__23736));
    InMux I__2815 (
            .O(N__23736),
            .I(N__23732));
    InMux I__2814 (
            .O(N__23735),
            .I(N__23729));
    LocalMux I__2813 (
            .O(N__23732),
            .I(N__23721));
    LocalMux I__2812 (
            .O(N__23729),
            .I(N__23721));
    CascadeMux I__2811 (
            .O(N__23728),
            .I(N__23718));
    InMux I__2810 (
            .O(N__23727),
            .I(N__23712));
    InMux I__2809 (
            .O(N__23726),
            .I(N__23712));
    Span4Mux_h I__2808 (
            .O(N__23721),
            .I(N__23709));
    InMux I__2807 (
            .O(N__23718),
            .I(N__23704));
    InMux I__2806 (
            .O(N__23717),
            .I(N__23704));
    LocalMux I__2805 (
            .O(N__23712),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ));
    Odrv4 I__2804 (
            .O(N__23709),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ));
    LocalMux I__2803 (
            .O(N__23704),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ));
    CascadeMux I__2802 (
            .O(N__23697),
            .I(\spi_master_inst.sclk_gen_u0.N_158_7_cascade_ ));
    InMux I__2801 (
            .O(N__23694),
            .I(N__23689));
    InMux I__2800 (
            .O(N__23693),
            .I(N__23683));
    InMux I__2799 (
            .O(N__23692),
            .I(N__23683));
    LocalMux I__2798 (
            .O(N__23689),
            .I(N__23679));
    InMux I__2797 (
            .O(N__23688),
            .I(N__23675));
    LocalMux I__2796 (
            .O(N__23683),
            .I(N__23672));
    InMux I__2795 (
            .O(N__23682),
            .I(N__23669));
    Span12Mux_s11_h I__2794 (
            .O(N__23679),
            .I(N__23666));
    InMux I__2793 (
            .O(N__23678),
            .I(N__23663));
    LocalMux I__2792 (
            .O(N__23675),
            .I(N__23660));
    Odrv4 I__2791 (
            .O(N__23672),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ));
    LocalMux I__2790 (
            .O(N__23669),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ));
    Odrv12 I__2789 (
            .O(N__23666),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ));
    LocalMux I__2788 (
            .O(N__23663),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ));
    Odrv12 I__2787 (
            .O(N__23660),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ));
    InMux I__2786 (
            .O(N__23649),
            .I(N__23646));
    LocalMux I__2785 (
            .O(N__23646),
            .I(\spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0 ));
    InMux I__2784 (
            .O(N__23643),
            .I(N__23636));
    InMux I__2783 (
            .O(N__23642),
            .I(N__23636));
    InMux I__2782 (
            .O(N__23641),
            .I(N__23633));
    LocalMux I__2781 (
            .O(N__23636),
            .I(\spi_master_inst.sclk_gen_u0.falling_count_start_iZ0 ));
    LocalMux I__2780 (
            .O(N__23633),
            .I(\spi_master_inst.sclk_gen_u0.falling_count_start_iZ0 ));
    CascadeMux I__2779 (
            .O(N__23628),
            .I(N__23625));
    InMux I__2778 (
            .O(N__23625),
            .I(N__23622));
    LocalMux I__2777 (
            .O(N__23622),
            .I(N__23619));
    Odrv4 I__2776 (
            .O(N__23619),
            .I(un3_trig_0_0));
    CascadeMux I__2775 (
            .O(N__23616),
            .I(un3_trig_0_0_cascade_));
    InMux I__2774 (
            .O(N__23613),
            .I(N__23610));
    LocalMux I__2773 (
            .O(N__23610),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2 ));
    InMux I__2772 (
            .O(N__23607),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4 ));
    InMux I__2771 (
            .O(N__23604),
            .I(N__23601));
    LocalMux I__2770 (
            .O(N__23601),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO ));
    InMux I__2769 (
            .O(N__23598),
            .I(N__23595));
    LocalMux I__2768 (
            .O(N__23595),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO ));
    InMux I__2767 (
            .O(N__23592),
            .I(N__23589));
    LocalMux I__2766 (
            .O(N__23589),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12 ));
    InMux I__2765 (
            .O(N__23586),
            .I(N__23583));
    LocalMux I__2764 (
            .O(N__23583),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2 ));
    InMux I__2763 (
            .O(N__23580),
            .I(N__23577));
    LocalMux I__2762 (
            .O(N__23577),
            .I(N__23574));
    Odrv12 I__2761 (
            .O(N__23574),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3 ));
    InMux I__2760 (
            .O(N__23571),
            .I(N__23568));
    LocalMux I__2759 (
            .O(N__23568),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4 ));
    InMux I__2758 (
            .O(N__23565),
            .I(N__23562));
    LocalMux I__2757 (
            .O(N__23562),
            .I(N__23559));
    Span4Mux_h I__2756 (
            .O(N__23559),
            .I(N__23556));
    Odrv4 I__2755 (
            .O(N__23556),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5 ));
    InMux I__2754 (
            .O(N__23553),
            .I(un1_button_debounce_counter_cry_21));
    InMux I__2753 (
            .O(N__23550),
            .I(bfn_8_20_0_));
    CascadeMux I__2752 (
            .O(N__23547),
            .I(N__23544));
    InMux I__2751 (
            .O(N__23544),
            .I(N__23540));
    InMux I__2750 (
            .O(N__23543),
            .I(N__23537));
    LocalMux I__2749 (
            .O(N__23540),
            .I(N__23534));
    LocalMux I__2748 (
            .O(N__23537),
            .I(button_debounce_counterZ0Z_23));
    Odrv4 I__2747 (
            .O(N__23534),
            .I(button_debounce_counterZ0Z_23));
    InMux I__2746 (
            .O(N__23529),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0 ));
    InMux I__2745 (
            .O(N__23526),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1 ));
    InMux I__2744 (
            .O(N__23523),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2 ));
    InMux I__2743 (
            .O(N__23520),
            .I(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3 ));
    CascadeMux I__2742 (
            .O(N__23517),
            .I(N__23513));
    InMux I__2741 (
            .O(N__23516),
            .I(N__23510));
    InMux I__2740 (
            .O(N__23513),
            .I(N__23507));
    LocalMux I__2739 (
            .O(N__23510),
            .I(button_debounce_counterZ0Z_13));
    LocalMux I__2738 (
            .O(N__23507),
            .I(button_debounce_counterZ0Z_13));
    InMux I__2737 (
            .O(N__23502),
            .I(un1_button_debounce_counter_cry_12));
    InMux I__2736 (
            .O(N__23499),
            .I(N__23495));
    InMux I__2735 (
            .O(N__23498),
            .I(N__23492));
    LocalMux I__2734 (
            .O(N__23495),
            .I(button_debounce_counterZ0Z_14));
    LocalMux I__2733 (
            .O(N__23492),
            .I(button_debounce_counterZ0Z_14));
    InMux I__2732 (
            .O(N__23487),
            .I(un1_button_debounce_counter_cry_13));
    InMux I__2731 (
            .O(N__23484),
            .I(N__23480));
    InMux I__2730 (
            .O(N__23483),
            .I(N__23477));
    LocalMux I__2729 (
            .O(N__23480),
            .I(button_debounce_counterZ0Z_15));
    LocalMux I__2728 (
            .O(N__23477),
            .I(button_debounce_counterZ0Z_15));
    InMux I__2727 (
            .O(N__23472),
            .I(un1_button_debounce_counter_cry_14));
    InMux I__2726 (
            .O(N__23469),
            .I(N__23465));
    InMux I__2725 (
            .O(N__23468),
            .I(N__23462));
    LocalMux I__2724 (
            .O(N__23465),
            .I(button_debounce_counterZ0Z_16));
    LocalMux I__2723 (
            .O(N__23462),
            .I(button_debounce_counterZ0Z_16));
    InMux I__2722 (
            .O(N__23457),
            .I(un1_button_debounce_counter_cry_15));
    InMux I__2721 (
            .O(N__23454),
            .I(N__23451));
    LocalMux I__2720 (
            .O(N__23451),
            .I(N__23447));
    InMux I__2719 (
            .O(N__23450),
            .I(N__23444));
    Odrv12 I__2718 (
            .O(N__23447),
            .I(button_debounce_counterZ0Z_17));
    LocalMux I__2717 (
            .O(N__23444),
            .I(button_debounce_counterZ0Z_17));
    InMux I__2716 (
            .O(N__23439),
            .I(bfn_8_19_0_));
    InMux I__2715 (
            .O(N__23436),
            .I(N__23433));
    LocalMux I__2714 (
            .O(N__23433),
            .I(N__23430));
    Span4Mux_v I__2713 (
            .O(N__23430),
            .I(N__23426));
    InMux I__2712 (
            .O(N__23429),
            .I(N__23423));
    Odrv4 I__2711 (
            .O(N__23426),
            .I(button_debounce_counterZ0Z_18));
    LocalMux I__2710 (
            .O(N__23423),
            .I(button_debounce_counterZ0Z_18));
    InMux I__2709 (
            .O(N__23418),
            .I(un1_button_debounce_counter_cry_17));
    InMux I__2708 (
            .O(N__23415),
            .I(N__23412));
    LocalMux I__2707 (
            .O(N__23412),
            .I(N__23408));
    InMux I__2706 (
            .O(N__23411),
            .I(N__23405));
    Odrv12 I__2705 (
            .O(N__23408),
            .I(button_debounce_counterZ0Z_19));
    LocalMux I__2704 (
            .O(N__23405),
            .I(button_debounce_counterZ0Z_19));
    InMux I__2703 (
            .O(N__23400),
            .I(un1_button_debounce_counter_cry_18));
    CascadeMux I__2702 (
            .O(N__23397),
            .I(N__23394));
    InMux I__2701 (
            .O(N__23394),
            .I(N__23391));
    LocalMux I__2700 (
            .O(N__23391),
            .I(N__23388));
    Span4Mux_v I__2699 (
            .O(N__23388),
            .I(N__23384));
    InMux I__2698 (
            .O(N__23387),
            .I(N__23381));
    Odrv4 I__2697 (
            .O(N__23384),
            .I(button_debounce_counterZ0Z_20));
    LocalMux I__2696 (
            .O(N__23381),
            .I(button_debounce_counterZ0Z_20));
    InMux I__2695 (
            .O(N__23376),
            .I(un1_button_debounce_counter_cry_19));
    InMux I__2694 (
            .O(N__23373),
            .I(un1_button_debounce_counter_cry_20));
    InMux I__2693 (
            .O(N__23370),
            .I(un1_button_debounce_counter_cry_4));
    InMux I__2692 (
            .O(N__23367),
            .I(N__23363));
    InMux I__2691 (
            .O(N__23366),
            .I(N__23360));
    LocalMux I__2690 (
            .O(N__23363),
            .I(button_debounce_counterZ0Z_6));
    LocalMux I__2689 (
            .O(N__23360),
            .I(button_debounce_counterZ0Z_6));
    InMux I__2688 (
            .O(N__23355),
            .I(un1_button_debounce_counter_cry_5));
    InMux I__2687 (
            .O(N__23352),
            .I(N__23348));
    InMux I__2686 (
            .O(N__23351),
            .I(N__23345));
    LocalMux I__2685 (
            .O(N__23348),
            .I(button_debounce_counterZ0Z_7));
    LocalMux I__2684 (
            .O(N__23345),
            .I(button_debounce_counterZ0Z_7));
    InMux I__2683 (
            .O(N__23340),
            .I(un1_button_debounce_counter_cry_6));
    InMux I__2682 (
            .O(N__23337),
            .I(N__23333));
    InMux I__2681 (
            .O(N__23336),
            .I(N__23330));
    LocalMux I__2680 (
            .O(N__23333),
            .I(button_debounce_counterZ0Z_8));
    LocalMux I__2679 (
            .O(N__23330),
            .I(button_debounce_counterZ0Z_8));
    InMux I__2678 (
            .O(N__23325),
            .I(un1_button_debounce_counter_cry_7));
    CascadeMux I__2677 (
            .O(N__23322),
            .I(N__23318));
    InMux I__2676 (
            .O(N__23321),
            .I(N__23315));
    InMux I__2675 (
            .O(N__23318),
            .I(N__23312));
    LocalMux I__2674 (
            .O(N__23315),
            .I(button_debounce_counterZ0Z_9));
    LocalMux I__2673 (
            .O(N__23312),
            .I(button_debounce_counterZ0Z_9));
    InMux I__2672 (
            .O(N__23307),
            .I(bfn_8_18_0_));
    InMux I__2671 (
            .O(N__23304),
            .I(N__23300));
    InMux I__2670 (
            .O(N__23303),
            .I(N__23297));
    LocalMux I__2669 (
            .O(N__23300),
            .I(button_debounce_counterZ0Z_10));
    LocalMux I__2668 (
            .O(N__23297),
            .I(button_debounce_counterZ0Z_10));
    InMux I__2667 (
            .O(N__23292),
            .I(un1_button_debounce_counter_cry_9));
    InMux I__2666 (
            .O(N__23289),
            .I(N__23285));
    InMux I__2665 (
            .O(N__23288),
            .I(N__23282));
    LocalMux I__2664 (
            .O(N__23285),
            .I(button_debounce_counterZ0Z_11));
    LocalMux I__2663 (
            .O(N__23282),
            .I(button_debounce_counterZ0Z_11));
    InMux I__2662 (
            .O(N__23277),
            .I(un1_button_debounce_counter_cry_10));
    InMux I__2661 (
            .O(N__23274),
            .I(N__23270));
    InMux I__2660 (
            .O(N__23273),
            .I(N__23267));
    LocalMux I__2659 (
            .O(N__23270),
            .I(button_debounce_counterZ0Z_12));
    LocalMux I__2658 (
            .O(N__23267),
            .I(button_debounce_counterZ0Z_12));
    InMux I__2657 (
            .O(N__23262),
            .I(un1_button_debounce_counter_cry_11));
    InMux I__2656 (
            .O(N__23259),
            .I(sCounter_cry_18));
    InMux I__2655 (
            .O(N__23256),
            .I(sCounter_cry_19));
    InMux I__2654 (
            .O(N__23253),
            .I(sCounter_cry_20));
    InMux I__2653 (
            .O(N__23250),
            .I(sCounter_cry_21));
    InMux I__2652 (
            .O(N__23247),
            .I(N__23231));
    InMux I__2651 (
            .O(N__23246),
            .I(N__23231));
    InMux I__2650 (
            .O(N__23245),
            .I(N__23231));
    InMux I__2649 (
            .O(N__23244),
            .I(N__23231));
    InMux I__2648 (
            .O(N__23243),
            .I(N__23206));
    InMux I__2647 (
            .O(N__23242),
            .I(N__23206));
    InMux I__2646 (
            .O(N__23241),
            .I(N__23206));
    InMux I__2645 (
            .O(N__23240),
            .I(N__23206));
    LocalMux I__2644 (
            .O(N__23231),
            .I(N__23203));
    InMux I__2643 (
            .O(N__23230),
            .I(N__23194));
    InMux I__2642 (
            .O(N__23229),
            .I(N__23194));
    InMux I__2641 (
            .O(N__23228),
            .I(N__23194));
    InMux I__2640 (
            .O(N__23227),
            .I(N__23194));
    InMux I__2639 (
            .O(N__23226),
            .I(N__23185));
    InMux I__2638 (
            .O(N__23225),
            .I(N__23185));
    InMux I__2637 (
            .O(N__23224),
            .I(N__23185));
    InMux I__2636 (
            .O(N__23223),
            .I(N__23185));
    InMux I__2635 (
            .O(N__23222),
            .I(N__23176));
    InMux I__2634 (
            .O(N__23221),
            .I(N__23176));
    InMux I__2633 (
            .O(N__23220),
            .I(N__23176));
    InMux I__2632 (
            .O(N__23219),
            .I(N__23176));
    InMux I__2631 (
            .O(N__23218),
            .I(N__23167));
    InMux I__2630 (
            .O(N__23217),
            .I(N__23167));
    InMux I__2629 (
            .O(N__23216),
            .I(N__23167));
    InMux I__2628 (
            .O(N__23215),
            .I(N__23167));
    LocalMux I__2627 (
            .O(N__23206),
            .I(LED_ACQ_c_i));
    Odrv4 I__2626 (
            .O(N__23203),
            .I(LED_ACQ_c_i));
    LocalMux I__2625 (
            .O(N__23194),
            .I(LED_ACQ_c_i));
    LocalMux I__2624 (
            .O(N__23185),
            .I(LED_ACQ_c_i));
    LocalMux I__2623 (
            .O(N__23176),
            .I(LED_ACQ_c_i));
    LocalMux I__2622 (
            .O(N__23167),
            .I(LED_ACQ_c_i));
    InMux I__2621 (
            .O(N__23154),
            .I(sCounter_cry_22));
    InMux I__2620 (
            .O(N__23151),
            .I(un1_button_debounce_counter_cry_1));
    InMux I__2619 (
            .O(N__23148),
            .I(un1_button_debounce_counter_cry_2));
    InMux I__2618 (
            .O(N__23145),
            .I(un1_button_debounce_counter_cry_3));
    InMux I__2617 (
            .O(N__23142),
            .I(sCounter_cry_9));
    InMux I__2616 (
            .O(N__23139),
            .I(sCounter_cry_10));
    InMux I__2615 (
            .O(N__23136),
            .I(sCounter_cry_11));
    InMux I__2614 (
            .O(N__23133),
            .I(sCounter_cry_12));
    InMux I__2613 (
            .O(N__23130),
            .I(sCounter_cry_13));
    InMux I__2612 (
            .O(N__23127),
            .I(sCounter_cry_14));
    InMux I__2611 (
            .O(N__23124),
            .I(bfn_8_16_0_));
    InMux I__2610 (
            .O(N__23121),
            .I(sCounter_cry_16));
    InMux I__2609 (
            .O(N__23118),
            .I(sCounter_cry_17));
    InMux I__2608 (
            .O(N__23115),
            .I(sCounter_cry_0));
    InMux I__2607 (
            .O(N__23112),
            .I(sCounter_cry_1));
    InMux I__2606 (
            .O(N__23109),
            .I(sCounter_cry_2));
    InMux I__2605 (
            .O(N__23106),
            .I(sCounter_cry_3));
    InMux I__2604 (
            .O(N__23103),
            .I(sCounter_cry_4));
    InMux I__2603 (
            .O(N__23100),
            .I(sCounter_cry_5));
    InMux I__2602 (
            .O(N__23097),
            .I(sCounter_cry_6));
    InMux I__2601 (
            .O(N__23094),
            .I(bfn_8_15_0_));
    InMux I__2600 (
            .O(N__23091),
            .I(sCounter_cry_8));
    InMux I__2599 (
            .O(N__23088),
            .I(N__23085));
    LocalMux I__2598 (
            .O(N__23085),
            .I(sEEPeriodZ0Z_20));
    CascadeMux I__2597 (
            .O(N__23082),
            .I(N__23079));
    InMux I__2596 (
            .O(N__23079),
            .I(N__23076));
    LocalMux I__2595 (
            .O(N__23076),
            .I(sEEPeriod_i_20));
    InMux I__2594 (
            .O(N__23073),
            .I(N__23070));
    LocalMux I__2593 (
            .O(N__23070),
            .I(sEEPeriodZ0Z_21));
    InMux I__2592 (
            .O(N__23067),
            .I(N__23064));
    LocalMux I__2591 (
            .O(N__23064),
            .I(sEEPeriod_i_21));
    InMux I__2590 (
            .O(N__23061),
            .I(N__23058));
    LocalMux I__2589 (
            .O(N__23058),
            .I(sEEPeriodZ0Z_22));
    InMux I__2588 (
            .O(N__23055),
            .I(N__23052));
    LocalMux I__2587 (
            .O(N__23052),
            .I(sEEPeriod_i_22));
    InMux I__2586 (
            .O(N__23049),
            .I(N__23046));
    LocalMux I__2585 (
            .O(N__23046),
            .I(sEEPeriodZ0Z_23));
    CascadeMux I__2584 (
            .O(N__23043),
            .I(N__23040));
    InMux I__2583 (
            .O(N__23040),
            .I(N__23037));
    LocalMux I__2582 (
            .O(N__23037),
            .I(sEEPeriod_i_23));
    InMux I__2581 (
            .O(N__23034),
            .I(bfn_8_13_0_));
    CascadeMux I__2580 (
            .O(N__23031),
            .I(N__23028));
    InMux I__2579 (
            .O(N__23028),
            .I(N__23025));
    LocalMux I__2578 (
            .O(N__23025),
            .I(un1_reset_rpi_inv_2_i_o3_15));
    CascadeMux I__2577 (
            .O(N__23022),
            .I(N__23019));
    InMux I__2576 (
            .O(N__23019),
            .I(N__23016));
    LocalMux I__2575 (
            .O(N__23016),
            .I(un1_reset_rpi_inv_2_i_o3_11));
    InMux I__2574 (
            .O(N__23013),
            .I(N__23010));
    LocalMux I__2573 (
            .O(N__23010),
            .I(sbuttonModeStatus_0_sqmuxa_17));
    InMux I__2572 (
            .O(N__23007),
            .I(bfn_8_14_0_));
    CascadeMux I__2571 (
            .O(N__23004),
            .I(N__23001));
    InMux I__2570 (
            .O(N__23001),
            .I(N__22998));
    LocalMux I__2569 (
            .O(N__22998),
            .I(sEEPeriod_i_12));
    CascadeMux I__2568 (
            .O(N__22995),
            .I(N__22992));
    InMux I__2567 (
            .O(N__22992),
            .I(N__22989));
    LocalMux I__2566 (
            .O(N__22989),
            .I(sEEPeriod_i_13));
    CascadeMux I__2565 (
            .O(N__22986),
            .I(N__22983));
    InMux I__2564 (
            .O(N__22983),
            .I(N__22980));
    LocalMux I__2563 (
            .O(N__22980),
            .I(sEEPeriod_i_14));
    CascadeMux I__2562 (
            .O(N__22977),
            .I(N__22974));
    InMux I__2561 (
            .O(N__22974),
            .I(N__22971));
    LocalMux I__2560 (
            .O(N__22971),
            .I(sEEPeriod_i_15));
    InMux I__2559 (
            .O(N__22968),
            .I(N__22965));
    LocalMux I__2558 (
            .O(N__22965),
            .I(sEEPeriodZ0Z_16));
    CascadeMux I__2557 (
            .O(N__22962),
            .I(N__22959));
    InMux I__2556 (
            .O(N__22959),
            .I(N__22956));
    LocalMux I__2555 (
            .O(N__22956),
            .I(sEEPeriod_i_16));
    InMux I__2554 (
            .O(N__22953),
            .I(N__22950));
    LocalMux I__2553 (
            .O(N__22950),
            .I(sEEPeriodZ0Z_17));
    CascadeMux I__2552 (
            .O(N__22947),
            .I(N__22944));
    InMux I__2551 (
            .O(N__22944),
            .I(N__22941));
    LocalMux I__2550 (
            .O(N__22941),
            .I(sEEPeriod_i_17));
    InMux I__2549 (
            .O(N__22938),
            .I(N__22935));
    LocalMux I__2548 (
            .O(N__22935),
            .I(sEEPeriodZ0Z_18));
    CascadeMux I__2547 (
            .O(N__22932),
            .I(N__22929));
    InMux I__2546 (
            .O(N__22929),
            .I(N__22926));
    LocalMux I__2545 (
            .O(N__22926),
            .I(sEEPeriod_i_18));
    InMux I__2544 (
            .O(N__22923),
            .I(N__22920));
    LocalMux I__2543 (
            .O(N__22920),
            .I(sEEPeriodZ0Z_19));
    CascadeMux I__2542 (
            .O(N__22917),
            .I(N__22914));
    InMux I__2541 (
            .O(N__22914),
            .I(N__22911));
    LocalMux I__2540 (
            .O(N__22911),
            .I(sEEPeriod_i_19));
    InMux I__2539 (
            .O(N__22908),
            .I(N__22905));
    LocalMux I__2538 (
            .O(N__22905),
            .I(sEEPeriodZ0Z_4));
    CascadeMux I__2537 (
            .O(N__22902),
            .I(N__22899));
    InMux I__2536 (
            .O(N__22899),
            .I(N__22896));
    LocalMux I__2535 (
            .O(N__22896),
            .I(sEEPeriod_i_4));
    InMux I__2534 (
            .O(N__22893),
            .I(N__22890));
    LocalMux I__2533 (
            .O(N__22890),
            .I(sEEPeriodZ0Z_5));
    CascadeMux I__2532 (
            .O(N__22887),
            .I(N__22884));
    InMux I__2531 (
            .O(N__22884),
            .I(N__22881));
    LocalMux I__2530 (
            .O(N__22881),
            .I(sEEPeriod_i_5));
    InMux I__2529 (
            .O(N__22878),
            .I(N__22875));
    LocalMux I__2528 (
            .O(N__22875),
            .I(sEEPeriodZ0Z_6));
    CascadeMux I__2527 (
            .O(N__22872),
            .I(N__22869));
    InMux I__2526 (
            .O(N__22869),
            .I(N__22866));
    LocalMux I__2525 (
            .O(N__22866),
            .I(sEEPeriod_i_6));
    InMux I__2524 (
            .O(N__22863),
            .I(N__22860));
    LocalMux I__2523 (
            .O(N__22860),
            .I(sEEPeriodZ0Z_7));
    CascadeMux I__2522 (
            .O(N__22857),
            .I(N__22854));
    InMux I__2521 (
            .O(N__22854),
            .I(N__22851));
    LocalMux I__2520 (
            .O(N__22851),
            .I(sEEPeriod_i_7));
    CascadeMux I__2519 (
            .O(N__22848),
            .I(N__22845));
    InMux I__2518 (
            .O(N__22845),
            .I(N__22842));
    LocalMux I__2517 (
            .O(N__22842),
            .I(sEEPeriod_i_8));
    CascadeMux I__2516 (
            .O(N__22839),
            .I(N__22836));
    InMux I__2515 (
            .O(N__22836),
            .I(N__22833));
    LocalMux I__2514 (
            .O(N__22833),
            .I(sEEPeriod_i_9));
    CascadeMux I__2513 (
            .O(N__22830),
            .I(N__22827));
    InMux I__2512 (
            .O(N__22827),
            .I(N__22824));
    LocalMux I__2511 (
            .O(N__22824),
            .I(sEEPeriod_i_10));
    CascadeMux I__2510 (
            .O(N__22821),
            .I(N__22818));
    InMux I__2509 (
            .O(N__22818),
            .I(N__22815));
    LocalMux I__2508 (
            .O(N__22815),
            .I(sEEPeriod_i_11));
    CascadeMux I__2507 (
            .O(N__22812),
            .I(g2_0_0_cascade_));
    InMux I__2506 (
            .O(N__22809),
            .I(N__22806));
    LocalMux I__2505 (
            .O(N__22806),
            .I(N__22803));
    Odrv4 I__2504 (
            .O(N__22803),
            .I(g1_0_0_0));
    InMux I__2503 (
            .O(N__22800),
            .I(N__22797));
    LocalMux I__2502 (
            .O(N__22797),
            .I(g1_0_1));
    InMux I__2501 (
            .O(N__22794),
            .I(N__22791));
    LocalMux I__2500 (
            .O(N__22791),
            .I(N__22788));
    Span4Mux_v I__2499 (
            .O(N__22788),
            .I(N__22785));
    Odrv4 I__2498 (
            .O(N__22785),
            .I(g0_2_0));
    InMux I__2497 (
            .O(N__22782),
            .I(N__22779));
    LocalMux I__2496 (
            .O(N__22779),
            .I(g1_4));
    CascadeMux I__2495 (
            .O(N__22776),
            .I(g2_0_cascade_));
    InMux I__2494 (
            .O(N__22773),
            .I(N__22770));
    LocalMux I__2493 (
            .O(N__22770),
            .I(sEEPeriodZ0Z_0));
    CascadeMux I__2492 (
            .O(N__22767),
            .I(N__22764));
    InMux I__2491 (
            .O(N__22764),
            .I(N__22761));
    LocalMux I__2490 (
            .O(N__22761),
            .I(sEEPeriod_i_0));
    InMux I__2489 (
            .O(N__22758),
            .I(N__22755));
    LocalMux I__2488 (
            .O(N__22755),
            .I(sEEPeriodZ0Z_1));
    CascadeMux I__2487 (
            .O(N__22752),
            .I(N__22749));
    InMux I__2486 (
            .O(N__22749),
            .I(N__22746));
    LocalMux I__2485 (
            .O(N__22746),
            .I(sEEPeriod_i_1));
    InMux I__2484 (
            .O(N__22743),
            .I(N__22740));
    LocalMux I__2483 (
            .O(N__22740),
            .I(sEEPeriodZ0Z_2));
    CascadeMux I__2482 (
            .O(N__22737),
            .I(N__22734));
    InMux I__2481 (
            .O(N__22734),
            .I(N__22731));
    LocalMux I__2480 (
            .O(N__22731),
            .I(sEEPeriod_i_2));
    InMux I__2479 (
            .O(N__22728),
            .I(N__22725));
    LocalMux I__2478 (
            .O(N__22725),
            .I(sEEPeriodZ0Z_3));
    CascadeMux I__2477 (
            .O(N__22722),
            .I(N__22719));
    InMux I__2476 (
            .O(N__22719),
            .I(N__22716));
    LocalMux I__2475 (
            .O(N__22716),
            .I(sEEPeriod_i_3));
    CascadeMux I__2474 (
            .O(N__22713),
            .I(N__22710));
    InMux I__2473 (
            .O(N__22710),
            .I(N__22707));
    LocalMux I__2472 (
            .O(N__22707),
            .I(g0_2_0_2));
    InMux I__2471 (
            .O(N__22704),
            .I(N__22701));
    LocalMux I__2470 (
            .O(N__22701),
            .I(N__22698));
    Span4Mux_v I__2469 (
            .O(N__22698),
            .I(N__22695));
    Odrv4 I__2468 (
            .O(N__22695),
            .I(g1_1));
    CascadeMux I__2467 (
            .O(N__22692),
            .I(g2_0_2_cascade_));
    InMux I__2466 (
            .O(N__22689),
            .I(N__22686));
    LocalMux I__2465 (
            .O(N__22686),
            .I(g1_0_3));
    InMux I__2464 (
            .O(N__22683),
            .I(N__22680));
    LocalMux I__2463 (
            .O(N__22680),
            .I(g0_2_0_1));
    CascadeMux I__2462 (
            .O(N__22677),
            .I(g2_0_1_cascade_));
    InMux I__2461 (
            .O(N__22674),
            .I(N__22671));
    LocalMux I__2460 (
            .O(N__22671),
            .I(N__22668));
    Odrv4 I__2459 (
            .O(N__22668),
            .I(g1_2));
    InMux I__2458 (
            .O(N__22665),
            .I(N__22662));
    LocalMux I__2457 (
            .O(N__22662),
            .I(g1_0_0_1));
    InMux I__2456 (
            .O(N__22659),
            .I(N__22656));
    LocalMux I__2455 (
            .O(N__22656),
            .I(g1_0_2));
    CascadeMux I__2454 (
            .O(N__22653),
            .I(N__22650));
    InMux I__2453 (
            .O(N__22650),
            .I(N__22647));
    LocalMux I__2452 (
            .O(N__22647),
            .I(N__22644));
    Odrv4 I__2451 (
            .O(N__22644),
            .I(g0_2_0_0));
    InMux I__2450 (
            .O(N__22641),
            .I(N__22631));
    InMux I__2449 (
            .O(N__22640),
            .I(N__22631));
    InMux I__2448 (
            .O(N__22639),
            .I(N__22624));
    InMux I__2447 (
            .O(N__22638),
            .I(N__22619));
    InMux I__2446 (
            .O(N__22637),
            .I(N__22619));
    CascadeMux I__2445 (
            .O(N__22636),
            .I(N__22614));
    LocalMux I__2444 (
            .O(N__22631),
            .I(N__22611));
    InMux I__2443 (
            .O(N__22630),
            .I(N__22606));
    InMux I__2442 (
            .O(N__22629),
            .I(N__22606));
    InMux I__2441 (
            .O(N__22628),
            .I(N__22601));
    InMux I__2440 (
            .O(N__22627),
            .I(N__22601));
    LocalMux I__2439 (
            .O(N__22624),
            .I(N__22598));
    LocalMux I__2438 (
            .O(N__22619),
            .I(N__22595));
    InMux I__2437 (
            .O(N__22618),
            .I(N__22590));
    InMux I__2436 (
            .O(N__22617),
            .I(N__22590));
    InMux I__2435 (
            .O(N__22614),
            .I(N__22587));
    Span4Mux_v I__2434 (
            .O(N__22611),
            .I(N__22576));
    LocalMux I__2433 (
            .O(N__22606),
            .I(N__22576));
    LocalMux I__2432 (
            .O(N__22601),
            .I(N__22576));
    Span4Mux_h I__2431 (
            .O(N__22598),
            .I(N__22576));
    Span4Mux_h I__2430 (
            .O(N__22595),
            .I(N__22576));
    LocalMux I__2429 (
            .O(N__22590),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ));
    LocalMux I__2428 (
            .O(N__22587),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ));
    Odrv4 I__2427 (
            .O(N__22576),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ));
    InMux I__2426 (
            .O(N__22569),
            .I(N__22566));
    LocalMux I__2425 (
            .O(N__22566),
            .I(N__22563));
    Span4Mux_v I__2424 (
            .O(N__22563),
            .I(N__22560));
    Odrv4 I__2423 (
            .O(N__22560),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12 ));
    InMux I__2422 (
            .O(N__22557),
            .I(N__22548));
    InMux I__2421 (
            .O(N__22556),
            .I(N__22548));
    InMux I__2420 (
            .O(N__22555),
            .I(N__22548));
    LocalMux I__2419 (
            .O(N__22548),
            .I(\spi_master_inst.sclk_gen_u0.N_150_0 ));
    InMux I__2418 (
            .O(N__22545),
            .I(N__22542));
    LocalMux I__2417 (
            .O(N__22542),
            .I(N__22539));
    Odrv4 I__2416 (
            .O(N__22539),
            .I(\spi_master_inst.sclk_gen_u0.N_36 ));
    CascadeMux I__2415 (
            .O(N__22536),
            .I(N__22533));
    InMux I__2414 (
            .O(N__22533),
            .I(N__22526));
    InMux I__2413 (
            .O(N__22532),
            .I(N__22526));
    InMux I__2412 (
            .O(N__22531),
            .I(N__22523));
    LocalMux I__2411 (
            .O(N__22526),
            .I(N__22520));
    LocalMux I__2410 (
            .O(N__22523),
            .I(N__22517));
    Span4Mux_v I__2409 (
            .O(N__22520),
            .I(N__22514));
    Span4Mux_h I__2408 (
            .O(N__22517),
            .I(N__22510));
    Span4Mux_h I__2407 (
            .O(N__22514),
            .I(N__22507));
    InMux I__2406 (
            .O(N__22513),
            .I(N__22504));
    Span4Mux_h I__2405 (
            .O(N__22510),
            .I(N__22501));
    Odrv4 I__2404 (
            .O(N__22507),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0 ));
    LocalMux I__2403 (
            .O(N__22504),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0 ));
    Odrv4 I__2402 (
            .O(N__22501),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0 ));
    InMux I__2401 (
            .O(N__22494),
            .I(N__22487));
    InMux I__2400 (
            .O(N__22493),
            .I(N__22487));
    InMux I__2399 (
            .O(N__22492),
            .I(N__22484));
    LocalMux I__2398 (
            .O(N__22487),
            .I(N__22480));
    LocalMux I__2397 (
            .O(N__22484),
            .I(N__22477));
    InMux I__2396 (
            .O(N__22483),
            .I(N__22474));
    Span4Mux_v I__2395 (
            .O(N__22480),
            .I(N__22469));
    Span4Mux_v I__2394 (
            .O(N__22477),
            .I(N__22469));
    LocalMux I__2393 (
            .O(N__22474),
            .I(\spi_master_inst.sclk_gen_u0.div_clk_iZ0 ));
    Odrv4 I__2392 (
            .O(N__22469),
            .I(\spi_master_inst.sclk_gen_u0.div_clk_iZ0 ));
    InMux I__2391 (
            .O(N__22464),
            .I(N__22461));
    LocalMux I__2390 (
            .O(N__22461),
            .I(\spi_master_inst.sclk_gen_u0.delay_clk_iZ0 ));
    InMux I__2389 (
            .O(N__22458),
            .I(N__22455));
    LocalMux I__2388 (
            .O(N__22455),
            .I(N__22452));
    Span4Mux_v I__2387 (
            .O(N__22452),
            .I(N__22449));
    Odrv4 I__2386 (
            .O(N__22449),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14 ));
    InMux I__2385 (
            .O(N__22446),
            .I(N__22443));
    LocalMux I__2384 (
            .O(N__22443),
            .I(N__22440));
    Odrv4 I__2383 (
            .O(N__22440),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0 ));
    InMux I__2382 (
            .O(N__22437),
            .I(N__22434));
    LocalMux I__2381 (
            .O(N__22434),
            .I(N__22431));
    Odrv4 I__2380 (
            .O(N__22431),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8 ));
    InMux I__2379 (
            .O(N__22428),
            .I(N__22425));
    LocalMux I__2378 (
            .O(N__22425),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9 ));
    InMux I__2377 (
            .O(N__22422),
            .I(N__22419));
    LocalMux I__2376 (
            .O(N__22419),
            .I(N__22416));
    Span4Mux_v I__2375 (
            .O(N__22416),
            .I(N__22413));
    Odrv4 I__2374 (
            .O(N__22413),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7 ));
    InMux I__2373 (
            .O(N__22410),
            .I(N__22407));
    LocalMux I__2372 (
            .O(N__22407),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1 ));
    InMux I__2371 (
            .O(N__22404),
            .I(N__22401));
    LocalMux I__2370 (
            .O(N__22401),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13 ));
    InMux I__2369 (
            .O(N__22398),
            .I(N__22395));
    LocalMux I__2368 (
            .O(N__22395),
            .I(N__22392));
    Span4Mux_h I__2367 (
            .O(N__22392),
            .I(N__22389));
    Odrv4 I__2366 (
            .O(N__22389),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10 ));
    InMux I__2365 (
            .O(N__22386),
            .I(sCounterRAM_cry_4));
    InMux I__2364 (
            .O(N__22383),
            .I(sCounterRAM_cry_5));
    InMux I__2363 (
            .O(N__22380),
            .I(N__22364));
    InMux I__2362 (
            .O(N__22379),
            .I(N__22364));
    InMux I__2361 (
            .O(N__22378),
            .I(N__22364));
    InMux I__2360 (
            .O(N__22377),
            .I(N__22364));
    InMux I__2359 (
            .O(N__22376),
            .I(N__22355));
    InMux I__2358 (
            .O(N__22375),
            .I(N__22355));
    InMux I__2357 (
            .O(N__22374),
            .I(N__22355));
    InMux I__2356 (
            .O(N__22373),
            .I(N__22355));
    LocalMux I__2355 (
            .O(N__22364),
            .I(un1_spi_data_miso_0_sqmuxa_1_i_0_N_3_0));
    LocalMux I__2354 (
            .O(N__22355),
            .I(un1_spi_data_miso_0_sqmuxa_1_i_0_N_3_0));
    InMux I__2353 (
            .O(N__22350),
            .I(sCounterRAM_cry_6));
    InMux I__2352 (
            .O(N__22347),
            .I(N__22344));
    LocalMux I__2351 (
            .O(N__22344),
            .I(sSPI_MSB0LSB1_RNIO3VPZ0Z1));
    CascadeMux I__2350 (
            .O(N__22341),
            .I(N__22338));
    InMux I__2349 (
            .O(N__22338),
            .I(N__22335));
    LocalMux I__2348 (
            .O(N__22335),
            .I(N__22332));
    Span4Mux_v I__2347 (
            .O(N__22332),
            .I(N__22329));
    Span4Mux_h I__2346 (
            .O(N__22329),
            .I(N__22326));
    Odrv4 I__2345 (
            .O(N__22326),
            .I(sbuttonModeStatus_0_sqmuxa_16));
    InMux I__2344 (
            .O(N__22323),
            .I(N__22320));
    LocalMux I__2343 (
            .O(N__22320),
            .I(N__22317));
    Span4Mux_v I__2342 (
            .O(N__22317),
            .I(N__22314));
    Odrv4 I__2341 (
            .O(N__22314),
            .I(sbuttonModeStatus_0_sqmuxa_14));
    InMux I__2340 (
            .O(N__22311),
            .I(N__22308));
    LocalMux I__2339 (
            .O(N__22308),
            .I(N__22305));
    Sp12to4 I__2338 (
            .O(N__22305),
            .I(N__22302));
    Odrv12 I__2337 (
            .O(N__22302),
            .I(sbuttonModeStatus_0_sqmuxa_15));
    CascadeMux I__2336 (
            .O(N__22299),
            .I(op_gt_op_gt_un13_striginternallto23_11_cascade_));
    InMux I__2335 (
            .O(N__22296),
            .I(N__22293));
    LocalMux I__2334 (
            .O(N__22293),
            .I(op_gt_op_gt_un13_striginternallto23_16));
    InMux I__2333 (
            .O(N__22290),
            .I(N__22284));
    InMux I__2332 (
            .O(N__22289),
            .I(N__22284));
    LocalMux I__2331 (
            .O(N__22284),
            .I(N__22281));
    Span4Mux_v I__2330 (
            .O(N__22281),
            .I(N__22277));
    InMux I__2329 (
            .O(N__22280),
            .I(N__22274));
    Odrv4 I__2328 (
            .O(N__22277),
            .I(sTrigInternalZ0));
    LocalMux I__2327 (
            .O(N__22274),
            .I(sTrigInternalZ0));
    CascadeMux I__2326 (
            .O(N__22269),
            .I(N__22266));
    InMux I__2325 (
            .O(N__22266),
            .I(N__22263));
    LocalMux I__2324 (
            .O(N__22263),
            .I(op_gt_op_gt_un13_striginternal_0));
    IoInMux I__2323 (
            .O(N__22260),
            .I(N__22257));
    LocalMux I__2322 (
            .O(N__22257),
            .I(N__22254));
    IoSpan4Mux I__2321 (
            .O(N__22254),
            .I(N__22251));
    Span4Mux_s2_h I__2320 (
            .O(N__22251),
            .I(N__22248));
    Sp12to4 I__2319 (
            .O(N__22248),
            .I(N__22245));
    Span12Mux_s11_v I__2318 (
            .O(N__22245),
            .I(N__22242));
    Odrv12 I__2317 (
            .O(N__22242),
            .I(LED_ACQ_obuf_RNOZ0));
    InMux I__2316 (
            .O(N__22239),
            .I(N__22236));
    LocalMux I__2315 (
            .O(N__22236),
            .I(op_gt_op_gt_un13_striginternallto23_18));
    InMux I__2314 (
            .O(N__22233),
            .I(bfn_7_16_0_));
    InMux I__2313 (
            .O(N__22230),
            .I(sCounterRAM_cry_0));
    InMux I__2312 (
            .O(N__22227),
            .I(sCounterRAM_cry_1));
    InMux I__2311 (
            .O(N__22224),
            .I(sCounterRAM_cry_2));
    InMux I__2310 (
            .O(N__22221),
            .I(sCounterRAM_cry_3));
    CascadeMux I__2309 (
            .O(N__22218),
            .I(sbuttonModeStatus_0_sqmuxa_22_cascade_));
    InMux I__2308 (
            .O(N__22215),
            .I(N__22212));
    LocalMux I__2307 (
            .O(N__22212),
            .I(N__22209));
    Span4Mux_v I__2306 (
            .O(N__22209),
            .I(N__22206));
    Span4Mux_v I__2305 (
            .O(N__22206),
            .I(N__22202));
    InMux I__2304 (
            .O(N__22205),
            .I(N__22199));
    Odrv4 I__2303 (
            .O(N__22202),
            .I(sbuttonModeStatusZ0));
    LocalMux I__2302 (
            .O(N__22199),
            .I(sbuttonModeStatusZ0));
    InMux I__2301 (
            .O(N__22194),
            .I(N__22191));
    LocalMux I__2300 (
            .O(N__22191),
            .I(N__22188));
    Odrv12 I__2299 (
            .O(N__22188),
            .I(g1_0_0_3));
    InMux I__2298 (
            .O(N__22185),
            .I(N__22182));
    LocalMux I__2297 (
            .O(N__22182),
            .I(un1_reset_rpi_inv_2_i_o3_16));
    CascadeMux I__2296 (
            .O(N__22179),
            .I(N__22176));
    InMux I__2295 (
            .O(N__22176),
            .I(N__22173));
    LocalMux I__2294 (
            .O(N__22173),
            .I(N__22170));
    Odrv4 I__2293 (
            .O(N__22170),
            .I(g0_2_0_4));
    InMux I__2292 (
            .O(N__22167),
            .I(N__22164));
    LocalMux I__2291 (
            .O(N__22164),
            .I(g2_0_4));
    InMux I__2290 (
            .O(N__22161),
            .I(N__22158));
    LocalMux I__2289 (
            .O(N__22158),
            .I(g2_0_3));
    CascadeMux I__2288 (
            .O(N__22155),
            .I(g1_0_1_1_cascade_));
    InMux I__2287 (
            .O(N__22152),
            .I(N__22149));
    LocalMux I__2286 (
            .O(N__22149),
            .I(g1_0_4));
    CascadeMux I__2285 (
            .O(N__22146),
            .I(N__22143));
    InMux I__2284 (
            .O(N__22143),
            .I(N__22140));
    LocalMux I__2283 (
            .O(N__22140),
            .I(op_gt_op_gt_un13_striginternallto23_13));
    CascadeMux I__2282 (
            .O(N__22137),
            .I(op_gt_op_gt_un13_striginternal_0_cascade_));
    InMux I__2281 (
            .O(N__22134),
            .I(N__22130));
    CascadeMux I__2280 (
            .O(N__22133),
            .I(N__22127));
    LocalMux I__2279 (
            .O(N__22130),
            .I(N__22124));
    InMux I__2278 (
            .O(N__22127),
            .I(N__22121));
    Span4Mux_v I__2277 (
            .O(N__22124),
            .I(N__22118));
    LocalMux I__2276 (
            .O(N__22121),
            .I(N__22115));
    Odrv4 I__2275 (
            .O(N__22118),
            .I(un3_trig_0_4));
    Odrv12 I__2274 (
            .O(N__22115),
            .I(un3_trig_0_4));
    InMux I__2273 (
            .O(N__22110),
            .I(N__22107));
    LocalMux I__2272 (
            .O(N__22107),
            .I(N__22104));
    Odrv12 I__2271 (
            .O(N__22104),
            .I(un1_reset_rpi_inv_2_i_o3_8));
    CascadeMux I__2270 (
            .O(N__22101),
            .I(un1_reset_rpi_inv_2_i_o3_18_cascade_));
    CascadeMux I__2269 (
            .O(N__22098),
            .I(N__22095));
    InMux I__2268 (
            .O(N__22095),
            .I(N__22092));
    LocalMux I__2267 (
            .O(N__22092),
            .I(N__22088));
    CascadeMux I__2266 (
            .O(N__22091),
            .I(N__22085));
    Span4Mux_v I__2265 (
            .O(N__22088),
            .I(N__22082));
    InMux I__2264 (
            .O(N__22085),
            .I(N__22079));
    Span4Mux_h I__2263 (
            .O(N__22082),
            .I(N__22076));
    LocalMux I__2262 (
            .O(N__22079),
            .I(N__22073));
    Odrv4 I__2261 (
            .O(N__22076),
            .I(un3_trig_0_5));
    Odrv12 I__2260 (
            .O(N__22073),
            .I(un3_trig_0_5));
    InMux I__2259 (
            .O(N__22068),
            .I(N__22065));
    LocalMux I__2258 (
            .O(N__22065),
            .I(un1_reset_rpi_inv_2_i_o3_13));
    CascadeMux I__2257 (
            .O(N__22062),
            .I(N__22059));
    InMux I__2256 (
            .O(N__22059),
            .I(N__22056));
    LocalMux I__2255 (
            .O(N__22056),
            .I(g0_2_0_3));
    CascadeMux I__2254 (
            .O(N__22053),
            .I(sTrigInternal_RNIOMLDZ0Z1_cascade_));
    InMux I__2253 (
            .O(N__22050),
            .I(N__22047));
    LocalMux I__2252 (
            .O(N__22047),
            .I(sTrigInternal_RNIOMLDZ0Z1));
    CascadeMux I__2251 (
            .O(N__22044),
            .I(sTrigInternal_RNOZ0Z_0_cascade_));
    InMux I__2250 (
            .O(N__22041),
            .I(N__22037));
    InMux I__2249 (
            .O(N__22040),
            .I(N__22034));
    LocalMux I__2248 (
            .O(N__22037),
            .I(N__22029));
    LocalMux I__2247 (
            .O(N__22034),
            .I(N__22029));
    Odrv4 I__2246 (
            .O(N__22029),
            .I(un3_trig_0));
    CascadeMux I__2245 (
            .O(N__22026),
            .I(sEETrigInternal_prev_RNISEUGZ0_cascade_));
    CascadeMux I__2244 (
            .O(N__22023),
            .I(N__22019));
    InMux I__2243 (
            .O(N__22022),
            .I(N__22014));
    InMux I__2242 (
            .O(N__22019),
            .I(N__22014));
    LocalMux I__2241 (
            .O(N__22014),
            .I(N__22011));
    Odrv12 I__2240 (
            .O(N__22011),
            .I(un3_trig_0_2));
    CascadeMux I__2239 (
            .O(N__22008),
            .I(N__22004));
    InMux I__2238 (
            .O(N__22007),
            .I(N__21999));
    InMux I__2237 (
            .O(N__22004),
            .I(N__21999));
    LocalMux I__2236 (
            .O(N__21999),
            .I(N__21996));
    Odrv4 I__2235 (
            .O(N__21996),
            .I(un3_trig_0_1));
    CascadeMux I__2234 (
            .O(N__21993),
            .I(g1_3_cascade_));
    InMux I__2233 (
            .O(N__21990),
            .I(N__21987));
    LocalMux I__2232 (
            .O(N__21987),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13 ));
    InMux I__2231 (
            .O(N__21984),
            .I(N__21981));
    LocalMux I__2230 (
            .O(N__21981),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1 ));
    InMux I__2229 (
            .O(N__21978),
            .I(N__21975));
    LocalMux I__2228 (
            .O(N__21975),
            .I(N__21972));
    Span4Mux_h I__2227 (
            .O(N__21972),
            .I(N__21969));
    Odrv4 I__2226 (
            .O(N__21969),
            .I(sEESingleContZ0));
    InMux I__2225 (
            .O(N__21966),
            .I(N__21961));
    InMux I__2224 (
            .O(N__21965),
            .I(N__21956));
    InMux I__2223 (
            .O(N__21964),
            .I(N__21956));
    LocalMux I__2222 (
            .O(N__21961),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3 ));
    LocalMux I__2221 (
            .O(N__21956),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3 ));
    InMux I__2220 (
            .O(N__21951),
            .I(N__21943));
    InMux I__2219 (
            .O(N__21950),
            .I(N__21943));
    InMux I__2218 (
            .O(N__21949),
            .I(N__21940));
    InMux I__2217 (
            .O(N__21948),
            .I(N__21937));
    LocalMux I__2216 (
            .O(N__21943),
            .I(\spi_master_inst.sclk_gen_u0.N_1515 ));
    LocalMux I__2215 (
            .O(N__21940),
            .I(\spi_master_inst.sclk_gen_u0.N_1515 ));
    LocalMux I__2214 (
            .O(N__21937),
            .I(\spi_master_inst.sclk_gen_u0.N_1515 ));
    CEMux I__2213 (
            .O(N__21930),
            .I(N__21927));
    LocalMux I__2212 (
            .O(N__21927),
            .I(N__21924));
    Odrv4 I__2211 (
            .O(N__21924),
            .I(sEESingleCont_1_sqmuxa));
    InMux I__2210 (
            .O(N__21921),
            .I(bfn_6_14_0_));
    IoInMux I__2209 (
            .O(N__21918),
            .I(N__21915));
    LocalMux I__2208 (
            .O(N__21915),
            .I(N__21912));
    Span4Mux_s1_h I__2207 (
            .O(N__21912),
            .I(N__21909));
    Span4Mux_h I__2206 (
            .O(N__21909),
            .I(N__21906));
    Span4Mux_h I__2205 (
            .O(N__21906),
            .I(N__21903));
    Odrv4 I__2204 (
            .O(N__21903),
            .I(pon_obuf_RNOZ0));
    InMux I__2203 (
            .O(N__21900),
            .I(N__21897));
    LocalMux I__2202 (
            .O(N__21897),
            .I(N__21894));
    Odrv12 I__2201 (
            .O(N__21894),
            .I(g1_0_5));
    InMux I__2200 (
            .O(N__21891),
            .I(N__21888));
    LocalMux I__2199 (
            .O(N__21888),
            .I(g1));
    InMux I__2198 (
            .O(N__21885),
            .I(N__21882));
    LocalMux I__2197 (
            .O(N__21882),
            .I(sEEPon_i_1));
    InMux I__2196 (
            .O(N__21879),
            .I(N__21876));
    LocalMux I__2195 (
            .O(N__21876),
            .I(N__21873));
    Odrv4 I__2194 (
            .O(N__21873),
            .I(sEEPonZ0Z_2));
    InMux I__2193 (
            .O(N__21870),
            .I(N__21867));
    LocalMux I__2192 (
            .O(N__21867),
            .I(sEEPon_i_2));
    InMux I__2191 (
            .O(N__21864),
            .I(N__21861));
    LocalMux I__2190 (
            .O(N__21861),
            .I(N__21858));
    Odrv4 I__2189 (
            .O(N__21858),
            .I(sEEPonZ0Z_3));
    CascadeMux I__2188 (
            .O(N__21855),
            .I(N__21852));
    InMux I__2187 (
            .O(N__21852),
            .I(N__21849));
    LocalMux I__2186 (
            .O(N__21849),
            .I(sEEPon_i_3));
    InMux I__2185 (
            .O(N__21846),
            .I(N__21843));
    LocalMux I__2184 (
            .O(N__21843),
            .I(N__21840));
    Odrv4 I__2183 (
            .O(N__21840),
            .I(sEEPonZ0Z_4));
    InMux I__2182 (
            .O(N__21837),
            .I(N__21834));
    LocalMux I__2181 (
            .O(N__21834),
            .I(sEEPon_i_4));
    InMux I__2180 (
            .O(N__21831),
            .I(N__21828));
    LocalMux I__2179 (
            .O(N__21828),
            .I(N__21825));
    Odrv4 I__2178 (
            .O(N__21825),
            .I(sEEPonZ0Z_5));
    InMux I__2177 (
            .O(N__21822),
            .I(N__21819));
    LocalMux I__2176 (
            .O(N__21819),
            .I(sEEPon_i_5));
    InMux I__2175 (
            .O(N__21816),
            .I(N__21813));
    LocalMux I__2174 (
            .O(N__21813),
            .I(N__21810));
    Span4Mux_v I__2173 (
            .O(N__21810),
            .I(N__21807));
    Odrv4 I__2172 (
            .O(N__21807),
            .I(sEEPonZ0Z_6));
    InMux I__2171 (
            .O(N__21804),
            .I(N__21801));
    LocalMux I__2170 (
            .O(N__21801),
            .I(sEEPon_i_6));
    InMux I__2169 (
            .O(N__21798),
            .I(N__21795));
    LocalMux I__2168 (
            .O(N__21795),
            .I(N__21792));
    Odrv4 I__2167 (
            .O(N__21792),
            .I(sEEPonZ0Z_7));
    InMux I__2166 (
            .O(N__21789),
            .I(N__21786));
    LocalMux I__2165 (
            .O(N__21786),
            .I(sEEPon_i_7));
    InMux I__2164 (
            .O(N__21783),
            .I(N__21780));
    LocalMux I__2163 (
            .O(N__21780),
            .I(sEEPonPoffZ0Z_1));
    InMux I__2162 (
            .O(N__21777),
            .I(N__21774));
    LocalMux I__2161 (
            .O(N__21774),
            .I(sEEPonPoffZ0Z_2));
    InMux I__2160 (
            .O(N__21771),
            .I(N__21768));
    LocalMux I__2159 (
            .O(N__21768),
            .I(sEEPonPoffZ0Z_3));
    InMux I__2158 (
            .O(N__21765),
            .I(N__21762));
    LocalMux I__2157 (
            .O(N__21762),
            .I(sEEPonPoffZ0Z_4));
    InMux I__2156 (
            .O(N__21759),
            .I(N__21756));
    LocalMux I__2155 (
            .O(N__21756),
            .I(sEEPonPoffZ0Z_5));
    InMux I__2154 (
            .O(N__21753),
            .I(N__21750));
    LocalMux I__2153 (
            .O(N__21750),
            .I(sEEPonPoffZ0Z_6));
    InMux I__2152 (
            .O(N__21747),
            .I(N__21744));
    LocalMux I__2151 (
            .O(N__21744),
            .I(sEEPonPoffZ0Z_7));
    InMux I__2150 (
            .O(N__21741),
            .I(N__21738));
    LocalMux I__2149 (
            .O(N__21738),
            .I(N__21735));
    Odrv12 I__2148 (
            .O(N__21735),
            .I(sEEPonZ0Z_0));
    InMux I__2147 (
            .O(N__21732),
            .I(N__21729));
    LocalMux I__2146 (
            .O(N__21729),
            .I(sEEPon_i_0));
    InMux I__2145 (
            .O(N__21726),
            .I(N__21723));
    LocalMux I__2144 (
            .O(N__21723),
            .I(N__21720));
    Odrv12 I__2143 (
            .O(N__21720),
            .I(sEEPonZ0Z_1));
    InMux I__2142 (
            .O(N__21717),
            .I(N__21714));
    LocalMux I__2141 (
            .O(N__21714),
            .I(sEEPonPoffZ0Z_0));
    InMux I__2140 (
            .O(N__21711),
            .I(N__21708));
    LocalMux I__2139 (
            .O(N__21708),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11 ));
    CascadeMux I__2138 (
            .O(N__21705),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15_cascade_ ));
    CascadeMux I__2137 (
            .O(N__21702),
            .I(N__21697));
    InMux I__2136 (
            .O(N__21701),
            .I(N__21689));
    InMux I__2135 (
            .O(N__21700),
            .I(N__21686));
    InMux I__2134 (
            .O(N__21697),
            .I(N__21683));
    InMux I__2133 (
            .O(N__21696),
            .I(N__21680));
    InMux I__2132 (
            .O(N__21695),
            .I(N__21673));
    InMux I__2131 (
            .O(N__21694),
            .I(N__21673));
    InMux I__2130 (
            .O(N__21693),
            .I(N__21673));
    InMux I__2129 (
            .O(N__21692),
            .I(N__21670));
    LocalMux I__2128 (
            .O(N__21689),
            .I(N__21667));
    LocalMux I__2127 (
            .O(N__21686),
            .I(N__21662));
    LocalMux I__2126 (
            .O(N__21683),
            .I(N__21662));
    LocalMux I__2125 (
            .O(N__21680),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ));
    LocalMux I__2124 (
            .O(N__21673),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ));
    LocalMux I__2123 (
            .O(N__21670),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ));
    Odrv4 I__2122 (
            .O(N__21667),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ));
    Odrv12 I__2121 (
            .O(N__21662),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ));
    InMux I__2120 (
            .O(N__21651),
            .I(N__21648));
    LocalMux I__2119 (
            .O(N__21648),
            .I(N__21645));
    Odrv4 I__2118 (
            .O(N__21645),
            .I(\spi_master_inst.spi_data_path_u1.N_1412 ));
    InMux I__2117 (
            .O(N__21642),
            .I(N__21637));
    InMux I__2116 (
            .O(N__21641),
            .I(N__21634));
    InMux I__2115 (
            .O(N__21640),
            .I(N__21631));
    LocalMux I__2114 (
            .O(N__21637),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3 ));
    LocalMux I__2113 (
            .O(N__21634),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3 ));
    LocalMux I__2112 (
            .O(N__21631),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3 ));
    InMux I__2111 (
            .O(N__21624),
            .I(N__21619));
    InMux I__2110 (
            .O(N__21623),
            .I(N__21616));
    InMux I__2109 (
            .O(N__21622),
            .I(N__21613));
    LocalMux I__2108 (
            .O(N__21619),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1 ));
    LocalMux I__2107 (
            .O(N__21616),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1 ));
    LocalMux I__2106 (
            .O(N__21613),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1 ));
    CascadeMux I__2105 (
            .O(N__21606),
            .I(N__21602));
    InMux I__2104 (
            .O(N__21605),
            .I(N__21598));
    InMux I__2103 (
            .O(N__21602),
            .I(N__21595));
    InMux I__2102 (
            .O(N__21601),
            .I(N__21592));
    LocalMux I__2101 (
            .O(N__21598),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2 ));
    LocalMux I__2100 (
            .O(N__21595),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2 ));
    LocalMux I__2099 (
            .O(N__21592),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2 ));
    InMux I__2098 (
            .O(N__21585),
            .I(N__21581));
    InMux I__2097 (
            .O(N__21584),
            .I(N__21578));
    LocalMux I__2096 (
            .O(N__21581),
            .I(\spi_master_inst.sclk_gen_u0.N_1666 ));
    LocalMux I__2095 (
            .O(N__21578),
            .I(\spi_master_inst.sclk_gen_u0.N_1666 ));
    CascadeMux I__2094 (
            .O(N__21573),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3_cascade_ ));
    InMux I__2093 (
            .O(N__21570),
            .I(N__21565));
    InMux I__2092 (
            .O(N__21569),
            .I(N__21562));
    InMux I__2091 (
            .O(N__21568),
            .I(N__21559));
    LocalMux I__2090 (
            .O(N__21565),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0 ));
    LocalMux I__2089 (
            .O(N__21562),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0 ));
    LocalMux I__2088 (
            .O(N__21559),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0 ));
    CascadeMux I__2087 (
            .O(N__21552),
            .I(\spi_master_inst.sclk_gen_u0.N_1515_cascade_ ));
    CascadeMux I__2086 (
            .O(N__21549),
            .I(\spi_master_inst.sclk_gen_u0.N_36_cascade_ ));
    InMux I__2085 (
            .O(N__21546),
            .I(N__21543));
    LocalMux I__2084 (
            .O(N__21543),
            .I(\spi_master_inst.sclk_gen_u0.N_48 ));
    CascadeMux I__2083 (
            .O(N__21540),
            .I(\spi_master_inst.sclk_gen_u0.N_5_cascade_ ));
    InMux I__2082 (
            .O(N__21537),
            .I(N__21533));
    InMux I__2081 (
            .O(N__21536),
            .I(N__21530));
    LocalMux I__2080 (
            .O(N__21533),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_start_iZ0 ));
    LocalMux I__2079 (
            .O(N__21530),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_start_iZ0 ));
    CascadeMux I__2078 (
            .O(N__21525),
            .I(N__21521));
    InMux I__2077 (
            .O(N__21524),
            .I(N__21517));
    InMux I__2076 (
            .O(N__21521),
            .I(N__21512));
    InMux I__2075 (
            .O(N__21520),
            .I(N__21512));
    LocalMux I__2074 (
            .O(N__21517),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1 ));
    LocalMux I__2073 (
            .O(N__21512),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1 ));
    InMux I__2072 (
            .O(N__21507),
            .I(N__21504));
    LocalMux I__2071 (
            .O(N__21504),
            .I(\spi_master_inst.spi_data_path_u1.N_1415 ));
    InMux I__2070 (
            .O(N__21501),
            .I(N__21498));
    LocalMux I__2069 (
            .O(N__21498),
            .I(N__21495));
    Span4Mux_h I__2068 (
            .O(N__21495),
            .I(N__21492));
    Odrv4 I__2067 (
            .O(N__21492),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6 ));
    CascadeMux I__2066 (
            .O(N__21489),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14_cascade_ ));
    InMux I__2065 (
            .O(N__21486),
            .I(N__21483));
    LocalMux I__2064 (
            .O(N__21483),
            .I(\spi_master_inst.spi_data_path_u1.N_1419 ));
    CascadeMux I__2063 (
            .O(N__21480),
            .I(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_ ));
    InMux I__2062 (
            .O(N__21477),
            .I(N__21474));
    LocalMux I__2061 (
            .O(N__21474),
            .I(\spi_master_inst.spi_data_path_u1.N_1422 ));
    InMux I__2060 (
            .O(N__21471),
            .I(N__21465));
    InMux I__2059 (
            .O(N__21470),
            .I(N__21465));
    LocalMux I__2058 (
            .O(N__21465),
            .I(\spi_master_inst.sclk_gen_u0.N_1520 ));
    InMux I__2057 (
            .O(N__21462),
            .I(N__21444));
    InMux I__2056 (
            .O(N__21461),
            .I(N__21444));
    InMux I__2055 (
            .O(N__21460),
            .I(N__21444));
    InMux I__2054 (
            .O(N__21459),
            .I(N__21444));
    InMux I__2053 (
            .O(N__21458),
            .I(N__21444));
    InMux I__2052 (
            .O(N__21457),
            .I(N__21437));
    InMux I__2051 (
            .O(N__21456),
            .I(N__21437));
    InMux I__2050 (
            .O(N__21455),
            .I(N__21437));
    LocalMux I__2049 (
            .O(N__21444),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_start_i_i ));
    LocalMux I__2048 (
            .O(N__21437),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_start_i_i ));
    InMux I__2047 (
            .O(N__21432),
            .I(bfn_5_13_0_));
    InMux I__2046 (
            .O(N__21429),
            .I(N__21426));
    LocalMux I__2045 (
            .O(N__21426),
            .I(\spi_master_inst.spi_data_path_u1.N_1423 ));
    InMux I__2044 (
            .O(N__21423),
            .I(N__21417));
    InMux I__2043 (
            .O(N__21422),
            .I(N__21417));
    LocalMux I__2042 (
            .O(N__21417),
            .I(N__21413));
    CascadeMux I__2041 (
            .O(N__21416),
            .I(N__21410));
    Span4Mux_v I__2040 (
            .O(N__21413),
            .I(N__21405));
    InMux I__2039 (
            .O(N__21410),
            .I(N__21402));
    InMux I__2038 (
            .O(N__21409),
            .I(N__21399));
    InMux I__2037 (
            .O(N__21408),
            .I(N__21396));
    Odrv4 I__2036 (
            .O(N__21405),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1 ));
    LocalMux I__2035 (
            .O(N__21402),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1 ));
    LocalMux I__2034 (
            .O(N__21399),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1 ));
    LocalMux I__2033 (
            .O(N__21396),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1 ));
    CascadeMux I__2032 (
            .O(N__21387),
            .I(N__21384));
    InMux I__2031 (
            .O(N__21384),
            .I(N__21381));
    LocalMux I__2030 (
            .O(N__21381),
            .I(\spi_master_inst.spi_data_path_u1.N_1416 ));
    InMux I__2029 (
            .O(N__21378),
            .I(N__21375));
    LocalMux I__2028 (
            .O(N__21375),
            .I(sEEPonPoff_i_0));
    InMux I__2027 (
            .O(N__21372),
            .I(N__21369));
    LocalMux I__2026 (
            .O(N__21369),
            .I(sEEPonPoff_i_1));
    InMux I__2025 (
            .O(N__21366),
            .I(N__21363));
    LocalMux I__2024 (
            .O(N__21363),
            .I(sEEPonPoff_i_2));
    CascadeMux I__2023 (
            .O(N__21360),
            .I(N__21357));
    InMux I__2022 (
            .O(N__21357),
            .I(N__21354));
    LocalMux I__2021 (
            .O(N__21354),
            .I(sEEPonPoff_i_3));
    InMux I__2020 (
            .O(N__21351),
            .I(N__21348));
    LocalMux I__2019 (
            .O(N__21348),
            .I(sEEPonPoff_i_4));
    CascadeMux I__2018 (
            .O(N__21345),
            .I(N__21342));
    InMux I__2017 (
            .O(N__21342),
            .I(N__21339));
    LocalMux I__2016 (
            .O(N__21339),
            .I(sEEPonPoff_i_5));
    InMux I__2015 (
            .O(N__21336),
            .I(N__21333));
    LocalMux I__2014 (
            .O(N__21333),
            .I(sEEPonPoff_i_6));
    InMux I__2013 (
            .O(N__21330),
            .I(N__21327));
    LocalMux I__2012 (
            .O(N__21327),
            .I(sEEPonPoff_i_7));
    CascadeMux I__2011 (
            .O(N__21324),
            .I(\spi_master_inst.sclk_gen_u0.N_1666_cascade_ ));
    InMux I__2010 (
            .O(N__21321),
            .I(N__21318));
    LocalMux I__2009 (
            .O(N__21318),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4 ));
    InMux I__2008 (
            .O(N__21315),
            .I(N__21309));
    InMux I__2007 (
            .O(N__21314),
            .I(N__21309));
    LocalMux I__2006 (
            .O(N__21309),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0 ));
    CascadeMux I__2005 (
            .O(N__21306),
            .I(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_ ));
    CascadeMux I__2004 (
            .O(N__21303),
            .I(\spi_master_inst.sclk_gen_u0.N_48_cascade_ ));
    InMux I__2003 (
            .O(N__21300),
            .I(N__21293));
    InMux I__2002 (
            .O(N__21299),
            .I(N__21290));
    CascadeMux I__2001 (
            .O(N__21298),
            .I(N__21287));
    InMux I__2000 (
            .O(N__21297),
            .I(N__21284));
    InMux I__1999 (
            .O(N__21296),
            .I(N__21281));
    LocalMux I__1998 (
            .O(N__21293),
            .I(N__21278));
    LocalMux I__1997 (
            .O(N__21290),
            .I(N__21275));
    InMux I__1996 (
            .O(N__21287),
            .I(N__21272));
    LocalMux I__1995 (
            .O(N__21284),
            .I(N__21265));
    LocalMux I__1994 (
            .O(N__21281),
            .I(N__21265));
    Span4Mux_h I__1993 (
            .O(N__21278),
            .I(N__21265));
    Span4Mux_h I__1992 (
            .O(N__21275),
            .I(N__21262));
    LocalMux I__1991 (
            .O(N__21272),
            .I(\spi_master_inst.ss_start_i ));
    Odrv4 I__1990 (
            .O(N__21265),
            .I(\spi_master_inst.ss_start_i ));
    Odrv4 I__1989 (
            .O(N__21262),
            .I(\spi_master_inst.ss_start_i ));
    InMux I__1988 (
            .O(N__21255),
            .I(bfn_5_5_0_));
    InMux I__1987 (
            .O(N__21252),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_0 ));
    InMux I__1986 (
            .O(N__21249),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_1 ));
    InMux I__1985 (
            .O(N__21246),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_2 ));
    InMux I__1984 (
            .O(N__21243),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_3 ));
    InMux I__1983 (
            .O(N__21240),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_4 ));
    InMux I__1982 (
            .O(N__21237),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_5 ));
    InMux I__1981 (
            .O(N__21234),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_6 ));
    InMux I__1980 (
            .O(N__21231),
            .I(N__21227));
    InMux I__1979 (
            .O(N__21230),
            .I(N__21224));
    LocalMux I__1978 (
            .O(N__21227),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6 ));
    LocalMux I__1977 (
            .O(N__21224),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6 ));
    InMux I__1976 (
            .O(N__21219),
            .I(N__21215));
    InMux I__1975 (
            .O(N__21218),
            .I(N__21212));
    LocalMux I__1974 (
            .O(N__21215),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5 ));
    LocalMux I__1973 (
            .O(N__21212),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5 ));
    CascadeMux I__1972 (
            .O(N__21207),
            .I(N__21203));
    InMux I__1971 (
            .O(N__21206),
            .I(N__21200));
    InMux I__1970 (
            .O(N__21203),
            .I(N__21197));
    LocalMux I__1969 (
            .O(N__21200),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7 ));
    LocalMux I__1968 (
            .O(N__21197),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7 ));
    InMux I__1967 (
            .O(N__21192),
            .I(N__21188));
    InMux I__1966 (
            .O(N__21191),
            .I(N__21185));
    LocalMux I__1965 (
            .O(N__21188),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4 ));
    LocalMux I__1964 (
            .O(N__21185),
            .I(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4 ));
    InMux I__1963 (
            .O(N__21180),
            .I(N__21177));
    LocalMux I__1962 (
            .O(N__21177),
            .I(N__21173));
    CascadeMux I__1961 (
            .O(N__21176),
            .I(N__21169));
    Span4Mux_v I__1960 (
            .O(N__21173),
            .I(N__21165));
    InMux I__1959 (
            .O(N__21172),
            .I(N__21162));
    InMux I__1958 (
            .O(N__21169),
            .I(N__21159));
    InMux I__1957 (
            .O(N__21168),
            .I(N__21156));
    Odrv4 I__1956 (
            .O(N__21165),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0 ));
    LocalMux I__1955 (
            .O(N__21162),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0 ));
    LocalMux I__1954 (
            .O(N__21159),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0 ));
    LocalMux I__1953 (
            .O(N__21156),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0 ));
    IoInMux I__1952 (
            .O(N__21147),
            .I(N__21144));
    LocalMux I__1951 (
            .O(N__21144),
            .I(N__21141));
    Span4Mux_s0_v I__1950 (
            .O(N__21141),
            .I(N__21138));
    Span4Mux_v I__1949 (
            .O(N__21138),
            .I(N__21135));
    Span4Mux_v I__1948 (
            .O(N__21135),
            .I(N__21132));
    Odrv4 I__1947 (
            .O(N__21132),
            .I(DAC_mosi_c));
    InMux I__1946 (
            .O(N__21129),
            .I(N__21126));
    LocalMux I__1945 (
            .O(N__21126),
            .I(N__21123));
    Span4Mux_h I__1944 (
            .O(N__21123),
            .I(N__21120));
    Odrv4 I__1943 (
            .O(N__21120),
            .I(\spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1 ));
    InMux I__1942 (
            .O(N__21117),
            .I(N__21114));
    LocalMux I__1941 (
            .O(N__21114),
            .I(N__21111));
    Span4Mux_v I__1940 (
            .O(N__21111),
            .I(N__21106));
    InMux I__1939 (
            .O(N__21110),
            .I(N__21103));
    InMux I__1938 (
            .O(N__21109),
            .I(N__21100));
    Odrv4 I__1937 (
            .O(N__21106),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5 ));
    LocalMux I__1936 (
            .O(N__21103),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5 ));
    LocalMux I__1935 (
            .O(N__21100),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5 ));
    InMux I__1934 (
            .O(N__21093),
            .I(N__21090));
    LocalMux I__1933 (
            .O(N__21090),
            .I(N__21087));
    Span4Mux_v I__1932 (
            .O(N__21087),
            .I(N__21082));
    InMux I__1931 (
            .O(N__21086),
            .I(N__21079));
    InMux I__1930 (
            .O(N__21085),
            .I(N__21076));
    Odrv4 I__1929 (
            .O(N__21082),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4 ));
    LocalMux I__1928 (
            .O(N__21079),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4 ));
    LocalMux I__1927 (
            .O(N__21076),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4 ));
    IoInMux I__1926 (
            .O(N__21069),
            .I(N__21066));
    LocalMux I__1925 (
            .O(N__21066),
            .I(N__21063));
    Span4Mux_s1_v I__1924 (
            .O(N__21063),
            .I(N__21060));
    Span4Mux_v I__1923 (
            .O(N__21060),
            .I(N__21056));
    InMux I__1922 (
            .O(N__21059),
            .I(N__21053));
    Span4Mux_v I__1921 (
            .O(N__21056),
            .I(N__21050));
    LocalMux I__1920 (
            .O(N__21053),
            .I(N__21047));
    Span4Mux_h I__1919 (
            .O(N__21050),
            .I(N__21042));
    Span4Mux_v I__1918 (
            .O(N__21047),
            .I(N__21042));
    Odrv4 I__1917 (
            .O(N__21042),
            .I(DAC_sclk_c));
    InMux I__1916 (
            .O(N__21039),
            .I(N__21036));
    LocalMux I__1915 (
            .O(N__21036),
            .I(N__21033));
    Odrv4 I__1914 (
            .O(N__21033),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO ));
    InMux I__1913 (
            .O(N__21030),
            .I(N__21023));
    InMux I__1912 (
            .O(N__21029),
            .I(N__21018));
    InMux I__1911 (
            .O(N__21028),
            .I(N__21018));
    InMux I__1910 (
            .O(N__21027),
            .I(N__21015));
    InMux I__1909 (
            .O(N__21026),
            .I(N__21012));
    LocalMux I__1908 (
            .O(N__21023),
            .I(N__21007));
    LocalMux I__1907 (
            .O(N__21018),
            .I(N__21007));
    LocalMux I__1906 (
            .O(N__21015),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6 ));
    LocalMux I__1905 (
            .O(N__21012),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6 ));
    Odrv4 I__1904 (
            .O(N__21007),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6 ));
    CascadeMux I__1903 (
            .O(N__21000),
            .I(N__20996));
    InMux I__1902 (
            .O(N__20999),
            .I(N__20987));
    InMux I__1901 (
            .O(N__20996),
            .I(N__20987));
    InMux I__1900 (
            .O(N__20995),
            .I(N__20987));
    CascadeMux I__1899 (
            .O(N__20994),
            .I(N__20981));
    LocalMux I__1898 (
            .O(N__20987),
            .I(N__20978));
    InMux I__1897 (
            .O(N__20986),
            .I(N__20975));
    CEMux I__1896 (
            .O(N__20985),
            .I(N__20972));
    InMux I__1895 (
            .O(N__20984),
            .I(N__20967));
    InMux I__1894 (
            .O(N__20981),
            .I(N__20967));
    Span4Mux_v I__1893 (
            .O(N__20978),
            .I(N__20964));
    LocalMux I__1892 (
            .O(N__20975),
            .I(N__20961));
    LocalMux I__1891 (
            .O(N__20972),
            .I(\spi_master_inst.o_sclk_RNIH6AC ));
    LocalMux I__1890 (
            .O(N__20967),
            .I(\spi_master_inst.o_sclk_RNIH6AC ));
    Odrv4 I__1889 (
            .O(N__20964),
            .I(\spi_master_inst.o_sclk_RNIH6AC ));
    Odrv4 I__1888 (
            .O(N__20961),
            .I(\spi_master_inst.o_sclk_RNIH6AC ));
    InMux I__1887 (
            .O(N__20952),
            .I(N__20949));
    LocalMux I__1886 (
            .O(N__20949),
            .I(N__20946));
    Odrv4 I__1885 (
            .O(N__20946),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO ));
    InMux I__1884 (
            .O(N__20943),
            .I(N__20940));
    LocalMux I__1883 (
            .O(N__20940),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO ));
    InMux I__1882 (
            .O(N__20937),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0 ));
    InMux I__1881 (
            .O(N__20934),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1 ));
    InMux I__1880 (
            .O(N__20931),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2 ));
    InMux I__1879 (
            .O(N__20928),
            .I(N__20924));
    InMux I__1878 (
            .O(N__20927),
            .I(N__20921));
    LocalMux I__1877 (
            .O(N__20924),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4 ));
    LocalMux I__1876 (
            .O(N__20921),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4 ));
    InMux I__1875 (
            .O(N__20916),
            .I(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3 ));
    InMux I__1874 (
            .O(N__20913),
            .I(bfn_3_5_0_));
    CascadeMux I__1873 (
            .O(N__20910),
            .I(N__20906));
    InMux I__1872 (
            .O(N__20909),
            .I(N__20903));
    InMux I__1871 (
            .O(N__20906),
            .I(N__20900));
    LocalMux I__1870 (
            .O(N__20903),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5 ));
    LocalMux I__1869 (
            .O(N__20900),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5 ));
    InMux I__1868 (
            .O(N__20895),
            .I(bfn_3_3_0_));
    CascadeMux I__1867 (
            .O(N__20892),
            .I(N__20889));
    InMux I__1866 (
            .O(N__20889),
            .I(N__20885));
    InMux I__1865 (
            .O(N__20888),
            .I(N__20882));
    LocalMux I__1864 (
            .O(N__20885),
            .I(N__20879));
    LocalMux I__1863 (
            .O(N__20882),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1 ));
    Odrv12 I__1862 (
            .O(N__20879),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1 ));
    InMux I__1861 (
            .O(N__20874),
            .I(N__20871));
    LocalMux I__1860 (
            .O(N__20871),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_s_1 ));
    InMux I__1859 (
            .O(N__20868),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0 ));
    InMux I__1858 (
            .O(N__20865),
            .I(N__20860));
    InMux I__1857 (
            .O(N__20864),
            .I(N__20857));
    InMux I__1856 (
            .O(N__20863),
            .I(N__20854));
    LocalMux I__1855 (
            .O(N__20860),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2 ));
    LocalMux I__1854 (
            .O(N__20857),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2 ));
    LocalMux I__1853 (
            .O(N__20854),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2 ));
    InMux I__1852 (
            .O(N__20847),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1 ));
    CascadeMux I__1851 (
            .O(N__20844),
            .I(N__20841));
    InMux I__1850 (
            .O(N__20841),
            .I(N__20836));
    InMux I__1849 (
            .O(N__20840),
            .I(N__20833));
    InMux I__1848 (
            .O(N__20839),
            .I(N__20830));
    LocalMux I__1847 (
            .O(N__20836),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3 ));
    LocalMux I__1846 (
            .O(N__20833),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3 ));
    LocalMux I__1845 (
            .O(N__20830),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3 ));
    InMux I__1844 (
            .O(N__20823),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2 ));
    InMux I__1843 (
            .O(N__20820),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3 ));
    InMux I__1842 (
            .O(N__20817),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4 ));
    InMux I__1841 (
            .O(N__20814),
            .I(N__20809));
    InMux I__1840 (
            .O(N__20813),
            .I(N__20806));
    InMux I__1839 (
            .O(N__20812),
            .I(N__20803));
    LocalMux I__1838 (
            .O(N__20809),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6 ));
    LocalMux I__1837 (
            .O(N__20806),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6 ));
    LocalMux I__1836 (
            .O(N__20803),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6 ));
    InMux I__1835 (
            .O(N__20796),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5 ));
    InMux I__1834 (
            .O(N__20793),
            .I(N__20779));
    InMux I__1833 (
            .O(N__20792),
            .I(N__20779));
    InMux I__1832 (
            .O(N__20791),
            .I(N__20779));
    InMux I__1831 (
            .O(N__20790),
            .I(N__20774));
    InMux I__1830 (
            .O(N__20789),
            .I(N__20774));
    InMux I__1829 (
            .O(N__20788),
            .I(N__20767));
    InMux I__1828 (
            .O(N__20787),
            .I(N__20767));
    InMux I__1827 (
            .O(N__20786),
            .I(N__20767));
    LocalMux I__1826 (
            .O(N__20779),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i ));
    LocalMux I__1825 (
            .O(N__20774),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i ));
    LocalMux I__1824 (
            .O(N__20767),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i ));
    InMux I__1823 (
            .O(N__20760),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6 ));
    CascadeMux I__1822 (
            .O(N__20757),
            .I(N__20752));
    InMux I__1821 (
            .O(N__20756),
            .I(N__20749));
    InMux I__1820 (
            .O(N__20755),
            .I(N__20746));
    InMux I__1819 (
            .O(N__20752),
            .I(N__20743));
    LocalMux I__1818 (
            .O(N__20749),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7 ));
    LocalMux I__1817 (
            .O(N__20746),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7 ));
    LocalMux I__1816 (
            .O(N__20743),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7 ));
    InMux I__1815 (
            .O(N__20736),
            .I(N__20732));
    InMux I__1814 (
            .O(N__20735),
            .I(N__20729));
    LocalMux I__1813 (
            .O(N__20732),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2 ));
    LocalMux I__1812 (
            .O(N__20729),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2 ));
    InMux I__1811 (
            .O(N__20724),
            .I(sRAM_pointer_read_cry_11));
    InMux I__1810 (
            .O(N__20721),
            .I(sRAM_pointer_read_cry_12));
    InMux I__1809 (
            .O(N__20718),
            .I(sRAM_pointer_read_cry_13));
    InMux I__1808 (
            .O(N__20715),
            .I(sRAM_pointer_read_cry_14));
    InMux I__1807 (
            .O(N__20712),
            .I(bfn_2_13_0_));
    InMux I__1806 (
            .O(N__20709),
            .I(sRAM_pointer_read_cry_16));
    InMux I__1805 (
            .O(N__20706),
            .I(sRAM_pointer_read_cry_17));
    CEMux I__1804 (
            .O(N__20703),
            .I(N__20694));
    CEMux I__1803 (
            .O(N__20702),
            .I(N__20694));
    CEMux I__1802 (
            .O(N__20701),
            .I(N__20694));
    GlobalMux I__1801 (
            .O(N__20694),
            .I(N__20691));
    gio2CtrlBuf I__1800 (
            .O(N__20691),
            .I(N_28_g));
    InMux I__1799 (
            .O(N__20688),
            .I(N__20685));
    LocalMux I__1798 (
            .O(N__20685),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0 ));
    CascadeMux I__1797 (
            .O(N__20682),
            .I(N__20679));
    InMux I__1796 (
            .O(N__20679),
            .I(N__20676));
    LocalMux I__1795 (
            .O(N__20676),
            .I(\spi_master_inst.sclk_gen_u0.sclk_count_i_s_0 ));
    InMux I__1794 (
            .O(N__20673),
            .I(sRAM_pointer_read_cry_1));
    InMux I__1793 (
            .O(N__20670),
            .I(sRAM_pointer_read_cry_2));
    InMux I__1792 (
            .O(N__20667),
            .I(sRAM_pointer_read_cry_3));
    InMux I__1791 (
            .O(N__20664),
            .I(sRAM_pointer_read_cry_4));
    InMux I__1790 (
            .O(N__20661),
            .I(sRAM_pointer_read_cry_5));
    InMux I__1789 (
            .O(N__20658),
            .I(sRAM_pointer_read_cry_6));
    InMux I__1788 (
            .O(N__20655),
            .I(bfn_2_12_0_));
    InMux I__1787 (
            .O(N__20652),
            .I(sRAM_pointer_read_cry_8));
    InMux I__1786 (
            .O(N__20649),
            .I(sRAM_pointer_read_cry_9));
    InMux I__1785 (
            .O(N__20646),
            .I(sRAM_pointer_read_cry_10));
    InMux I__1784 (
            .O(N__20643),
            .I(N__20640));
    LocalMux I__1783 (
            .O(N__20640),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3 ));
    CascadeMux I__1782 (
            .O(N__20637),
            .I(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3_cascade_ ));
    InMux I__1781 (
            .O(N__20634),
            .I(N__20631));
    LocalMux I__1780 (
            .O(N__20631),
            .I(\spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1 ));
    InMux I__1779 (
            .O(N__20628),
            .I(N__20622));
    InMux I__1778 (
            .O(N__20627),
            .I(N__20622));
    LocalMux I__1777 (
            .O(N__20622),
            .I(\spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i ));
    CascadeMux I__1776 (
            .O(N__20619),
            .I(\spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i_cascade_ ));
    InMux I__1775 (
            .O(N__20616),
            .I(bfn_2_11_0_));
    InMux I__1774 (
            .O(N__20613),
            .I(sRAM_pointer_read_cry_0));
    InMux I__1773 (
            .O(N__20610),
            .I(N__20607));
    LocalMux I__1772 (
            .O(N__20607),
            .I(N__20604));
    Span4Mux_v I__1771 (
            .O(N__20604),
            .I(N__20601));
    Span4Mux_h I__1770 (
            .O(N__20601),
            .I(N__20598));
    Odrv4 I__1769 (
            .O(N__20598),
            .I(button_mode_c));
    IoInMux I__1768 (
            .O(N__20595),
            .I(N__20592));
    LocalMux I__1767 (
            .O(N__20592),
            .I(N__20589));
    Span4Mux_s0_h I__1766 (
            .O(N__20589),
            .I(N__20586));
    Span4Mux_v I__1765 (
            .O(N__20586),
            .I(N__20583));
    Span4Mux_v I__1764 (
            .O(N__20583),
            .I(N__20580));
    Span4Mux_h I__1763 (
            .O(N__20580),
            .I(N__20577));
    Odrv4 I__1762 (
            .O(N__20577),
            .I(button_mode_ibuf_RNIN5KZ0Z7));
    IoInMux I__1761 (
            .O(N__20574),
            .I(N__20571));
    LocalMux I__1760 (
            .O(N__20571),
            .I(N__20568));
    Span12Mux_s7_v I__1759 (
            .O(N__20568),
            .I(N__20565));
    Odrv12 I__1758 (
            .O(N__20565),
            .I(DAC_cs_c));
    IoInMux I__1757 (
            .O(N__20562),
            .I(N__20559));
    LocalMux I__1756 (
            .O(N__20559),
            .I(N__20556));
    Span4Mux_s0_h I__1755 (
            .O(N__20556),
            .I(N__20553));
    Span4Mux_h I__1754 (
            .O(N__20553),
            .I(N__20550));
    Sp12to4 I__1753 (
            .O(N__20550),
            .I(N__20547));
    Span12Mux_v I__1752 (
            .O(N__20547),
            .I(N__20544));
    Span12Mux_h I__1751 (
            .O(N__20544),
            .I(N__20541));
    Odrv12 I__1750 (
            .O(N__20541),
            .I(\pll128M2_inst.pll_clk128 ));
    IoInMux I__1749 (
            .O(N__20538),
            .I(N__20535));
    LocalMux I__1748 (
            .O(N__20535),
            .I(N__20532));
    Span4Mux_s3_v I__1747 (
            .O(N__20532),
            .I(N__20529));
    Sp12to4 I__1746 (
            .O(N__20529),
            .I(N__20526));
    Span12Mux_h I__1745 (
            .O(N__20526),
            .I(N__20523));
    Span12Mux_v I__1744 (
            .O(N__20523),
            .I(N__20520));
    Odrv12 I__1743 (
            .O(N__20520),
            .I(clk_c));
    IoInMux I__1742 (
            .O(N__20517),
            .I(N__20514));
    LocalMux I__1741 (
            .O(N__20514),
            .I(N__20511));
    Odrv4 I__1740 (
            .O(N__20511),
            .I(\pll128M2_inst.pll_clk64_0 ));
    INV \INVspi_slave_inst.tx_data_count_neg_sclk_i_0C  (
            .O(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .I(N__30702));
    INV \INVspi_slave_inst.tx_done_neg_sclk_iC  (
            .O(\INVspi_slave_inst.tx_done_neg_sclk_iC_net ),
            .I(N__30701));
    INV \INVspi_slave_inst.rx_done_neg_sclk_iC  (
            .O(\INVspi_slave_inst.rx_done_neg_sclk_iC_net ),
            .I(N__30699));
    INV \INVspi_slave_inst.rx_data_count_neg_sclk_i_0C  (
            .O(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .I(N__30698));
    defparam IN_MUX_bfv_22_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_10_0_));
    defparam IN_MUX_bfv_22_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_11_0_ (
            .carryinitin(un2_scounterdac_cry_8),
            .carryinitout(bfn_22_11_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(un1_sacqtime_cry_7),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(un1_sacqtime_cry_15),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(un1_sacqtime_cry_23),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_9_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_3_0_));
    defparam IN_MUX_bfv_3_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_4_0_));
    defparam IN_MUX_bfv_3_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_5_0_ (
            .carryinitin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO ),
            .carryinitout(bfn_3_5_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_6_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_12_0_ (
            .carryinitin(un7_spon_cry_7),
            .carryinitout(bfn_6_12_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(un7_spon_cry_15),
            .carryinitout(bfn_6_13_0_));
    defparam IN_MUX_bfv_6_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_14_0_ (
            .carryinitin(un7_spon_cry_23),
            .carryinitout(bfn_6_14_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(un5_sdacdyn_cry_7),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(un5_sdacdyn_cry_15),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(un5_sdacdyn_cry_23),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(un4_spoff_cry_7),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(un4_spoff_cry_15),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(un4_spoff_cry_23),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(un4_speriod_cry_7),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(un4_speriod_cry_15),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(un4_speriod_cry_23),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(un4_sacqtime_cry_7),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(un4_sacqtime_cry_15),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(un4_sacqtime_cry_23),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(un1_spoff_cry_7),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(un1_spoff_cry_15),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(un1_spoff_cry_23),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(un10_trig_prev_cry_7),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_15_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_2_0_));
    defparam IN_MUX_bfv_10_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_2_0_));
    defparam IN_MUX_bfv_3_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_3_0_));
    defparam IN_MUX_bfv_5_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_5_0_));
    defparam IN_MUX_bfv_10_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_6_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(un1_button_debounce_counter_cry_8),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(un1_button_debounce_counter_cry_16),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(sRAM_pointer_write_cry_7),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(sRAM_pointer_write_cry_15),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(sRAM_pointer_read_cry_7),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(sRAM_pointer_read_cry_15),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(sCounter_cry_7),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(sCounter_cry_15),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_15_0_));
    ICE_GB reset_rpi_ibuf_RNIIUT3_0 (
            .USERSIGNALTOGLOBALBUFFER(N__27288),
            .GLOBALBUFFEROUTPUT(LED3_c_i_g));
    ICE_GB sEEPointerReset_RNI2CQM_0 (
            .USERSIGNALTOGLOBALBUFFER(N__26601),
            .GLOBALBUFFEROUTPUT(N_26_g));
    ICE_GB \pll128M2_inst.PLLOUTCOREB_derived_clock_RNI5L14  (
            .USERSIGNALTOGLOBALBUFFER(N__20517),
            .GLOBALBUFFEROUTPUT(pll_clk64_0_g));
    ICE_GB spi_sclk_inferred_clock_RNIH8F3 (
            .USERSIGNALTOGLOBALBUFFER(N__28701),
            .GLOBALBUFFEROUTPUT(spi_sclk_g));
    ICE_GB sEEPointerReset_RNILL2C1_0 (
            .USERSIGNALTOGLOBALBUFFER(N__27849),
            .GLOBALBUFFEROUTPUT(N_28_g));
    ICE_GB \pll128M2_inst.PLLOUTCOREA_derived_clock_RNI4765  (
            .USERSIGNALTOGLOBALBUFFER(N__20562),
            .GLOBALBUFFEROUTPUT(pll_clk128_g));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB sCounterDAC_RNIBR1C_0_0 (
            .USERSIGNALTOGLOBALBUFFER(N__53346),
            .GLOBALBUFFEROUTPUT(op_eq_scounterdac10_g));
    ICE_GB button_mode_ibuf_RNIN5K7_0 (
            .USERSIGNALTOGLOBALBUFFER(N__20595),
            .GLOBALBUFFEROUTPUT(N_3089_g));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam button_mode_ibuf_RNIN5K7_LC_1_19_4.C_ON=1'b0;
    defparam button_mode_ibuf_RNIN5K7_LC_1_19_4.SEQ_MODE=4'b0000;
    defparam button_mode_ibuf_RNIN5K7_LC_1_19_4.LUT_INIT=16'b0000000010101010;
    LogicCell40 button_mode_ibuf_RNIN5K7_LC_1_19_4 (
            .in0(N__32691),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20610),
            .lcout(button_mode_ibuf_RNIN5KZ0Z7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.o_slave_csn_0_LC_2_2_6 .C_ON=1'b0;
    defparam \spi_master_inst.o_slave_csn_0_LC_2_2_6 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.o_slave_csn_0_LC_2_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.o_slave_csn_0_LC_2_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21300),
            .lcout(DAC_cs_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53259),
            .ce(),
            .sr(N__53148));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIIUTC1_7_LC_2_3_0 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIIUTC1_7_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIIUTC1_7_LC_2_3_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIIUTC1_7_LC_2_3_0  (
            .in0(N__20812),
            .in1(N__21109),
            .in2(N__20757),
            .in3(N__21085),
            .lcout(\spi_master_inst.sclk_gen_u0.un1_sclk_count_start_ilto7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_1_LC_2_3_3 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_1_LC_2_3_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_1_LC_2_3_3 .LUT_INIT=16'b1100111110101010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_1_LC_2_3_3  (
            .in0(N__20874),
            .in1(N__20628),
            .in2(N__22536),
            .in3(N__20790),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53265),
            .ce(),
            .sr(N__53147));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_0_LC_2_3_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_0_LC_2_3_7 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_0_LC_2_3_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_0_LC_2_3_7  (
            .in0(N__22532),
            .in1(N__20627),
            .in2(N__20682),
            .in3(N__20789),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53265),
            .ce(),
            .sr(N__53147));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52_2_LC_2_4_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52_2_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52_2_LC_2_4_0 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52_2_LC_2_4_0  (
            .in0(N__22637),
            .in1(N__21299),
            .in2(N__21702),
            .in3(N__20643),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIGUQ52Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_RNI06S51_5_LC_2_4_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_RNI06S51_5_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_RNI06S51_5_LC_2_4_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_RNI06S51_5_LC_2_4_1  (
            .in0(N__20927),
            .in1(N__21408),
            .in2(N__20910),
            .in3(N__21168),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3 ),
            .ltout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIL1LO1_2_LC_2_4_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIL1LO1_2_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIL1LO1_2_LC_2_4_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIL1LO1_2_LC_2_4_2  (
            .in0(N__22638),
            .in1(_gnd_net_),
            .in2(N__20637),
            .in3(N__21700),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIL2KE2_1_LC_2_4_6 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIL2KE2_1_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIL2KE2_1_LC_2_4_6 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_RNIL2KE2_1_LC_2_4_6  (
            .in0(N__20839),
            .in1(N__20864),
            .in2(N__20892),
            .in3(N__20634),
            .lcout(\spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i ),
            .ltout(\spi_master_inst.sclk_gen_u0.un1_sclk_count_start_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_RNIPPNJ2_LC_2_4_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_RNIPPNJ2_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_RNIPPNJ2_LC_2_4_7 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_start_i_RNIPPNJ2_LC_2_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20619),
            .in3(N__22531),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_i_0_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_0_LC_2_5_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_0_LC_2_5_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_0_LC_2_5_1 .LUT_INIT=16'b0001111101000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_0_LC_2_5_1  (
            .in0(N__21026),
            .in1(N__20736),
            .in2(N__20994),
            .in3(N__21172),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53272),
            .ce(),
            .sr(N__53144));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_1_LC_2_5_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_1_LC_2_5_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_1_LC_2_5_2 .LUT_INIT=16'b0001010011110000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_1_LC_2_5_2  (
            .in0(N__21027),
            .in1(N__20943),
            .in2(N__21416),
            .in3(N__20984),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53272),
            .ce(),
            .sr(N__53144));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_6_LC_2_5_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_6_LC_2_5_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_6_LC_2_5_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_6_LC_2_5_7  (
            .in0(N__25752),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53272),
            .ce(),
            .sr(N__53144));
    defparam sRAM_pointer_read_0_LC_2_11_0.C_ON=1'b1;
    defparam sRAM_pointer_read_0_LC_2_11_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_0_LC_2_11_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_0_LC_2_11_0 (
            .in0(N__33548),
            .in1(N__29750),
            .in2(_gnd_net_),
            .in3(N__20616),
            .lcout(sRAM_pointer_readZ0Z_0),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(sRAM_pointer_read_cry_0),
            .clk(N__47843),
            .ce(N__20701),
            .sr(N__53118));
    defparam sRAM_pointer_read_1_LC_2_11_1.C_ON=1'b1;
    defparam sRAM_pointer_read_1_LC_2_11_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_1_LC_2_11_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_1_LC_2_11_1 (
            .in0(N__33544),
            .in1(N__29675),
            .in2(_gnd_net_),
            .in3(N__20613),
            .lcout(sRAM_pointer_readZ0Z_1),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_0),
            .carryout(sRAM_pointer_read_cry_1),
            .clk(N__47843),
            .ce(N__20701),
            .sr(N__53118));
    defparam sRAM_pointer_read_2_LC_2_11_2.C_ON=1'b1;
    defparam sRAM_pointer_read_2_LC_2_11_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_2_LC_2_11_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_2_LC_2_11_2 (
            .in0(N__33549),
            .in1(N__28067),
            .in2(_gnd_net_),
            .in3(N__20673),
            .lcout(sRAM_pointer_readZ0Z_2),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_1),
            .carryout(sRAM_pointer_read_cry_2),
            .clk(N__47843),
            .ce(N__20701),
            .sr(N__53118));
    defparam sRAM_pointer_read_3_LC_2_11_3.C_ON=1'b1;
    defparam sRAM_pointer_read_3_LC_2_11_3.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_3_LC_2_11_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_3_LC_2_11_3 (
            .in0(N__33545),
            .in1(N__28673),
            .in2(_gnd_net_),
            .in3(N__20670),
            .lcout(sRAM_pointer_readZ0Z_3),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_2),
            .carryout(sRAM_pointer_read_cry_3),
            .clk(N__47843),
            .ce(N__20701),
            .sr(N__53118));
    defparam sRAM_pointer_read_4_LC_2_11_4.C_ON=1'b1;
    defparam sRAM_pointer_read_4_LC_2_11_4.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_4_LC_2_11_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_4_LC_2_11_4 (
            .in0(N__33550),
            .in1(N__28637),
            .in2(_gnd_net_),
            .in3(N__20667),
            .lcout(sRAM_pointer_readZ0Z_4),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_3),
            .carryout(sRAM_pointer_read_cry_4),
            .clk(N__47843),
            .ce(N__20701),
            .sr(N__53118));
    defparam sRAM_pointer_read_5_LC_2_11_5.C_ON=1'b1;
    defparam sRAM_pointer_read_5_LC_2_11_5.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_5_LC_2_11_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_5_LC_2_11_5 (
            .in0(N__33546),
            .in1(N__28592),
            .in2(_gnd_net_),
            .in3(N__20664),
            .lcout(sRAM_pointer_readZ0Z_5),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_4),
            .carryout(sRAM_pointer_read_cry_5),
            .clk(N__47843),
            .ce(N__20701),
            .sr(N__53118));
    defparam sRAM_pointer_read_6_LC_2_11_6.C_ON=1'b1;
    defparam sRAM_pointer_read_6_LC_2_11_6.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_6_LC_2_11_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_6_LC_2_11_6 (
            .in0(N__33551),
            .in1(N__28547),
            .in2(_gnd_net_),
            .in3(N__20661),
            .lcout(sRAM_pointer_readZ0Z_6),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_5),
            .carryout(sRAM_pointer_read_cry_6),
            .clk(N__47843),
            .ce(N__20701),
            .sr(N__53118));
    defparam sRAM_pointer_read_7_LC_2_11_7.C_ON=1'b1;
    defparam sRAM_pointer_read_7_LC_2_11_7.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_7_LC_2_11_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_7_LC_2_11_7 (
            .in0(N__33547),
            .in1(N__28499),
            .in2(_gnd_net_),
            .in3(N__20658),
            .lcout(sRAM_pointer_readZ0Z_7),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_6),
            .carryout(sRAM_pointer_read_cry_7),
            .clk(N__47843),
            .ce(N__20701),
            .sr(N__53118));
    defparam sRAM_pointer_read_8_LC_2_12_0.C_ON=1'b1;
    defparam sRAM_pointer_read_8_LC_2_12_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_8_LC_2_12_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_8_LC_2_12_0 (
            .in0(N__33459),
            .in1(N__28451),
            .in2(_gnd_net_),
            .in3(N__20655),
            .lcout(sRAM_pointer_readZ0Z_8),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(sRAM_pointer_read_cry_8),
            .clk(N__47852),
            .ce(N__20702),
            .sr(N__53105));
    defparam sRAM_pointer_read_9_LC_2_12_1.C_ON=1'b1;
    defparam sRAM_pointer_read_9_LC_2_12_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_9_LC_2_12_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_9_LC_2_12_1 (
            .in0(N__33446),
            .in1(N__28403),
            .in2(_gnd_net_),
            .in3(N__20652),
            .lcout(sRAM_pointer_readZ0Z_9),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_8),
            .carryout(sRAM_pointer_read_cry_9),
            .clk(N__47852),
            .ce(N__20702),
            .sr(N__53105));
    defparam sRAM_pointer_read_10_LC_2_12_2.C_ON=1'b1;
    defparam sRAM_pointer_read_10_LC_2_12_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_10_LC_2_12_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_10_LC_2_12_2 (
            .in0(N__33456),
            .in1(N__29630),
            .in2(_gnd_net_),
            .in3(N__20649),
            .lcout(sRAM_pointer_readZ0Z_10),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_9),
            .carryout(sRAM_pointer_read_cry_10),
            .clk(N__47852),
            .ce(N__20702),
            .sr(N__53105));
    defparam sRAM_pointer_read_11_LC_2_12_3.C_ON=1'b1;
    defparam sRAM_pointer_read_11_LC_2_12_3.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_11_LC_2_12_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_11_LC_2_12_3 (
            .in0(N__33443),
            .in1(N__30392),
            .in2(_gnd_net_),
            .in3(N__20646),
            .lcout(sRAM_pointer_readZ0Z_11),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_10),
            .carryout(sRAM_pointer_read_cry_11),
            .clk(N__47852),
            .ce(N__20702),
            .sr(N__53105));
    defparam sRAM_pointer_read_12_LC_2_12_4.C_ON=1'b1;
    defparam sRAM_pointer_read_12_LC_2_12_4.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_12_LC_2_12_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_12_LC_2_12_4 (
            .in0(N__33457),
            .in1(N__30338),
            .in2(_gnd_net_),
            .in3(N__20724),
            .lcout(sRAM_pointer_readZ0Z_12),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_11),
            .carryout(sRAM_pointer_read_cry_12),
            .clk(N__47852),
            .ce(N__20702),
            .sr(N__53105));
    defparam sRAM_pointer_read_13_LC_2_12_5.C_ON=1'b1;
    defparam sRAM_pointer_read_13_LC_2_12_5.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_13_LC_2_12_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_13_LC_2_12_5 (
            .in0(N__33444),
            .in1(N__30302),
            .in2(_gnd_net_),
            .in3(N__20721),
            .lcout(sRAM_pointer_readZ0Z_13),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_12),
            .carryout(sRAM_pointer_read_cry_13),
            .clk(N__47852),
            .ce(N__20702),
            .sr(N__53105));
    defparam sRAM_pointer_read_14_LC_2_12_6.C_ON=1'b1;
    defparam sRAM_pointer_read_14_LC_2_12_6.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_14_LC_2_12_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_14_LC_2_12_6 (
            .in0(N__33458),
            .in1(N__28289),
            .in2(_gnd_net_),
            .in3(N__20718),
            .lcout(sRAM_pointer_readZ0Z_14),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_13),
            .carryout(sRAM_pointer_read_cry_14),
            .clk(N__47852),
            .ce(N__20702),
            .sr(N__53105));
    defparam sRAM_pointer_read_15_LC_2_12_7.C_ON=1'b1;
    defparam sRAM_pointer_read_15_LC_2_12_7.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_15_LC_2_12_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_15_LC_2_12_7 (
            .in0(N__33445),
            .in1(N__28241),
            .in2(_gnd_net_),
            .in3(N__20715),
            .lcout(sRAM_pointer_readZ0Z_15),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_14),
            .carryout(sRAM_pointer_read_cry_15),
            .clk(N__47852),
            .ce(N__20702),
            .sr(N__53105));
    defparam sRAM_pointer_read_16_LC_2_13_0.C_ON=1'b1;
    defparam sRAM_pointer_read_16_LC_2_13_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_16_LC_2_13_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_16_LC_2_13_0 (
            .in0(N__33503),
            .in1(N__28199),
            .in2(_gnd_net_),
            .in3(N__20712),
            .lcout(sRAM_pointer_readZ0Z_16),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(sRAM_pointer_read_cry_16),
            .clk(N__47853),
            .ce(N__20703),
            .sr(N__53089));
    defparam sRAM_pointer_read_17_LC_2_13_1.C_ON=1'b1;
    defparam sRAM_pointer_read_17_LC_2_13_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_17_LC_2_13_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_17_LC_2_13_1 (
            .in0(N__33484),
            .in1(N__28151),
            .in2(_gnd_net_),
            .in3(N__20709),
            .lcout(sRAM_pointer_readZ0Z_17),
            .ltout(),
            .carryin(sRAM_pointer_read_cry_16),
            .carryout(sRAM_pointer_read_cry_17),
            .clk(N__47853),
            .ce(N__20703),
            .sr(N__53089));
    defparam sRAM_pointer_read_18_LC_2_13_2.C_ON=1'b0;
    defparam sRAM_pointer_read_18_LC_2_13_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_read_18_LC_2_13_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_read_18_LC_2_13_2 (
            .in0(N__33504),
            .in1(N__28109),
            .in2(_gnd_net_),
            .in3(N__20706),
            .lcout(sRAM_pointer_readZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47853),
            .ce(N__20703),
            .sr(N__53089));
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_RNO_0_LC_3_2_4 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_RNO_0_LC_3_2_4 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_RNO_0_LC_3_2_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \spi_master_inst.sclk_gen_u0.div_clk_i_RNO_0_LC_3_2_4  (
            .in0(N__20863),
            .in1(N__20755),
            .in2(N__20844),
            .in3(N__20813),
            .lcout(\spi_master_inst.sclk_gen_u0.div_clk_i2lto7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_0_LC_3_3_0 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_0_LC_3_3_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_0_LC_3_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_0_LC_3_3_0  (
            .in0(_gnd_net_),
            .in1(N__20688),
            .in2(_gnd_net_),
            .in3(N__20895),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_i_s_0 ),
            .ltout(),
            .carryin(bfn_3_3_0_),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_1_LC_3_3_1 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_1_LC_3_3_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_1_LC_3_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_RNO_0_1_LC_3_3_1  (
            .in0(_gnd_net_),
            .in1(N__20888),
            .in2(_gnd_net_),
            .in3(N__20868),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_i_s_1 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_0 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_2_LC_3_3_2 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_2_LC_3_3_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_2_LC_3_3_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_2_LC_3_3_2  (
            .in0(N__20791),
            .in1(N__20865),
            .in2(_gnd_net_),
            .in3(N__20847),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_2 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_1 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2 ),
            .clk(N__53260),
            .ce(),
            .sr(N__53146));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_3_LC_3_3_3 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_3_LC_3_3_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_3_LC_3_3_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_3_LC_3_3_3  (
            .in0(N__20786),
            .in1(N__20840),
            .in2(_gnd_net_),
            .in3(N__20823),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_2 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3 ),
            .clk(N__53260),
            .ce(),
            .sr(N__53146));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_4_LC_3_3_4 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_4_LC_3_3_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_4_LC_3_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_4_LC_3_3_4  (
            .in0(N__20792),
            .in1(N__21086),
            .in2(_gnd_net_),
            .in3(N__20820),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_3 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4 ),
            .clk(N__53260),
            .ce(),
            .sr(N__53146));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_5_LC_3_3_5 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_5_LC_3_3_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_5_LC_3_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_5_LC_3_3_5  (
            .in0(N__20787),
            .in1(N__21110),
            .in2(_gnd_net_),
            .in3(N__20817),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_5 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_4 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5 ),
            .clk(N__53260),
            .ce(),
            .sr(N__53146));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_6_LC_3_3_6 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_6_LC_3_3_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_6_LC_3_3_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_6_LC_3_3_6  (
            .in0(N__20793),
            .in1(N__20814),
            .in2(_gnd_net_),
            .in3(N__20796),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_6 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_5 ),
            .carryout(\spi_master_inst.sclk_gen_u0.sclk_count_i_cry_6 ),
            .clk(N__53260),
            .ce(),
            .sr(N__53146));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_7_LC_3_3_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_7_LC_3_3_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_i_7_LC_3_3_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_i_7_LC_3_3_7  (
            .in0(N__20788),
            .in1(N__20756),
            .in2(_gnd_net_),
            .in3(N__20760),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53260),
            .ce(),
            .sr(N__53146));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_c_LC_3_4_0 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_c_LC_3_4_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_c_LC_3_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_c_LC_3_4_0  (
            .in0(_gnd_net_),
            .in1(N__20735),
            .in2(N__21176),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_4_0_),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_LUT4_0_LC_3_4_1 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_LUT4_0_LC_3_4_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_LUT4_0_LC_3_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_LUT4_0_LC_3_4_1  (
            .in0(_gnd_net_),
            .in1(N__21409),
            .in2(_gnd_net_),
            .in3(N__20937),
            .lcout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_0 ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_LUT4_0_LC_3_4_2 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_LUT4_0_LC_3_4_2 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_LUT4_0_LC_3_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_LUT4_0_LC_3_4_2  (
            .in0(_gnd_net_),
            .in1(N__21701),
            .in2(_gnd_net_),
            .in3(N__20934),
            .lcout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_1 ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_LUT4_0_LC_3_4_3 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_LUT4_0_LC_3_4_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_LUT4_0_LC_3_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_LUT4_0_LC_3_4_3  (
            .in0(_gnd_net_),
            .in1(N__22639),
            .in2(_gnd_net_),
            .in3(N__20931),
            .lcout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_2 ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_4_LC_3_4_4 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_4_LC_3_4_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_4_LC_3_4_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_4_LC_3_4_4  (
            .in0(N__20986),
            .in1(N__20928),
            .in2(_gnd_net_),
            .in3(N__20916),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_3 ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4 ),
            .clk(N__53266),
            .ce(),
            .sr(N__53145));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_0_LC_3_4_5 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_0_LC_3_4_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_0_LC_3_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_0_LC_3_4_5  (
            .in0(_gnd_net_),
            .in1(N__37824),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4 ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_1_LC_3_4_6 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_1_LC_3_4_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_1_LC_3_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_1_LC_3_4_6  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__37907),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_0_THRU_CO ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_2_LC_3_4_7 .C_ON=1'b1;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_2_LC_3_4_7 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_2_LC_3_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_c_THRU_CRY_2_LC_3_4_7  (
            .in0(_gnd_net_),
            .in1(N__37828),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_1_THRU_CO ),
            .carryout(\spi_master_inst.spi_data_path_u1.un1_tx_data_count_neg_sclk_i_cry_4_THRU_CRY_2_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_5_LC_3_5_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_5_LC_3_5_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_5_LC_3_5_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_er_5_LC_3_5_0  (
            .in0(_gnd_net_),
            .in1(N__20909),
            .in2(_gnd_net_),
            .in3(N__20913),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53270),
            .ce(N__20985),
            .sr(N__53143));
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_RNIH6AC_LC_3_6_3 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_RNIH6AC_LC_3_6_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_RNIH6AC_LC_3_6_3 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.o_sclk_RNIH6AC_LC_3_6_3  (
            .in0(N__22492),
            .in1(N__23688),
            .in2(_gnd_net_),
            .in3(N__21059),
            .lcout(\spi_master_inst.o_sclk_RNIH6AC ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_ft_ibuf_RNI4OFN_LC_3_7_4.C_ON=1'b0;
    defparam trig_ft_ibuf_RNI4OFN_LC_3_7_4.SEQ_MODE=4'b0000;
    defparam trig_ft_ibuf_RNI4OFN_LC_3_7_4.LUT_INIT=16'b0000000000010001;
    LogicCell40 trig_ft_ibuf_RNI4OFN_LC_3_7_4 (
            .in0(N__23892),
            .in1(N__23964),
            .in2(_gnd_net_),
            .in3(N__24040),
            .lcout(un3_trig_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_3_8_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_3_8_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_3_8_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_3_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_ft_ibuf_RNI4OFN_0_LC_3_10_3.C_ON=1'b0;
    defparam trig_ft_ibuf_RNI4OFN_0_LC_3_10_3.SEQ_MODE=4'b0000;
    defparam trig_ft_ibuf_RNI4OFN_0_LC_3_10_3.LUT_INIT=16'b0000000000010001;
    LogicCell40 trig_ft_ibuf_RNI4OFN_0_LC_3_10_3 (
            .in0(N__23931),
            .in1(N__23907),
            .in2(_gnd_net_),
            .in3(N__24024),
            .lcout(un3_trig_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI70MD9_0_LC_5_3_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI70MD9_0_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI70MD9_0_LC_5_3_4 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI70MD9_0_LC_5_3_4  (
            .in0(N__21297),
            .in1(N__21429),
            .in2(N__21387),
            .in3(N__21180),
            .lcout(DAC_mosi_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_LC_5_4_1 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_LC_5_4_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.div_clk_i_LC_5_4_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.div_clk_i_LC_5_4_1  (
            .in0(N__21129),
            .in1(N__21117),
            .in2(_gnd_net_),
            .in3(N__21093),
            .lcout(\spi_master_inst.sclk_gen_u0.div_clk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53255),
            .ce(),
            .sr(N__53142));
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_LC_5_4_3 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_LC_5_4_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.o_sclk_LC_5_4_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.o_sclk_LC_5_4_3  (
            .in0(_gnd_net_),
            .in1(N__22483),
            .in2(_gnd_net_),
            .in3(N__23694),
            .lcout(DAC_sclk_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53255),
            .ce(),
            .sr(N__53142));
    defparam \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_i_LC_5_4_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_i_LC_5_4_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_i_LC_5_4_4 .LUT_INIT=16'b1111100011011000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_i_LC_5_4_4  (
            .in0(N__20995),
            .in1(N__21028),
            .in2(N__27026),
            .in3(N__21296),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_done_neg_sclk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53255),
            .ce(),
            .sr(N__53142));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_2_LC_5_4_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_2_LC_5_4_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_2_LC_5_4_6 .LUT_INIT=16'b0001110001001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_2_LC_5_4_6  (
            .in0(N__21030),
            .in1(N__21692),
            .in2(N__21000),
            .in3(N__21039),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53255),
            .ce(),
            .sr(N__53142));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_3_LC_5_4_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_3_LC_5_4_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_3_LC_5_4_7 .LUT_INIT=16'b0011010001110000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_3_LC_5_4_7  (
            .in0(N__21029),
            .in1(N__20999),
            .in2(N__22636),
            .in3(N__20952),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53255),
            .ce(),
            .sr(N__53142));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_0_LC_5_5_0 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_0_LC_5_5_0 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_0_LC_5_5_0 .LUT_INIT=16'b1011101111101110;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_0_LC_5_5_0  (
            .in0(N__21460),
            .in1(N__21570),
            .in2(_gnd_net_),
            .in3(N__21255),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_5_0_),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_0 ),
            .clk(N__53261),
            .ce(),
            .sr(N__53141));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_1_LC_5_5_1 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_1_LC_5_5_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_1_LC_5_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_1_LC_5_5_1  (
            .in0(N__21455),
            .in1(N__21624),
            .in2(_gnd_net_),
            .in3(N__21252),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_1 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_0 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_1 ),
            .clk(N__53261),
            .ce(),
            .sr(N__53141));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_2_LC_5_5_2 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_2_LC_5_5_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_2_LC_5_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_2_LC_5_5_2  (
            .in0(N__21461),
            .in1(N__21605),
            .in2(_gnd_net_),
            .in3(N__21249),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_2 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_1 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_2 ),
            .clk(N__53261),
            .ce(),
            .sr(N__53141));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_3_LC_5_5_3 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_3_LC_5_5_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_3_LC_5_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_3_LC_5_5_3  (
            .in0(N__21456),
            .in1(N__21642),
            .in2(_gnd_net_),
            .in3(N__21246),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_2 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_3 ),
            .clk(N__53261),
            .ce(),
            .sr(N__53141));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_4_LC_5_5_4 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_4_LC_5_5_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_4_LC_5_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_4_LC_5_5_4  (
            .in0(N__21462),
            .in1(N__21192),
            .in2(_gnd_net_),
            .in3(N__21243),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_3 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_4 ),
            .clk(N__53261),
            .ce(),
            .sr(N__53141));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_5_LC_5_5_5 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_5_LC_5_5_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_5_LC_5_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_5_LC_5_5_5  (
            .in0(N__21457),
            .in1(N__21219),
            .in2(_gnd_net_),
            .in3(N__21240),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_5 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_4 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_5 ),
            .clk(N__53261),
            .ce(),
            .sr(N__53141));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_6_LC_5_5_6 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_6_LC_5_5_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_6_LC_5_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_6_LC_5_5_6  (
            .in0(N__21458),
            .in1(N__21231),
            .in2(_gnd_net_),
            .in3(N__21237),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_6 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_5 ),
            .carryout(\spi_master_inst.sclk_gen_u0.delay_count_i_cry_6 ),
            .clk(N__53261),
            .ce(),
            .sr(N__53141));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_7_LC_5_5_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_7_LC_5_5_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_7_LC_5_5_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_7_LC_5_5_7  (
            .in0(N__21206),
            .in1(N__21459),
            .in2(_gnd_net_),
            .in3(N__21234),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53261),
            .ce(),
            .sr(N__53141));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIQU1N1_7_LC_5_6_0 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIQU1N1_7_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIQU1N1_7_LC_5_6_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_RNIQU1N1_7_LC_5_6_0  (
            .in0(N__21230),
            .in1(N__21218),
            .in2(N__21207),
            .in3(N__21191),
            .lcout(\spi_master_inst.sclk_gen_u0.N_1666 ),
            .ltout(\spi_master_inst.sclk_gen_u0.N_1666_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_0_LC_5_6_1 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_0_LC_5_6_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_0_LC_5_6_1 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_0_LC_5_6_1  (
            .in0(N__21321),
            .in1(N__21315),
            .in2(N__21324),
            .in3(N__21471),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53267),
            .ce(),
            .sr(N__53136));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIAE1N1_0_LC_5_6_2 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIAE1N1_0_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNIAE1N1_0_LC_5_6_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_RNIAE1N1_0_LC_5_6_2  (
            .in0(N__21569),
            .in1(N__21623),
            .in2(N__21606),
            .in3(N__21641),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4 ),
            .ltout(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0IPL3_0_LC_5_6_3 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0IPL3_0_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0IPL3_0_LC_5_6_3 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0IPL3_0_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(N__21314),
            .in2(N__21306),
            .in3(N__21585),
            .lcout(\spi_master_inst.sclk_gen_u0.N_48 ),
            .ltout(\spi_master_inst.sclk_gen_u0.N_48_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_4_LC_5_6_4 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_4_LC_5_6_4 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_4_LC_5_6_4 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_4_LC_5_6_4  (
            .in0(N__23727),
            .in1(_gnd_net_),
            .in2(N__21303),
            .in3(N__27003),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53267),
            .ce(),
            .sr(N__53136));
    defparam \spi_master_inst.sclk_gen_u0.o_ss_start_LC_5_6_5 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.o_ss_start_LC_5_6_5 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.sclk_gen_u0.o_ss_start_LC_5_6_5 .LUT_INIT=16'b1111111101110100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.o_ss_start_LC_5_6_5  (
            .in0(N__27002),
            .in1(N__23726),
            .in2(N__21298),
            .in3(N__21470),
            .lcout(\spi_master_inst.ss_start_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53267),
            .ce(),
            .sr(N__53136));
    defparam trig_ft_ibuf_RNI4OFN_2_LC_5_7_0.C_ON=1'b0;
    defparam trig_ft_ibuf_RNI4OFN_2_LC_5_7_0.SEQ_MODE=4'b0000;
    defparam trig_ft_ibuf_RNI4OFN_2_LC_5_7_0.LUT_INIT=16'b0000000000010001;
    LogicCell40 trig_ft_ibuf_RNI4OFN_2_LC_5_7_0 (
            .in0(N__23901),
            .in1(N__23965),
            .in2(_gnd_net_),
            .in3(N__24041),
            .lcout(un3_trig_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_ft_ibuf_RNI4OFN_3_LC_5_7_5.C_ON=1'b0;
    defparam trig_ft_ibuf_RNI4OFN_3_LC_5_7_5.SEQ_MODE=4'b0000;
    defparam trig_ft_ibuf_RNI4OFN_3_LC_5_7_5.LUT_INIT=16'b0000000000000101;
    LogicCell40 trig_ft_ibuf_RNI4OFN_3_LC_5_7_5 (
            .in0(N__23966),
            .in1(_gnd_net_),
            .in2(N__24056),
            .in3(N__23902),
            .lcout(un3_trig_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sSingleCont_LC_5_8_7.C_ON=1'b0;
    defparam sSingleCont_LC_5_8_7.SEQ_MODE=4'b1010;
    defparam sSingleCont_LC_5_8_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 sSingleCont_LC_5_8_7 (
            .in0(_gnd_net_),
            .in1(N__22215),
            .in2(_gnd_net_),
            .in3(N__21978),
            .lcout(LED_MODE_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53273),
            .ce(),
            .sr(N__53119));
    defparam sSPI_MSB0LSB1_LC_5_9_7.C_ON=1'b0;
    defparam sSPI_MSB0LSB1_LC_5_9_7.SEQ_MODE=4'b1010;
    defparam sSPI_MSB0LSB1_LC_5_9_7.LUT_INIT=16'b1101001001011010;
    LogicCell40 sSPI_MSB0LSB1_LC_5_9_7 (
            .in0(N__27911),
            .in1(N__32215),
            .in2(N__27956),
            .in3(N__31977),
            .lcout(sSPI_MSB0LSBZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47842),
            .ce(),
            .sr(N__53106));
    defparam un4_spoff_cry_0_c_inv_LC_5_10_0.C_ON=1'b1;
    defparam un4_spoff_cry_0_c_inv_LC_5_10_0.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_0_c_inv_LC_5_10_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_spoff_cry_0_c_inv_LC_5_10_0 (
            .in0(_gnd_net_),
            .in1(N__21378),
            .in2(N__34245),
            .in3(N__21717),
            .lcout(sEEPonPoff_i_0),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(un4_spoff_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_1_c_inv_LC_5_10_1.C_ON=1'b1;
    defparam un4_spoff_cry_1_c_inv_LC_5_10_1.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_1_c_inv_LC_5_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_spoff_cry_1_c_inv_LC_5_10_1 (
            .in0(_gnd_net_),
            .in1(N__21372),
            .in2(N__35064),
            .in3(N__21783),
            .lcout(sEEPonPoff_i_1),
            .ltout(),
            .carryin(un4_spoff_cry_0),
            .carryout(un4_spoff_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_2_c_inv_LC_5_10_2.C_ON=1'b1;
    defparam un4_spoff_cry_2_c_inv_LC_5_10_2.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_2_c_inv_LC_5_10_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_spoff_cry_2_c_inv_LC_5_10_2 (
            .in0(N__21777),
            .in1(N__21366),
            .in2(N__34968),
            .in3(_gnd_net_),
            .lcout(sEEPonPoff_i_2),
            .ltout(),
            .carryin(un4_spoff_cry_1),
            .carryout(un4_spoff_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_3_c_inv_LC_5_10_3.C_ON=1'b1;
    defparam un4_spoff_cry_3_c_inv_LC_5_10_3.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_3_c_inv_LC_5_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_spoff_cry_3_c_inv_LC_5_10_3 (
            .in0(_gnd_net_),
            .in1(N__34857),
            .in2(N__21360),
            .in3(N__21771),
            .lcout(sEEPonPoff_i_3),
            .ltout(),
            .carryin(un4_spoff_cry_2),
            .carryout(un4_spoff_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_4_c_inv_LC_5_10_4.C_ON=1'b1;
    defparam un4_spoff_cry_4_c_inv_LC_5_10_4.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_4_c_inv_LC_5_10_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_spoff_cry_4_c_inv_LC_5_10_4 (
            .in0(_gnd_net_),
            .in1(N__21351),
            .in2(N__36883),
            .in3(N__21765),
            .lcout(sEEPonPoff_i_4),
            .ltout(),
            .carryin(un4_spoff_cry_3),
            .carryout(un4_spoff_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_5_c_inv_LC_5_10_5.C_ON=1'b1;
    defparam un4_spoff_cry_5_c_inv_LC_5_10_5.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_5_c_inv_LC_5_10_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_spoff_cry_5_c_inv_LC_5_10_5 (
            .in0(_gnd_net_),
            .in1(N__34728),
            .in2(N__21345),
            .in3(N__21759),
            .lcout(sEEPonPoff_i_5),
            .ltout(),
            .carryin(un4_spoff_cry_4),
            .carryout(un4_spoff_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_6_c_inv_LC_5_10_6.C_ON=1'b1;
    defparam un4_spoff_cry_6_c_inv_LC_5_10_6.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_6_c_inv_LC_5_10_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_spoff_cry_6_c_inv_LC_5_10_6 (
            .in0(N__21753),
            .in1(N__21336),
            .in2(N__34620),
            .in3(_gnd_net_),
            .lcout(sEEPonPoff_i_6),
            .ltout(),
            .carryin(un4_spoff_cry_5),
            .carryout(un4_spoff_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_7_c_inv_LC_5_10_7.C_ON=1'b1;
    defparam un4_spoff_cry_7_c_inv_LC_5_10_7.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_7_c_inv_LC_5_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_spoff_cry_7_c_inv_LC_5_10_7 (
            .in0(_gnd_net_),
            .in1(N__21330),
            .in2(N__34494),
            .in3(N__21747),
            .lcout(sEEPonPoff_i_7),
            .ltout(),
            .carryin(un4_spoff_cry_6),
            .carryout(un4_spoff_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_8_c_LC_5_11_0.C_ON=1'b1;
    defparam un4_spoff_cry_8_c_LC_5_11_0.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_8_c_LC_5_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_8_c_LC_5_11_0 (
            .in0(_gnd_net_),
            .in1(N__37841),
            .in2(N__35889),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(un4_spoff_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_9_c_LC_5_11_1.C_ON=1'b1;
    defparam un4_spoff_cry_9_c_LC_5_11_1.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_9_c_LC_5_11_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_9_c_LC_5_11_1 (
            .in0(_gnd_net_),
            .in1(N__35763),
            .in2(N__37911),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_8),
            .carryout(un4_spoff_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_10_c_LC_5_11_2.C_ON=1'b1;
    defparam un4_spoff_cry_10_c_LC_5_11_2.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_10_c_LC_5_11_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_10_c_LC_5_11_2 (
            .in0(_gnd_net_),
            .in1(N__37829),
            .in2(N__35654),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_9),
            .carryout(un4_spoff_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_11_c_LC_5_11_3.C_ON=1'b1;
    defparam un4_spoff_cry_11_c_LC_5_11_3.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_11_c_LC_5_11_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_11_c_LC_5_11_3 (
            .in0(_gnd_net_),
            .in1(N__35541),
            .in2(N__37908),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_10),
            .carryout(un4_spoff_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_12_c_LC_5_11_4.C_ON=1'b1;
    defparam un4_spoff_cry_12_c_LC_5_11_4.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_12_c_LC_5_11_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_12_c_LC_5_11_4 (
            .in0(_gnd_net_),
            .in1(N__37833),
            .in2(N__35418),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_11),
            .carryout(un4_spoff_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_13_c_LC_5_11_5.C_ON=1'b1;
    defparam un4_spoff_cry_13_c_LC_5_11_5.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_13_c_LC_5_11_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_13_c_LC_5_11_5 (
            .in0(_gnd_net_),
            .in1(N__35311),
            .in2(N__37909),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_12),
            .carryout(un4_spoff_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_14_c_LC_5_11_6.C_ON=1'b1;
    defparam un4_spoff_cry_14_c_LC_5_11_6.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_14_c_LC_5_11_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_14_c_LC_5_11_6 (
            .in0(_gnd_net_),
            .in1(N__37837),
            .in2(N__35208),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_13),
            .carryout(un4_spoff_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_15_c_LC_5_11_7.C_ON=1'b1;
    defparam un4_spoff_cry_15_c_LC_5_11_7.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_15_c_LC_5_11_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_15_c_LC_5_11_7 (
            .in0(_gnd_net_),
            .in1(N__36659),
            .in2(N__37910),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_14),
            .carryout(un4_spoff_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_16_c_LC_5_12_0.C_ON=1'b1;
    defparam un4_spoff_cry_16_c_LC_5_12_0.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_16_c_LC_5_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_16_c_LC_5_12_0 (
            .in0(_gnd_net_),
            .in1(N__37865),
            .in2(N__36546),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(un4_spoff_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_17_c_LC_5_12_1.C_ON=1'b1;
    defparam un4_spoff_cry_17_c_LC_5_12_1.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_17_c_LC_5_12_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_17_c_LC_5_12_1 (
            .in0(_gnd_net_),
            .in1(N__36444),
            .in2(N__37929),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_16),
            .carryout(un4_spoff_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_18_c_LC_5_12_2.C_ON=1'b1;
    defparam un4_spoff_cry_18_c_LC_5_12_2.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_18_c_LC_5_12_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_18_c_LC_5_12_2 (
            .in0(_gnd_net_),
            .in1(N__37869),
            .in2(N__36346),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_17),
            .carryout(un4_spoff_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_19_c_LC_5_12_3.C_ON=1'b1;
    defparam un4_spoff_cry_19_c_LC_5_12_3.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_19_c_LC_5_12_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_19_c_LC_5_12_3 (
            .in0(_gnd_net_),
            .in1(N__36254),
            .in2(N__37930),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_18),
            .carryout(un4_spoff_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_20_c_LC_5_12_4.C_ON=1'b1;
    defparam un4_spoff_cry_20_c_LC_5_12_4.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_20_c_LC_5_12_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_20_c_LC_5_12_4 (
            .in0(_gnd_net_),
            .in1(N__37873),
            .in2(N__36169),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_19),
            .carryout(un4_spoff_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIR3KA_20_LC_5_12_5.C_ON=1'b1;
    defparam sCounter_RNIR3KA_20_LC_5_12_5.SEQ_MODE=4'b0000;
    defparam sCounter_RNIR3KA_20_LC_5_12_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 sCounter_RNIR3KA_20_LC_5_12_5 (
            .in0(_gnd_net_),
            .in1(N__36072),
            .in2(N__37928),
            .in3(N__36158),
            .lcout(un1_reset_rpi_inv_2_i_o3_8),
            .ltout(),
            .carryin(un4_spoff_cry_20),
            .carryout(un4_spoff_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_22_c_LC_5_12_6.C_ON=1'b1;
    defparam un4_spoff_cry_22_c_LC_5_12_6.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_22_c_LC_5_12_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_22_c_LC_5_12_6 (
            .in0(_gnd_net_),
            .in1(N__37874),
            .in2(N__36000),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_21),
            .carryout(un4_spoff_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_23_c_LC_5_12_7.C_ON=1'b1;
    defparam un4_spoff_cry_23_c_LC_5_12_7.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_23_c_LC_5_12_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_spoff_cry_23_c_LC_5_12_7 (
            .in0(_gnd_net_),
            .in1(N__37088),
            .in2(N__37931),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_spoff_cry_22),
            .carryout(un4_spoff_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_spoff_cry_23_THRU_LUT4_0_LC_5_13_0.C_ON=1'b0;
    defparam un4_spoff_cry_23_THRU_LUT4_0_LC_5_13_0.SEQ_MODE=4'b0000;
    defparam un4_spoff_cry_23_THRU_LUT4_0_LC_5_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un4_spoff_cry_23_THRU_LUT4_0_LC_5_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21432),
            .lcout(un4_spoff_cry_23_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIUNHB4_1_LC_6_3_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIUNHB4_1_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIUNHB4_1_LC_6_3_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIUNHB4_1_LC_6_3_0  (
            .in0(N__21486),
            .in1(N__21477),
            .in2(_gnd_net_),
            .in3(N__21423),
            .lcout(\spi_master_inst.spi_data_path_u1.N_1423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI60IB4_1_LC_6_3_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI60IB4_1_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI60IB4_1_LC_6_3_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI60IB4_1_LC_6_3_2  (
            .in0(N__21651),
            .in1(N__21507),
            .in2(_gnd_net_),
            .in3(N__21422),
            .lcout(\spi_master_inst.spi_data_path_u1.N_1416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI73G42_2_LC_6_4_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI73G42_2_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI73G42_2_LC_6_4_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI73G42_2_LC_6_4_0  (
            .in0(N__21694),
            .in1(N__21990),
            .in2(_gnd_net_),
            .in3(N__21984),
            .lcout(\spi_master_inst.spi_data_path_u1.N_1415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4Q_14_LC_6_4_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4Q_14_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4Q_14_LC_6_4_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4Q_14_LC_6_4_1  (
            .in0(N__22458),
            .in1(N__21501),
            .in2(_gnd_net_),
            .in3(N__22628),
            .lcout(),
            .ltout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIOJ4QZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIICLT1_2_LC_6_4_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIICLT1_2_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIICLT1_2_LC_6_4_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIICLT1_2_LC_6_4_2  (
            .in0(N__21695),
            .in1(_gnd_net_),
            .in2(N__21489),
            .in3(N__22398),
            .lcout(\spi_master_inst.spi_data_path_u1.N_1419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01_0_LC_6_4_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01_0_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01_0_LC_6_4_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01_0_LC_6_4_6  (
            .in0(N__22627),
            .in1(N__22437),
            .in2(_gnd_net_),
            .in3(N__22446),
            .lcout(),
            .ltout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI52V01Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI3VF42_2_LC_6_4_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI3VF42_2_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI3VF42_2_LC_6_4_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNI3VF42_2_LC_6_4_7  (
            .in0(N__22569),
            .in1(_gnd_net_),
            .in2(N__21480),
            .in3(N__21693),
            .lcout(\spi_master_inst.spi_data_path_u1.N_1422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI1JPL3_1_LC_6_5_1 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI1JPL3_1_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI1JPL3_1_LC_6_5_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI1JPL3_1_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(N__21524),
            .in2(_gnd_net_),
            .in3(N__21948),
            .lcout(\spi_master_inst.sclk_gen_u0.N_1520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4Q_11_LC_6_5_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4Q_11_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4Q_11_LC_6_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4Q_11_LC_6_5_3  (
            .in0(N__23772),
            .in1(N__23580),
            .in2(_gnd_net_),
            .in3(N__22617),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIID4QZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNI6TQC_LC_6_5_5 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNI6TQC_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNI6TQC_LC_6_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNI6TQC_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21536),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_start_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4Q_15_LC_6_5_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4Q_15_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4Q_15_LC_6_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4Q_15_LC_6_5_6  (
            .in0(N__22618),
            .in1(N__22422),
            .in2(_gnd_net_),
            .in3(N__23781),
            .lcout(),
            .ltout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIQL4QZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIMGLT1_2_LC_6_5_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIMGLT1_2_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIMGLT1_2_LC_6_5_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_data_count_neg_sclk_i_RNIMGLT1_2_LC_6_5_7  (
            .in0(N__21711),
            .in1(_gnd_net_),
            .in2(N__21705),
            .in3(N__21696),
            .lcout(\spi_master_inst.spi_data_path_u1.N_1412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI6OGR_1_LC_6_6_0 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI6OGR_1_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI6OGR_1_LC_6_6_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_RNI6OGR_1_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__21640),
            .in2(_gnd_net_),
            .in3(N__21622),
            .lcout(),
            .ltout(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_o2_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4D3E3_0_LC_6_6_1 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4D3E3_0_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4D3E3_0_LC_6_6_1 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_i_RNI4D3E3_0_LC_6_6_1  (
            .in0(N__21601),
            .in1(N__21584),
            .in2(N__21573),
            .in3(N__21568),
            .lcout(\spi_master_inst.sclk_gen_u0.N_1515 ),
            .ltout(\spi_master_inst.sclk_gen_u0.N_1515_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0RFT3_1_LC_6_6_2 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0RFT3_1_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0RFT3_1_LC_6_6_2 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI0RFT3_1_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__21964),
            .in2(N__21552),
            .in3(N__21520),
            .lcout(\spi_master_inst.sclk_gen_u0.N_36 ),
            .ltout(\spi_master_inst.sclk_gen_u0.N_36_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNO_0_LC_6_6_3 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNO_0_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNO_0_LC_6_6_3 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_start_i_RNO_0_LC_6_6_3  (
            .in0(N__23717),
            .in1(N__27000),
            .in2(N__21549),
            .in3(N__21546),
            .lcout(),
            .ltout(\spi_master_inst.sclk_gen_u0.N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_LC_6_6_4 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_LC_6_6_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_count_start_i_LC_6_6_4 .LUT_INIT=16'b0000111110001101;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_count_start_i_LC_6_6_4  (
            .in0(N__23692),
            .in1(N__21537),
            .in2(N__21540),
            .in3(N__23756),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_count_start_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53256),
            .ce(),
            .sr(N__53120));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_1_LC_6_6_5 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_1_LC_6_6_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_1_LC_6_6_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_1_LC_6_6_5  (
            .in0(N__23757),
            .in1(N__23693),
            .in2(N__21525),
            .in3(N__21950),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53256),
            .ce(),
            .sr(N__53120));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_3_LC_6_6_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_3_LC_6_6_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_3_LC_6_6_7 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_3_LC_6_6_7  (
            .in0(N__21965),
            .in1(N__27001),
            .in2(N__23728),
            .in3(N__21951),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53256),
            .ce(),
            .sr(N__53120));
    defparam sTrigCounter_RNO_2_0_LC_6_7_3.C_ON=1'b0;
    defparam sTrigCounter_RNO_2_0_LC_6_7_3.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_2_0_LC_6_7_3.LUT_INIT=16'b1010100011111100;
    LogicCell40 sTrigCounter_RNO_2_0_LC_6_7_3 (
            .in0(N__24927),
            .in1(N__24488),
            .in2(N__22091),
            .in3(N__29094),
            .lcout(g1_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_ft_ibuf_RNI4OFN_5_LC_6_7_7.C_ON=1'b0;
    defparam trig_ft_ibuf_RNI4OFN_5_LC_6_7_7.SEQ_MODE=4'b0000;
    defparam trig_ft_ibuf_RNI4OFN_5_LC_6_7_7.LUT_INIT=16'b0000000000010001;
    LogicCell40 trig_ft_ibuf_RNI4OFN_5_LC_6_7_7 (
            .in0(N__24057),
            .in1(N__23900),
            .in2(_gnd_net_),
            .in3(N__23970),
            .lcout(un3_trig_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPon_0_LC_6_8_0.C_ON=1'b0;
    defparam sEEPon_0_LC_6_8_0.SEQ_MODE=4'b1010;
    defparam sEEPon_0_LC_6_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_0_LC_6_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51258),
            .lcout(sEEPonZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47836),
            .ce(N__30896),
            .sr(N__53091));
    defparam sEEPon_1_LC_6_8_1.C_ON=1'b0;
    defparam sEEPon_1_LC_6_8_1.SEQ_MODE=4'b1010;
    defparam sEEPon_1_LC_6_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_1_LC_6_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50675),
            .lcout(sEEPonZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47836),
            .ce(N__30896),
            .sr(N__53091));
    defparam sEEPon_7_LC_6_8_2.C_ON=1'b0;
    defparam sEEPon_7_LC_6_8_2.SEQ_MODE=4'b1010;
    defparam sEEPon_7_LC_6_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_7_LC_6_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48798),
            .lcout(sEEPonZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47836),
            .ce(N__30896),
            .sr(N__53091));
    defparam sEEPon_3_LC_6_8_3.C_ON=1'b0;
    defparam sEEPon_3_LC_6_8_3.SEQ_MODE=4'b1010;
    defparam sEEPon_3_LC_6_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_3_LC_6_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49821),
            .lcout(sEEPonZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47836),
            .ce(N__30896),
            .sr(N__53091));
    defparam sEEPon_4_LC_6_8_4.C_ON=1'b0;
    defparam sEEPon_4_LC_6_8_4.SEQ_MODE=4'b1011;
    defparam sEEPon_4_LC_6_8_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPon_4_LC_6_8_4 (
            .in0(N__49345),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPonZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47836),
            .ce(N__30896),
            .sr(N__53091));
    defparam sEEPon_6_LC_6_8_6.C_ON=1'b0;
    defparam sEEPon_6_LC_6_8_6.SEQ_MODE=4'b1010;
    defparam sEEPon_6_LC_6_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_6_LC_6_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48306),
            .lcout(sEEPonZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47836),
            .ce(N__30896),
            .sr(N__53091));
    defparam sEEPon_5_LC_6_9_3.C_ON=1'b0;
    defparam sEEPon_5_LC_6_9_3.SEQ_MODE=4'b1010;
    defparam sEEPon_5_LC_6_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_5_LC_6_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47118),
            .lcout(sEEPonZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47827),
            .ce(N__30900),
            .sr(N__53080));
    defparam sEEPon_2_LC_6_9_5.C_ON=1'b0;
    defparam sEEPon_2_LC_6_9_5.SEQ_MODE=4'b1011;
    defparam sEEPon_2_LC_6_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPon_2_LC_6_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50283),
            .lcout(sEEPonZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47827),
            .ce(N__30900),
            .sr(N__53080));
    defparam sEEPonPoff_0_LC_6_10_0.C_ON=1'b0;
    defparam sEEPonPoff_0_LC_6_10_0.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_0_LC_6_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_0_LC_6_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51232),
            .lcout(sEEPonPoffZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47819),
            .ce(N__30810),
            .sr(N__53068));
    defparam sEEPonPoff_1_LC_6_10_1.C_ON=1'b0;
    defparam sEEPonPoff_1_LC_6_10_1.SEQ_MODE=4'b1011;
    defparam sEEPonPoff_1_LC_6_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_1_LC_6_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50676),
            .lcout(sEEPonPoffZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47819),
            .ce(N__30810),
            .sr(N__53068));
    defparam sEEPonPoff_2_LC_6_10_2.C_ON=1'b0;
    defparam sEEPonPoff_2_LC_6_10_2.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_2_LC_6_10_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPonPoff_2_LC_6_10_2 (
            .in0(N__50285),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPonPoffZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47819),
            .ce(N__30810),
            .sr(N__53068));
    defparam sEEPonPoff_3_LC_6_10_3.C_ON=1'b0;
    defparam sEEPonPoff_3_LC_6_10_3.SEQ_MODE=4'b1011;
    defparam sEEPonPoff_3_LC_6_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_3_LC_6_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49823),
            .lcout(sEEPonPoffZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47819),
            .ce(N__30810),
            .sr(N__53068));
    defparam sEEPonPoff_4_LC_6_10_4.C_ON=1'b0;
    defparam sEEPonPoff_4_LC_6_10_4.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_4_LC_6_10_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPonPoff_4_LC_6_10_4 (
            .in0(N__49347),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPonPoffZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47819),
            .ce(N__30810),
            .sr(N__53068));
    defparam sEEPonPoff_5_LC_6_10_5.C_ON=1'b0;
    defparam sEEPonPoff_5_LC_6_10_5.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_5_LC_6_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_5_LC_6_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47072),
            .lcout(sEEPonPoffZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47819),
            .ce(N__30810),
            .sr(N__53068));
    defparam sEEPonPoff_6_LC_6_10_6.C_ON=1'b0;
    defparam sEEPonPoff_6_LC_6_10_6.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_6_LC_6_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPonPoff_6_LC_6_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48336),
            .lcout(sEEPonPoffZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47819),
            .ce(N__30810),
            .sr(N__53068));
    defparam sEEPonPoff_7_LC_6_10_7.C_ON=1'b0;
    defparam sEEPonPoff_7_LC_6_10_7.SEQ_MODE=4'b1010;
    defparam sEEPonPoff_7_LC_6_10_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPonPoff_7_LC_6_10_7 (
            .in0(N__48593),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPonPoffZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47819),
            .ce(N__30810),
            .sr(N__53068));
    defparam un7_spon_cry_0_c_inv_LC_6_11_0.C_ON=1'b1;
    defparam un7_spon_cry_0_c_inv_LC_6_11_0.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_0_c_inv_LC_6_11_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 un7_spon_cry_0_c_inv_LC_6_11_0 (
            .in0(N__21741),
            .in1(N__21732),
            .in2(N__34243),
            .in3(_gnd_net_),
            .lcout(sEEPon_i_0),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(un7_spon_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_1_c_inv_LC_6_11_1.C_ON=1'b1;
    defparam un7_spon_cry_1_c_inv_LC_6_11_1.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_1_c_inv_LC_6_11_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un7_spon_cry_1_c_inv_LC_6_11_1 (
            .in0(_gnd_net_),
            .in1(N__21885),
            .in2(N__35063),
            .in3(N__21726),
            .lcout(sEEPon_i_1),
            .ltout(),
            .carryin(un7_spon_cry_0),
            .carryout(un7_spon_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_2_c_inv_LC_6_11_2.C_ON=1'b1;
    defparam un7_spon_cry_2_c_inv_LC_6_11_2.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_2_c_inv_LC_6_11_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 un7_spon_cry_2_c_inv_LC_6_11_2 (
            .in0(N__21879),
            .in1(N__21870),
            .in2(N__34964),
            .in3(_gnd_net_),
            .lcout(sEEPon_i_2),
            .ltout(),
            .carryin(un7_spon_cry_1),
            .carryout(un7_spon_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_3_c_inv_LC_6_11_3.C_ON=1'b1;
    defparam un7_spon_cry_3_c_inv_LC_6_11_3.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_3_c_inv_LC_6_11_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un7_spon_cry_3_c_inv_LC_6_11_3 (
            .in0(_gnd_net_),
            .in1(N__34851),
            .in2(N__21855),
            .in3(N__21864),
            .lcout(sEEPon_i_3),
            .ltout(),
            .carryin(un7_spon_cry_2),
            .carryout(un7_spon_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_4_c_inv_LC_6_11_4.C_ON=1'b1;
    defparam un7_spon_cry_4_c_inv_LC_6_11_4.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_4_c_inv_LC_6_11_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un7_spon_cry_4_c_inv_LC_6_11_4 (
            .in0(_gnd_net_),
            .in1(N__21837),
            .in2(N__36882),
            .in3(N__21846),
            .lcout(sEEPon_i_4),
            .ltout(),
            .carryin(un7_spon_cry_3),
            .carryout(un7_spon_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_5_c_inv_LC_6_11_5.C_ON=1'b1;
    defparam un7_spon_cry_5_c_inv_LC_6_11_5.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_5_c_inv_LC_6_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un7_spon_cry_5_c_inv_LC_6_11_5 (
            .in0(_gnd_net_),
            .in1(N__21822),
            .in2(N__34727),
            .in3(N__21831),
            .lcout(sEEPon_i_5),
            .ltout(),
            .carryin(un7_spon_cry_4),
            .carryout(un7_spon_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_6_c_inv_LC_6_11_6.C_ON=1'b1;
    defparam un7_spon_cry_6_c_inv_LC_6_11_6.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_6_c_inv_LC_6_11_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un7_spon_cry_6_c_inv_LC_6_11_6 (
            .in0(_gnd_net_),
            .in1(N__21804),
            .in2(N__34619),
            .in3(N__21816),
            .lcout(sEEPon_i_6),
            .ltout(),
            .carryin(un7_spon_cry_5),
            .carryout(un7_spon_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_7_c_inv_LC_6_11_7.C_ON=1'b1;
    defparam un7_spon_cry_7_c_inv_LC_6_11_7.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_7_c_inv_LC_6_11_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un7_spon_cry_7_c_inv_LC_6_11_7 (
            .in0(N__21798),
            .in1(N__21789),
            .in2(N__34489),
            .in3(_gnd_net_),
            .lcout(sEEPon_i_7),
            .ltout(),
            .carryin(un7_spon_cry_6),
            .carryout(un7_spon_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_8_c_LC_6_12_0.C_ON=1'b1;
    defparam un7_spon_cry_8_c_LC_6_12_0.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_8_c_LC_6_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_8_c_LC_6_12_0 (
            .in0(_gnd_net_),
            .in1(N__37944),
            .in2(N__35881),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_12_0_),
            .carryout(un7_spon_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_9_c_LC_6_12_1.C_ON=1'b1;
    defparam un7_spon_cry_9_c_LC_6_12_1.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_9_c_LC_6_12_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_9_c_LC_6_12_1 (
            .in0(_gnd_net_),
            .in1(N__35767),
            .in2(N__37971),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_8),
            .carryout(un7_spon_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_10_c_LC_6_12_2.C_ON=1'b1;
    defparam un7_spon_cry_10_c_LC_6_12_2.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_10_c_LC_6_12_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_10_c_LC_6_12_2 (
            .in0(_gnd_net_),
            .in1(N__37932),
            .in2(N__35655),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_9),
            .carryout(un7_spon_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_11_c_LC_6_12_3.C_ON=1'b1;
    defparam un7_spon_cry_11_c_LC_6_12_3.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_11_c_LC_6_12_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_11_c_LC_6_12_3 (
            .in0(_gnd_net_),
            .in1(N__35536),
            .in2(N__37968),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_10),
            .carryout(un7_spon_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_12_c_LC_6_12_4.C_ON=1'b1;
    defparam un7_spon_cry_12_c_LC_6_12_4.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_12_c_LC_6_12_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_12_c_LC_6_12_4 (
            .in0(_gnd_net_),
            .in1(N__37936),
            .in2(N__35414),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_11),
            .carryout(un7_spon_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_13_c_LC_6_12_5.C_ON=1'b1;
    defparam un7_spon_cry_13_c_LC_6_12_5.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_13_c_LC_6_12_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_13_c_LC_6_12_5 (
            .in0(_gnd_net_),
            .in1(N__35315),
            .in2(N__37969),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_12),
            .carryout(un7_spon_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_14_c_LC_6_12_6.C_ON=1'b1;
    defparam un7_spon_cry_14_c_LC_6_12_6.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_14_c_LC_6_12_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_14_c_LC_6_12_6 (
            .in0(_gnd_net_),
            .in1(N__37940),
            .in2(N__35204),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_13),
            .carryout(un7_spon_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_15_c_LC_6_12_7.C_ON=1'b1;
    defparam un7_spon_cry_15_c_LC_6_12_7.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_15_c_LC_6_12_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_15_c_LC_6_12_7 (
            .in0(_gnd_net_),
            .in1(N__36655),
            .in2(N__37970),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_14),
            .carryout(un7_spon_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_16_c_LC_6_13_0.C_ON=1'b1;
    defparam un7_spon_cry_16_c_LC_6_13_0.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_16_c_LC_6_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_16_c_LC_6_13_0 (
            .in0(_gnd_net_),
            .in1(N__37912),
            .in2(N__36545),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(un7_spon_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_17_c_LC_6_13_1.C_ON=1'b1;
    defparam un7_spon_cry_17_c_LC_6_13_1.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_17_c_LC_6_13_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_17_c_LC_6_13_1 (
            .in0(_gnd_net_),
            .in1(N__36441),
            .in2(N__37964),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_16),
            .carryout(un7_spon_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_18_c_LC_6_13_2.C_ON=1'b1;
    defparam un7_spon_cry_18_c_LC_6_13_2.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_18_c_LC_6_13_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_18_c_LC_6_13_2 (
            .in0(_gnd_net_),
            .in1(N__37916),
            .in2(N__36348),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_17),
            .carryout(un7_spon_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_19_c_LC_6_13_3.C_ON=1'b1;
    defparam un7_spon_cry_19_c_LC_6_13_3.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_19_c_LC_6_13_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_19_c_LC_6_13_3 (
            .in0(_gnd_net_),
            .in1(N__36251),
            .in2(N__37965),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_18),
            .carryout(un7_spon_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_20_c_LC_6_13_4.C_ON=1'b1;
    defparam un7_spon_cry_20_c_LC_6_13_4.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_20_c_LC_6_13_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_20_c_LC_6_13_4 (
            .in0(_gnd_net_),
            .in1(N__37920),
            .in2(N__36171),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_19),
            .carryout(un7_spon_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_21_c_LC_6_13_5.C_ON=1'b1;
    defparam un7_spon_cry_21_c_LC_6_13_5.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_21_c_LC_6_13_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_21_c_LC_6_13_5 (
            .in0(_gnd_net_),
            .in1(N__36079),
            .in2(N__37966),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_20),
            .carryout(un7_spon_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_22_c_LC_6_13_6.C_ON=1'b1;
    defparam un7_spon_cry_22_c_LC_6_13_6.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_22_c_LC_6_13_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_22_c_LC_6_13_6 (
            .in0(_gnd_net_),
            .in1(N__37924),
            .in2(N__35996),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_21),
            .carryout(un7_spon_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un7_spon_cry_23_c_LC_6_13_7.C_ON=1'b1;
    defparam un7_spon_cry_23_c_LC_6_13_7.SEQ_MODE=4'b0000;
    defparam un7_spon_cry_23_c_LC_6_13_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un7_spon_cry_23_c_LC_6_13_7 (
            .in0(_gnd_net_),
            .in1(N__37079),
            .in2(N__37967),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un7_spon_cry_22),
            .carryout(un7_spon_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pon_obuf_RNO_LC_6_14_0.C_ON=1'b0;
    defparam pon_obuf_RNO_LC_6_14_0.SEQ_MODE=4'b0000;
    defparam pon_obuf_RNO_LC_6_14_0.LUT_INIT=16'b0000000011101110;
    LogicCell40 pon_obuf_RNO_LC_6_14_0 (
            .in0(N__36956),
            .in1(N__36840),
            .in2(_gnd_net_),
            .in3(N__21921),
            .lcout(pon_obuf_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_0_LC_6_15_3.C_ON=1'b0;
    defparam sTrigCounter_0_LC_6_15_3.SEQ_MODE=4'b1000;
    defparam sTrigCounter_0_LC_6_15_3.LUT_INIT=16'b1100110010011100;
    LogicCell40 sTrigCounter_0_LC_6_15_3 (
            .in0(N__22167),
            .in1(N__31350),
            .in2(N__32590),
            .in3(N__21891),
            .lcout(sTrigCounterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47844),
            .ce(),
            .sr(N__27541));
    defparam sTrigCounter_RNO_0_0_LC_6_16_2.C_ON=1'b0;
    defparam sTrigCounter_RNO_0_0_LC_6_16_2.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_0_0_LC_6_16_2.LUT_INIT=16'b0100110011001100;
    LogicCell40 sTrigCounter_RNO_0_0_LC_6_16_2 (
            .in0(N__24384),
            .in1(N__21900),
            .in2(N__24310),
            .in3(N__24720),
            .lcout(g1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sSPI_MSB0LSB1_RNIFIB13_LC_6_17_4.C_ON=1'b0;
    defparam sSPI_MSB0LSB1_RNIFIB13_LC_6_17_4.SEQ_MODE=4'b0000;
    defparam sSPI_MSB0LSB1_RNIFIB13_LC_6_17_4.LUT_INIT=16'b1011101000010000;
    LogicCell40 sSPI_MSB0LSB1_RNIFIB13_LC_6_17_4 (
            .in0(N__32175),
            .in1(N__27981),
            .in2(N__27912),
            .in3(N__22347),
            .lcout(un1_spi_data_miso_0_sqmuxa_1_i_0_N_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4Q_13_LC_7_4_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4Q_13_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4Q_13_LC_7_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4Q_13_LC_7_4_5  (
            .in0(N__22630),
            .in1(N__23565),
            .in2(_gnd_net_),
            .in3(N__22404),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIMH4QZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01_1_LC_7_4_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01_1_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01_1_LC_7_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01_1_LC_7_4_6  (
            .in0(N__22410),
            .in1(N__22428),
            .in2(_gnd_net_),
            .in3(N__22629),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNI74V01Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEESingleCont_er_LC_7_5_3.C_ON=1'b0;
    defparam sEESingleCont_er_LC_7_5_3.SEQ_MODE=4'b1010;
    defparam sEESingleCont_er_LC_7_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEESingleCont_er_LC_7_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51203),
            .lcout(sEESingleContZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47849),
            .ce(N__21930),
            .sr(N__53121));
    defparam sTrigCounter_RNO_5_5_LC_7_6_0.C_ON=1'b0;
    defparam sTrigCounter_RNO_5_5_LC_7_6_0.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_5_5_LC_7_6_0.LUT_INIT=16'b1111110001010100;
    LogicCell40 sTrigCounter_RNO_5_5_LC_7_6_0 (
            .in0(N__29106),
            .in1(N__24507),
            .in2(N__23628),
            .in3(N__24942),
            .lcout(g0_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI3LPL3_3_LC_7_6_3 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI3LPL3_3_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI3LPL3_3_LC_7_6_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_RNI3LPL3_3_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__21966),
            .in2(_gnd_net_),
            .in3(N__21949),
            .lcout(\spi_master_inst.sclk_gen_u0.N_150_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEESingleCont_er_RNO_LC_7_6_7.C_ON=1'b0;
    defparam sEESingleCont_er_RNO_LC_7_6_7.SEQ_MODE=4'b0000;
    defparam sEESingleCont_er_RNO_LC_7_6_7.LUT_INIT=16'b0000001000000000;
    LogicCell40 sEESingleCont_er_RNO_LC_7_6_7 (
            .in0(N__43287),
            .in1(N__31107),
            .in2(N__44469),
            .in3(N__44751),
            .lcout(sEESingleCont_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_4_2_LC_7_7_1.C_ON=1'b0;
    defparam sTrigCounter_RNO_4_2_LC_7_7_1.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_4_2_LC_7_7_1.LUT_INIT=16'b1111010111000100;
    LogicCell40 sTrigCounter_RNO_4_2_LC_7_7_1 (
            .in0(N__29101),
            .in1(N__24429),
            .in2(N__24938),
            .in3(N__24467),
            .lcout(g0_2_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_prev_LC_7_7_2.C_ON=1'b0;
    defparam trig_prev_LC_7_7_2.SEQ_MODE=4'b1010;
    defparam trig_prev_LC_7_7_2.LUT_INIT=16'b1111111111101110;
    LogicCell40 trig_prev_LC_7_7_2 (
            .in0(N__23972),
            .in1(N__23899),
            .in2(_gnd_net_),
            .in3(N__24059),
            .lcout(trig_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47837),
            .ce(),
            .sr(N__53092));
    defparam trig_ft_ibuf_RNIM2UO_LC_7_7_3.C_ON=1'b0;
    defparam trig_ft_ibuf_RNIM2UO_LC_7_7_3.SEQ_MODE=4'b0000;
    defparam trig_ft_ibuf_RNIM2UO_LC_7_7_3.LUT_INIT=16'b1111111100000001;
    LogicCell40 trig_ft_ibuf_RNIM2UO_LC_7_7_3 (
            .in0(N__24058),
            .in1(N__23971),
            .in2(N__23906),
            .in3(N__24464),
            .lcout(N_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_3_3_LC_7_7_4.C_ON=1'b0;
    defparam sTrigCounter_RNO_3_3_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_3_3_LC_7_7_4.LUT_INIT=16'b1100100011111010;
    LogicCell40 sTrigCounter_RNO_3_3_LC_7_7_4 (
            .in0(N__24465),
            .in1(N__24910),
            .in2(N__22023),
            .in3(N__29099),
            .lcout(g1_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_4_3_LC_7_7_5.C_ON=1'b0;
    defparam sTrigCounter_RNO_4_3_LC_7_7_5.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_4_3_LC_7_7_5.LUT_INIT=16'b1111010111000100;
    LogicCell40 sTrigCounter_RNO_4_3_LC_7_7_5 (
            .in0(N__29102),
            .in1(N__22022),
            .in2(N__24939),
            .in3(N__24468),
            .lcout(g0_2_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_3_4_LC_7_7_6.C_ON=1'b0;
    defparam sTrigCounter_RNO_3_4_LC_7_7_6.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_3_4_LC_7_7_6.LUT_INIT=16'b1100100011111010;
    LogicCell40 sTrigCounter_RNO_3_4_LC_7_7_6 (
            .in0(N__24466),
            .in1(N__24911),
            .in2(N__22008),
            .in3(N__29100),
            .lcout(g1_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_5_4_LC_7_7_7.C_ON=1'b0;
    defparam sTrigCounter_RNO_5_4_LC_7_7_7.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_5_4_LC_7_7_7.LUT_INIT=16'b1111010111000100;
    LogicCell40 sTrigCounter_RNO_5_4_LC_7_7_7 (
            .in0(N__29103),
            .in1(N__22007),
            .in2(N__24940),
            .in3(N__24469),
            .lcout(g0_2_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_4_5_LC_7_8_0.C_ON=1'b0;
    defparam sTrigCounter_RNO_4_5_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_4_5_LC_7_8_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 sTrigCounter_RNO_4_5_LC_7_8_0 (
            .in0(N__24229),
            .in1(N__24203),
            .in2(N__32623),
            .in3(N__24602),
            .lcout(),
            .ltout(g1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_1_5_LC_7_8_1.C_ON=1'b0;
    defparam sTrigCounter_RNO_1_5_LC_7_8_1.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_1_5_LC_7_8_1.LUT_INIT=16'b1100000000000000;
    LogicCell40 sTrigCounter_RNO_1_5_LC_7_8_1 (
            .in0(_gnd_net_),
            .in1(N__31299),
            .in2(N__21993),
            .in3(N__31387),
            .lcout(g1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPointerReset_LC_7_8_5.C_ON=1'b0;
    defparam sEEPointerReset_LC_7_8_5.SEQ_MODE=4'b1000;
    defparam sEEPointerReset_LC_7_8_5.LUT_INIT=16'b1000100011110000;
    LogicCell40 sEEPointerReset_LC_7_8_5 (
            .in0(N__51257),
            .in1(N__43855),
            .in2(N__33391),
            .in3(N__28959),
            .lcout(sEEPointerResetZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47828),
            .ce(),
            .sr(_gnd_net_));
    defparam sPeriod_prev_RNIRSLG_LC_7_8_6.C_ON=1'b0;
    defparam sPeriod_prev_RNIRSLG_LC_7_8_6.SEQ_MODE=4'b0000;
    defparam sPeriod_prev_RNIRSLG_LC_7_8_6.LUT_INIT=16'b0011001111111111;
    LogicCell40 sPeriod_prev_RNIRSLG_LC_7_8_6 (
            .in0(_gnd_net_),
            .in1(N__24257),
            .in2(_gnd_net_),
            .in3(N__24361),
            .lcout(un1_reset_rpi_inv_2_i_o3_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPeriod_0_LC_7_9_0.C_ON=1'b0;
    defparam sEEPeriod_0_LC_7_9_0.SEQ_MODE=4'b1010;
    defparam sEEPeriod_0_LC_7_9_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPeriod_0_LC_7_9_0 (
            .in0(N__51259),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47820),
            .ce(N__24519),
            .sr(N__53069));
    defparam sEEPeriod_1_LC_7_9_1.C_ON=1'b0;
    defparam sEEPeriod_1_LC_7_9_1.SEQ_MODE=4'b1010;
    defparam sEEPeriod_1_LC_7_9_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPeriod_1_LC_7_9_1 (
            .in0(N__50592),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47820),
            .ce(N__24519),
            .sr(N__53069));
    defparam sEEPeriod_2_LC_7_9_2.C_ON=1'b0;
    defparam sEEPeriod_2_LC_7_9_2.SEQ_MODE=4'b1010;
    defparam sEEPeriod_2_LC_7_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_2_LC_7_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50282),
            .lcout(sEEPeriodZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47820),
            .ce(N__24519),
            .sr(N__53069));
    defparam sEEPeriod_3_LC_7_9_3.C_ON=1'b0;
    defparam sEEPeriod_3_LC_7_9_3.SEQ_MODE=4'b1010;
    defparam sEEPeriod_3_LC_7_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_3_LC_7_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49820),
            .lcout(sEEPeriodZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47820),
            .ce(N__24519),
            .sr(N__53069));
    defparam sEEPeriod_4_LC_7_9_4.C_ON=1'b0;
    defparam sEEPeriod_4_LC_7_9_4.SEQ_MODE=4'b1010;
    defparam sEEPeriod_4_LC_7_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_4_LC_7_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49354),
            .lcout(sEEPeriodZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47820),
            .ce(N__24519),
            .sr(N__53069));
    defparam sEEPeriod_5_LC_7_9_5.C_ON=1'b0;
    defparam sEEPeriod_5_LC_7_9_5.SEQ_MODE=4'b1011;
    defparam sEEPeriod_5_LC_7_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_5_LC_7_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47063),
            .lcout(sEEPeriodZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47820),
            .ce(N__24519),
            .sr(N__53069));
    defparam sEEPeriod_6_LC_7_9_6.C_ON=1'b0;
    defparam sEEPeriod_6_LC_7_9_6.SEQ_MODE=4'b1010;
    defparam sEEPeriod_6_LC_7_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_6_LC_7_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48153),
            .lcout(sEEPeriodZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47820),
            .ce(N__24519),
            .sr(N__53069));
    defparam sEEPeriod_7_LC_7_9_7.C_ON=1'b0;
    defparam sEEPeriod_7_LC_7_9_7.SEQ_MODE=4'b1011;
    defparam sEEPeriod_7_LC_7_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_7_LC_7_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48776),
            .lcout(sEEPeriodZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47820),
            .ce(N__24519),
            .sr(N__53069));
    defparam sTrigCounter_RNO_3_1_LC_7_10_0.C_ON=1'b0;
    defparam sTrigCounter_RNO_3_1_LC_7_10_0.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_3_1_LC_7_10_0.LUT_INIT=16'b1100100011111010;
    LogicCell40 sTrigCounter_RNO_3_1_LC_7_10_0 (
            .in0(N__24490),
            .in1(N__24878),
            .in2(N__22133),
            .in3(N__29097),
            .lcout(g1_0_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigInternal_prev_LC_7_10_1.C_ON=1'b0;
    defparam sEETrigInternal_prev_LC_7_10_1.SEQ_MODE=4'b1010;
    defparam sEETrigInternal_prev_LC_7_10_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEETrigInternal_prev_LC_7_10_1 (
            .in0(N__29098),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEETrigInternal_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47812),
            .ce(),
            .sr(N__53058));
    defparam sEETrigInternal_prev_RNISEUG_LC_7_10_2.C_ON=1'b0;
    defparam sEETrigInternal_prev_RNISEUG_LC_7_10_2.SEQ_MODE=4'b0000;
    defparam sEETrigInternal_prev_RNISEUG_LC_7_10_2.LUT_INIT=16'b0011001100000000;
    LogicCell40 sEETrigInternal_prev_RNISEUG_LC_7_10_2 (
            .in0(_gnd_net_),
            .in1(N__24874),
            .in2(_gnd_net_),
            .in3(N__29095),
            .lcout(),
            .ltout(sEETrigInternal_prev_RNISEUGZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigInternal_RNIOMLD1_LC_7_10_3.C_ON=1'b0;
    defparam sTrigInternal_RNIOMLD1_LC_7_10_3.SEQ_MODE=4'b0000;
    defparam sTrigInternal_RNIOMLD1_LC_7_10_3.LUT_INIT=16'b0000001100000010;
    LogicCell40 sTrigInternal_RNIOMLD1_LC_7_10_3 (
            .in0(N__22040),
            .in1(N__22280),
            .in2(N__22026),
            .in3(N__24491),
            .lcout(sTrigInternal_RNIOMLDZ0Z1),
            .ltout(sTrigInternal_RNIOMLDZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigInternal_RNO_0_LC_7_10_4.C_ON=1'b0;
    defparam sTrigInternal_RNO_0_LC_7_10_4.SEQ_MODE=4'b0000;
    defparam sTrigInternal_RNO_0_LC_7_10_4.LUT_INIT=16'b0100010011100100;
    LogicCell40 sTrigInternal_RNO_0_LC_7_10_4 (
            .in0(N__36958),
            .in1(N__36859),
            .in2(N__22053),
            .in3(N__24816),
            .lcout(),
            .ltout(sTrigInternal_RNOZ0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigInternal_LC_7_10_5.C_ON=1'b0;
    defparam sTrigInternal_LC_7_10_5.SEQ_MODE=4'b1010;
    defparam sTrigInternal_LC_7_10_5.LUT_INIT=16'b0000011100000011;
    LogicCell40 sTrigInternal_LC_7_10_5 (
            .in0(N__24740),
            .in1(N__22050),
            .in2(N__22044),
            .in3(N__24718),
            .lcout(sTrigInternalZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47812),
            .ce(),
            .sr(N__53058));
    defparam trig_prev_RNIIHS91_LC_7_10_7.C_ON=1'b0;
    defparam trig_prev_RNIIHS91_LC_7_10_7.SEQ_MODE=4'b0000;
    defparam trig_prev_RNIIHS91_LC_7_10_7.LUT_INIT=16'b1111010111000100;
    LogicCell40 trig_prev_RNIIHS91_LC_7_10_7 (
            .in0(N__29096),
            .in1(N__22041),
            .in2(N__24909),
            .in3(N__24489),
            .lcout(N_127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPeriod_16_LC_7_11_0.C_ON=1'b0;
    defparam sEEPeriod_16_LC_7_11_0.SEQ_MODE=4'b1011;
    defparam sEEPeriod_16_LC_7_11_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPeriod_16_LC_7_11_0 (
            .in0(N__51260),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47803),
            .ce(N__28923),
            .sr(N__53048));
    defparam sEEPeriod_17_LC_7_11_1.C_ON=1'b0;
    defparam sEEPeriod_17_LC_7_11_1.SEQ_MODE=4'b1010;
    defparam sEEPeriod_17_LC_7_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_17_LC_7_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50599),
            .lcout(sEEPeriodZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47803),
            .ce(N__28923),
            .sr(N__53048));
    defparam sEEPeriod_18_LC_7_11_2.C_ON=1'b0;
    defparam sEEPeriod_18_LC_7_11_2.SEQ_MODE=4'b1010;
    defparam sEEPeriod_18_LC_7_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_18_LC_7_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50284),
            .lcout(sEEPeriodZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47803),
            .ce(N__28923),
            .sr(N__53048));
    defparam sEEPeriod_19_LC_7_11_3.C_ON=1'b0;
    defparam sEEPeriod_19_LC_7_11_3.SEQ_MODE=4'b1010;
    defparam sEEPeriod_19_LC_7_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_19_LC_7_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49822),
            .lcout(sEEPeriodZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47803),
            .ce(N__28923),
            .sr(N__53048));
    defparam sEEPeriod_20_LC_7_11_4.C_ON=1'b0;
    defparam sEEPeriod_20_LC_7_11_4.SEQ_MODE=4'b1010;
    defparam sEEPeriod_20_LC_7_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_20_LC_7_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49346),
            .lcout(sEEPeriodZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47803),
            .ce(N__28923),
            .sr(N__53048));
    defparam sEEPeriod_21_LC_7_11_5.C_ON=1'b0;
    defparam sEEPeriod_21_LC_7_11_5.SEQ_MODE=4'b1010;
    defparam sEEPeriod_21_LC_7_11_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPeriod_21_LC_7_11_5 (
            .in0(N__47064),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47803),
            .ce(N__28923),
            .sr(N__53048));
    defparam sEEPeriod_22_LC_7_11_6.C_ON=1'b0;
    defparam sEEPeriod_22_LC_7_11_6.SEQ_MODE=4'b1010;
    defparam sEEPeriod_22_LC_7_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_22_LC_7_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48305),
            .lcout(sEEPeriodZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47803),
            .ce(N__28923),
            .sr(N__53048));
    defparam sEEPeriod_23_LC_7_11_7.C_ON=1'b0;
    defparam sEEPeriod_23_LC_7_11_7.SEQ_MODE=4'b1010;
    defparam sEEPeriod_23_LC_7_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_23_LC_7_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48769),
            .lcout(sEEPeriodZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47803),
            .ce(N__28923),
            .sr(N__53048));
    defparam sTrigCounter_RNO_4_1_LC_7_12_0.C_ON=1'b0;
    defparam sTrigCounter_RNO_4_1_LC_7_12_0.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_4_1_LC_7_12_0.LUT_INIT=16'b1111010111000100;
    LogicCell40 sTrigCounter_RNO_4_1_LC_7_12_0 (
            .in0(N__29105),
            .in1(N__22134),
            .in2(N__24945),
            .in3(N__24509),
            .lcout(g0_2_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNI743O1_18_LC_7_12_1.C_ON=1'b0;
    defparam sCounter_RNI743O1_18_LC_7_12_1.SEQ_MODE=4'b0000;
    defparam sCounter_RNI743O1_18_LC_7_12_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNI743O1_18_LC_7_12_1 (
            .in0(N__22110),
            .in1(N__36253),
            .in2(N__23031),
            .in3(N__36332),
            .lcout(),
            .ltout(un1_reset_rpi_inv_2_i_o3_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIRQR25_10_LC_7_12_2.C_ON=1'b0;
    defparam sCounter_RNIRQR25_10_LC_7_12_2.SEQ_MODE=4'b0000;
    defparam sCounter_RNIRQR25_10_LC_7_12_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNIRQR25_10_LC_7_12_2 (
            .in0(N__22068),
            .in1(N__24972),
            .in2(N__22101),
            .in3(N__22185),
            .lcout(N_1479),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_3_0_LC_7_12_3.C_ON=1'b0;
    defparam sTrigCounter_RNO_3_0_LC_7_12_3.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_3_0_LC_7_12_3.LUT_INIT=16'b1100100011111010;
    LogicCell40 sTrigCounter_RNO_3_0_LC_7_12_3 (
            .in0(N__24508),
            .in1(N__24934),
            .in2(N__22098),
            .in3(N__29104),
            .lcout(g0_2_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_1_2_LC_7_12_5.C_ON=1'b0;
    defparam sTrigCounter_RNO_1_2_LC_7_12_5.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_1_2_LC_7_12_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 sTrigCounter_RNO_1_2_LC_7_12_5 (
            .in0(N__31280),
            .in1(N__32595),
            .in2(_gnd_net_),
            .in3(N__31363),
            .lcout(g1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNI6K4L_16_LC_7_12_7.C_ON=1'b0;
    defparam sCounter_RNI6K4L_16_LC_7_12_7.SEQ_MODE=4'b0000;
    defparam sCounter_RNI6K4L_16_LC_7_12_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNI6K4L_16_LC_7_12_7 (
            .in0(N__36529),
            .in1(N__36654),
            .in2(N__35202),
            .in3(N__36430),
            .lcout(un1_reset_rpi_inv_2_i_o3_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_2_1_LC_7_13_1.C_ON=1'b0;
    defparam sTrigCounter_RNO_2_1_LC_7_13_1.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_2_1_LC_7_13_1.LUT_INIT=16'b0100010011100100;
    LogicCell40 sTrigCounter_RNO_2_1_LC_7_13_1 (
            .in0(N__36934),
            .in1(N__36813),
            .in2(N__22062),
            .in3(N__24798),
            .lcout(g2_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_2_LC_7_13_2.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_2_LC_7_13_2.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_2_LC_7_13_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_2_LC_7_13_2 (
            .in0(N__22311),
            .in1(N__22323),
            .in2(N__22341),
            .in3(N__25185),
            .lcout(),
            .ltout(sbuttonModeStatus_0_sqmuxa_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_LC_7_13_3.C_ON=1'b0;
    defparam sbuttonModeStatus_LC_7_13_3.SEQ_MODE=4'b1000;
    defparam sbuttonModeStatus_LC_7_13_3.LUT_INIT=16'b0110110011001100;
    LogicCell40 sbuttonModeStatus_LC_7_13_3 (
            .in0(N__23013),
            .in1(N__22205),
            .in2(N__22218),
            .in3(N__25248),
            .lcout(sbuttonModeStatusZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53276),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_1_1_LC_7_13_5.C_ON=1'b0;
    defparam sTrigCounter_RNO_1_1_LC_7_13_5.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_1_1_LC_7_13_5.LUT_INIT=16'b0100110011001100;
    LogicCell40 sTrigCounter_RNO_1_1_LC_7_13_5 (
            .in0(N__24380),
            .in1(N__22194),
            .in2(N__24309),
            .in3(N__24719),
            .lcout(g1_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIOUF02_23_LC_7_13_7.C_ON=1'b0;
    defparam sCounter_RNIOUF02_23_LC_7_13_7.SEQ_MODE=4'b0000;
    defparam sCounter_RNIOUF02_23_LC_7_13_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNIOUF02_23_LC_7_13_7 (
            .in0(N__37075),
            .in1(N__34452),
            .in2(N__23022),
            .in3(N__34574),
            .lcout(un1_reset_rpi_inv_2_i_o3_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIJ0NP_17_LC_7_14_1.C_ON=1'b0;
    defparam sCounter_RNIJ0NP_17_LC_7_14_1.SEQ_MODE=4'b0000;
    defparam sCounter_RNIJ0NP_17_LC_7_14_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNIJ0NP_17_LC_7_14_1 (
            .in0(N__36629),
            .in1(N__35163),
            .in2(N__36443),
            .in3(N__36805),
            .lcout(op_gt_op_gt_un13_striginternallto23_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_1_0_LC_7_14_2.C_ON=1'b0;
    defparam sTrigCounter_RNO_1_0_LC_7_14_2.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_1_0_LC_7_14_2.LUT_INIT=16'b0010001011100010;
    LogicCell40 sTrigCounter_RNO_1_0_LC_7_14_2 (
            .in0(N__36806),
            .in1(N__36955),
            .in2(N__22179),
            .in3(N__24797),
            .lcout(g2_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_0_1_LC_7_14_4.C_ON=1'b0;
    defparam sTrigCounter_RNO_0_1_LC_7_14_4.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_0_1_LC_7_14_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 sTrigCounter_RNO_0_1_LC_7_14_4 (
            .in0(N__32631),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31349),
            .lcout(),
            .ltout(g1_0_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_1_LC_7_14_5.C_ON=1'b0;
    defparam sTrigCounter_1_LC_7_14_5.SEQ_MODE=4'b1000;
    defparam sTrigCounter_1_LC_7_14_5.LUT_INIT=16'b1010101010011010;
    LogicCell40 sTrigCounter_1_LC_7_14_5 (
            .in0(N__31262),
            .in1(N__22161),
            .in2(N__22155),
            .in3(N__22152),
            .lcout(sTrigCounterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47829),
            .ce(),
            .sr(N__27543));
    defparam sCounter_RNIVUR25_10_LC_7_15_0.C_ON=1'b0;
    defparam sCounter_RNIVUR25_10_LC_7_15_0.SEQ_MODE=4'b0000;
    defparam sCounter_RNIVUR25_10_LC_7_15_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 sCounter_RNIVUR25_10_LC_7_15_0 (
            .in0(N__24987),
            .in1(N__22239),
            .in2(N__22146),
            .in3(N__22296),
            .lcout(op_gt_op_gt_un13_striginternal_0),
            .ltout(op_gt_op_gt_un13_striginternal_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigInternal_RNIMEFL5_LC_7_15_1.C_ON=1'b0;
    defparam sTrigInternal_RNIMEFL5_LC_7_15_1.SEQ_MODE=4'b0000;
    defparam sTrigInternal_RNIMEFL5_LC_7_15_1.LUT_INIT=16'b0111011101110101;
    LogicCell40 sTrigInternal_RNIMEFL5_LC_7_15_1 (
            .in0(N__32633),
            .in1(N__22289),
            .in2(N__22137),
            .in3(N__24799),
            .lcout(LED_ACQ_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIAME71_8_LC_7_15_2.C_ON=1'b0;
    defparam sCounter_RNIAME71_8_LC_7_15_2.SEQ_MODE=4'b0000;
    defparam sCounter_RNIAME71_8_LC_7_15_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNIAME71_8_LC_7_15_2 (
            .in0(N__35738),
            .in1(N__34454),
            .in2(N__34594),
            .in3(N__35849),
            .lcout(),
            .ltout(op_gt_op_gt_un13_striginternallto23_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIQVE02_16_LC_7_15_3.C_ON=1'b0;
    defparam sCounter_RNIQVE02_16_LC_7_15_3.SEQ_MODE=4'b0000;
    defparam sCounter_RNIQVE02_16_LC_7_15_3.LUT_INIT=16'b0000000000010000;
    LogicCell40 sCounter_RNIQVE02_16_LC_7_15_3 (
            .in0(N__36525),
            .in1(N__34700),
            .in2(N__22299),
            .in3(N__34834),
            .lcout(op_gt_op_gt_un13_striginternallto23_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LED_ACQ_obuf_RNO_LC_7_15_4.C_ON=1'b0;
    defparam LED_ACQ_obuf_RNO_LC_7_15_4.SEQ_MODE=4'b0000;
    defparam LED_ACQ_obuf_RNO_LC_7_15_4.LUT_INIT=16'b1000100010001100;
    LogicCell40 LED_ACQ_obuf_RNO_LC_7_15_4 (
            .in0(N__22290),
            .in1(N__32632),
            .in2(N__22269),
            .in3(N__24822),
            .lcout(LED_ACQ_obuf_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNISQHJ1_18_LC_7_15_5.C_ON=1'b0;
    defparam sCounter_RNISQHJ1_18_LC_7_15_5.SEQ_MODE=4'b0000;
    defparam sCounter_RNISQHJ1_18_LC_7_15_5.LUT_INIT=16'b0000000000100000;
    LogicCell40 sCounter_RNISQHJ1_18_LC_7_15_5 (
            .in0(N__25488),
            .in1(N__36228),
            .in2(N__24960),
            .in3(N__36309),
            .lcout(op_gt_op_gt_un13_striginternallto23_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterRAM_0_LC_7_16_0.C_ON=1'b1;
    defparam sCounterRAM_0_LC_7_16_0.SEQ_MODE=4'b1010;
    defparam sCounterRAM_0_LC_7_16_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_0_LC_7_16_0 (
            .in0(N__22373),
            .in1(N__27392),
            .in2(_gnd_net_),
            .in3(N__22233),
            .lcout(sCounterRAMZ0Z_0),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(sCounterRAM_cry_0),
            .clk(N__47845),
            .ce(),
            .sr(N__53007));
    defparam sCounterRAM_1_LC_7_16_1.C_ON=1'b1;
    defparam sCounterRAM_1_LC_7_16_1.SEQ_MODE=4'b1010;
    defparam sCounterRAM_1_LC_7_16_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_1_LC_7_16_1 (
            .in0(N__22377),
            .in1(N__28013),
            .in2(_gnd_net_),
            .in3(N__22230),
            .lcout(sCounterRAMZ0Z_1),
            .ltout(),
            .carryin(sCounterRAM_cry_0),
            .carryout(sCounterRAM_cry_1),
            .clk(N__47845),
            .ce(),
            .sr(N__53007));
    defparam sCounterRAM_2_LC_7_16_2.C_ON=1'b1;
    defparam sCounterRAM_2_LC_7_16_2.SEQ_MODE=4'b1010;
    defparam sCounterRAM_2_LC_7_16_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_2_LC_7_16_2 (
            .in0(N__22374),
            .in1(N__28034),
            .in2(_gnd_net_),
            .in3(N__22227),
            .lcout(sCounterRAMZ0Z_2),
            .ltout(),
            .carryin(sCounterRAM_cry_1),
            .carryout(sCounterRAM_cry_2),
            .clk(N__47845),
            .ce(),
            .sr(N__53007));
    defparam sCounterRAM_3_LC_7_16_3.C_ON=1'b1;
    defparam sCounterRAM_3_LC_7_16_3.SEQ_MODE=4'b1010;
    defparam sCounterRAM_3_LC_7_16_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_3_LC_7_16_3 (
            .in0(N__22378),
            .in1(N__25307),
            .in2(_gnd_net_),
            .in3(N__22224),
            .lcout(sCounterRAMZ0Z_3),
            .ltout(),
            .carryin(sCounterRAM_cry_2),
            .carryout(sCounterRAM_cry_3),
            .clk(N__47845),
            .ce(),
            .sr(N__53007));
    defparam sCounterRAM_4_LC_7_16_4.C_ON=1'b1;
    defparam sCounterRAM_4_LC_7_16_4.SEQ_MODE=4'b1010;
    defparam sCounterRAM_4_LC_7_16_4.LUT_INIT=16'b0000010101010000;
    LogicCell40 sCounterRAM_4_LC_7_16_4 (
            .in0(N__22375),
            .in1(_gnd_net_),
            .in2(N__27437),
            .in3(N__22221),
            .lcout(sCounterRAMZ0Z_4),
            .ltout(),
            .carryin(sCounterRAM_cry_3),
            .carryout(sCounterRAM_cry_4),
            .clk(N__47845),
            .ce(),
            .sr(N__53007));
    defparam sCounterRAM_5_LC_7_16_5.C_ON=1'b1;
    defparam sCounterRAM_5_LC_7_16_5.SEQ_MODE=4'b1010;
    defparam sCounterRAM_5_LC_7_16_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_5_LC_7_16_5 (
            .in0(N__22379),
            .in1(N__27452),
            .in2(_gnd_net_),
            .in3(N__22386),
            .lcout(sCounterRAMZ0Z_5),
            .ltout(),
            .carryin(sCounterRAM_cry_4),
            .carryout(sCounterRAM_cry_5),
            .clk(N__47845),
            .ce(),
            .sr(N__53007));
    defparam sCounterRAM_6_LC_7_16_6.C_ON=1'b1;
    defparam sCounterRAM_6_LC_7_16_6.SEQ_MODE=4'b1010;
    defparam sCounterRAM_6_LC_7_16_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_6_LC_7_16_6 (
            .in0(N__22376),
            .in1(N__25323),
            .in2(_gnd_net_),
            .in3(N__22383),
            .lcout(sCounterRAMZ0Z_6),
            .ltout(),
            .carryin(sCounterRAM_cry_5),
            .carryout(sCounterRAM_cry_6),
            .clk(N__47845),
            .ce(),
            .sr(N__53007));
    defparam sCounterRAM_7_LC_7_16_7.C_ON=1'b0;
    defparam sCounterRAM_7_LC_7_16_7.SEQ_MODE=4'b1010;
    defparam sCounterRAM_7_LC_7_16_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterRAM_7_LC_7_16_7 (
            .in0(N__22380),
            .in1(N__27410),
            .in2(_gnd_net_),
            .in3(N__22350),
            .lcout(sCounterRAMZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47845),
            .ce(),
            .sr(N__53007));
    defparam RAM_DATA_cl_10_15_LC_7_17_0.C_ON=1'b0;
    defparam RAM_DATA_cl_10_15_LC_7_17_0.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_10_15_LC_7_17_0.LUT_INIT=16'b0010000000000000;
    LogicCell40 RAM_DATA_cl_10_15_LC_7_17_0 (
            .in0(N__31944),
            .in1(N__26610),
            .in2(N__32676),
            .in3(N__32177),
            .lcout(RAM_DATA_cl_10Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47850),
            .ce(),
            .sr(N__52999));
    defparam sADC_clk_LC_7_17_2.C_ON=1'b0;
    defparam sADC_clk_LC_7_17_2.SEQ_MODE=4'b1010;
    defparam sADC_clk_LC_7_17_2.LUT_INIT=16'b0010100000000000;
    LogicCell40 sADC_clk_LC_7_17_2 (
            .in0(N__31943),
            .in1(N__27602),
            .in2(N__38229),
            .in3(N__32176),
            .lcout(ADC_clk_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47850),
            .ce(),
            .sr(N__52999));
    defparam sSPI_MSB0LSB1_RNIO3VP1_LC_7_17_5.C_ON=1'b0;
    defparam sSPI_MSB0LSB1_RNIO3VP1_LC_7_17_5.SEQ_MODE=4'b0000;
    defparam sSPI_MSB0LSB1_RNIO3VP1_LC_7_17_5.LUT_INIT=16'b0101010100001100;
    LogicCell40 sSPI_MSB0LSB1_RNIO3VP1_LC_7_17_5 (
            .in0(N__31693),
            .in1(N__27907),
            .in2(N__27980),
            .in3(N__31942),
            .lcout(sSPI_MSB0LSB1_RNIO3VPZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_7_LC_7_18_0.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_7_LC_7_18_0.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_7_LC_7_18_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_7_LC_7_18_0 (
            .in0(N__23468),
            .in1(N__23483),
            .in2(N__23547),
            .in3(N__23498),
            .lcout(sbuttonModeStatus_0_sqmuxa_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_5_LC_7_18_4.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_5_LC_7_18_4.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_5_LC_7_18_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_5_LC_7_18_4 (
            .in0(N__23336),
            .in1(N__23351),
            .in2(N__23322),
            .in3(N__23366),
            .lcout(sbuttonModeStatus_0_sqmuxa_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_6_LC_7_18_5.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_6_LC_7_18_5.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_6_LC_7_18_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_6_LC_7_18_5 (
            .in0(N__23273),
            .in1(N__23288),
            .in2(N__23517),
            .in3(N__23303),
            .lcout(sbuttonModeStatus_0_sqmuxa_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_14_LC_8_3_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_14_LC_8_3_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_14_LC_8_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_14_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25704),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53246),
            .ce(),
            .sr(N__53131));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_0_LC_8_4_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_0_LC_8_4_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_0_LC_8_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_0_LC_8_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28890),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53249),
            .ce(),
            .sr(N__53122));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_8_LC_8_4_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_8_LC_8_4_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_8_LC_8_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_8_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28866),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53249),
            .ce(),
            .sr(N__53122));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_9_LC_8_4_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_9_LC_8_4_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_9_LC_8_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_9_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28854),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53249),
            .ce(),
            .sr(N__53122));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_7_LC_8_4_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_7_LC_8_4_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_7_LC_8_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_7_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28878),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53249),
            .ce(),
            .sr(N__53122));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_1_LC_8_4_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_1_LC_8_4_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_1_LC_8_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_1_LC_8_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25740),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53249),
            .ce(),
            .sr(N__53122));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_13_LC_8_4_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_13_LC_8_4_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_13_LC_8_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_13_LC_8_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28752),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53249),
            .ce(),
            .sr(N__53122));
    defparam sPeriod_prev_LC_8_5_0.C_ON=1'b0;
    defparam sPeriod_prev_LC_8_5_0.SEQ_MODE=4'b1010;
    defparam sPeriod_prev_LC_8_5_0.LUT_INIT=16'b0000000011101110;
    LogicCell40 sPeriod_prev_LC_8_5_0 (
            .in0(N__36972),
            .in1(N__36877),
            .in2(_gnd_net_),
            .in3(N__24825),
            .lcout(sPeriod_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47846),
            .ce(),
            .sr(N__53107));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4Q_10_LC_8_5_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4Q_10_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4Q_10_LC_8_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4Q_10_LC_8_5_3  (
            .in0(N__23763),
            .in1(N__23586),
            .in2(_gnd_net_),
            .in3(N__22640),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIGB4QZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4Q_12_LC_8_5_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4Q_12_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4Q_12_LC_8_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4Q_12_LC_8_5_4  (
            .in0(N__22641),
            .in1(N__23571),
            .in2(_gnd_net_),
            .in3(N__23592),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_i_RNIKF4QZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_done_reg2_i_LC_8_5_6 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_reg2_i_LC_8_5_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_done_reg2_i_LC_8_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_done_reg2_i_LC_8_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28812),
            .lcout(\spi_slave_inst.rx_done_reg2_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47846),
            .ce(),
            .sr(N__53107));
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_LC_8_6_1 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_LC_8_6_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_LC_8_6_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.falling_count_start_i_LC_8_6_1  (
            .in0(N__23643),
            .in1(N__23649),
            .in2(_gnd_net_),
            .in3(N__22555),
            .lcout(\spi_master_inst.sclk_gen_u0.falling_count_start_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53253),
            .ce(),
            .sr(N__53093));
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_2_LC_8_6_2 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_2_LC_8_6_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.spim_clk_state_i_2_LC_8_6_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spim_clk_state_i_2_LC_8_6_2  (
            .in0(N__22556),
            .in1(N__23682),
            .in2(_gnd_net_),
            .in3(N__23750),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53253),
            .ce(),
            .sr(N__53093));
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_LC_8_6_4 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_LC_8_6_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.sclk_count_start_i_LC_8_6_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.sclk_count_start_i_LC_8_6_4  (
            .in0(N__22557),
            .in1(N__22513),
            .in2(N__23739),
            .in3(N__22545),
            .lcout(\spi_master_inst.sclk_gen_u0.sclk_count_start_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53253),
            .ce(),
            .sr(N__53093));
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_RNISHDJ_LC_8_6_6 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_RNISHDJ_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_RNISHDJ_LC_8_6_6 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_clk_i_RNISHDJ_LC_8_6_6  (
            .in0(N__22464),
            .in1(N__22493),
            .in2(_gnd_net_),
            .in3(N__23642),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_ie_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_LC_8_6_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_LC_8_6_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.delay_clk_i_LC_8_6_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.delay_clk_i_LC_8_6_7  (
            .in0(N__22494),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_master_inst.sclk_gen_u0.delay_clk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53253),
            .ce(),
            .sr(N__53093));
    defparam sEETrigCounter_4_LC_8_7_0.C_ON=1'b0;
    defparam sEETrigCounter_4_LC_8_7_0.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_4_LC_8_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_4_LC_8_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49361),
            .lcout(sEETrigCounterZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47830),
            .ce(N__31020),
            .sr(N__53081));
    defparam sEETrigCounter_5_LC_8_7_1.C_ON=1'b0;
    defparam sEETrigCounter_5_LC_8_7_1.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_5_LC_8_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_5_LC_8_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46970),
            .lcout(sEETrigCounterZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47830),
            .ce(N__31020),
            .sr(N__53081));
    defparam sEETrigCounter_6_LC_8_7_2.C_ON=1'b0;
    defparam sEETrigCounter_6_LC_8_7_2.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_6_LC_8_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_6_LC_8_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48146),
            .lcout(sEETrigCounterZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47830),
            .ce(N__31020),
            .sr(N__53081));
    defparam sEETrigCounter_7_LC_8_7_3.C_ON=1'b0;
    defparam sEETrigCounter_7_LC_8_7_3.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_7_LC_8_7_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEETrigCounter_7_LC_8_7_3 (
            .in0(N__48736),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEETrigCounterZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47830),
            .ce(N__31020),
            .sr(N__53081));
    defparam sTrigCounter_RNO_2_2_LC_8_8_0.C_ON=1'b0;
    defparam sTrigCounter_RNO_2_2_LC_8_8_0.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_2_2_LC_8_8_0.LUT_INIT=16'b0100010011100100;
    LogicCell40 sTrigCounter_RNO_2_2_LC_8_8_0 (
            .in0(N__36973),
            .in1(N__36848),
            .in2(N__22713),
            .in3(N__24818),
            .lcout(),
            .ltout(g2_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_2_LC_8_8_1.C_ON=1'b0;
    defparam sTrigCounter_2_LC_8_8_1.SEQ_MODE=4'b1000;
    defparam sTrigCounter_2_LC_8_8_1.LUT_INIT=16'b1010101010100110;
    LogicCell40 sTrigCounter_2_LC_8_8_1 (
            .in0(N__24611),
            .in1(N__22704),
            .in2(N__22692),
            .in3(N__22689),
            .lcout(sTrigCounterZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47821),
            .ce(),
            .sr(N__27542));
    defparam sTrigCounter_RNO_0_2_LC_8_8_2.C_ON=1'b0;
    defparam sTrigCounter_RNO_0_2_LC_8_8_2.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_0_2_LC_8_8_2.LUT_INIT=16'b0111111100000000;
    LogicCell40 sTrigCounter_RNO_0_2_LC_8_8_2 (
            .in0(N__24357),
            .in1(N__24259),
            .in2(N__24714),
            .in3(N__24405),
            .lcout(g1_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_2_3_LC_8_8_3.C_ON=1'b0;
    defparam sTrigCounter_RNO_2_3_LC_8_8_3.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_2_3_LC_8_8_3.LUT_INIT=16'b0100010011110000;
    LogicCell40 sTrigCounter_RNO_2_3_LC_8_8_3 (
            .in0(N__24817),
            .in1(N__22683),
            .in2(N__36873),
            .in3(N__36974),
            .lcout(),
            .ltout(g2_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_3_LC_8_8_4.C_ON=1'b0;
    defparam sTrigCounter_3_LC_8_8_4.SEQ_MODE=4'b1000;
    defparam sTrigCounter_3_LC_8_8_4.LUT_INIT=16'b1100110011000110;
    LogicCell40 sTrigCounter_3_LC_8_8_4 (
            .in0(N__22674),
            .in1(N__24204),
            .in2(N__22677),
            .in3(N__22659),
            .lcout(sTrigCounterZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47821),
            .ce(),
            .sr(N__27542));
    defparam sTrigCounter_RNO_1_3_LC_8_8_5.C_ON=1'b0;
    defparam sTrigCounter_RNO_1_3_LC_8_8_5.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_1_3_LC_8_8_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 sTrigCounter_RNO_1_3_LC_8_8_5 (
            .in0(N__24610),
            .in1(N__31300),
            .in2(N__32594),
            .in3(N__31388),
            .lcout(g1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_0_3_LC_8_8_6.C_ON=1'b0;
    defparam sTrigCounter_RNO_0_3_LC_8_8_6.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_0_3_LC_8_8_6.LUT_INIT=16'b0010101010101010;
    LogicCell40 sTrigCounter_RNO_0_3_LC_8_8_6 (
            .in0(N__22665),
            .in1(N__24258),
            .in2(N__24376),
            .in3(N__24703),
            .lcout(g1_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_2_4_LC_8_9_0.C_ON=1'b0;
    defparam sTrigCounter_RNO_2_4_LC_8_9_0.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_2_4_LC_8_9_0.LUT_INIT=16'b0100010011100100;
    LogicCell40 sTrigCounter_RNO_2_4_LC_8_9_0 (
            .in0(N__36959),
            .in1(N__36860),
            .in2(N__22653),
            .in3(N__24824),
            .lcout(),
            .ltout(g2_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_4_LC_8_9_1.C_ON=1'b0;
    defparam sTrigCounter_4_LC_8_9_1.SEQ_MODE=4'b1000;
    defparam sTrigCounter_4_LC_8_9_1.LUT_INIT=16'b1010101010100110;
    LogicCell40 sTrigCounter_4_LC_8_9_1 (
            .in0(N__24230),
            .in1(N__24567),
            .in2(N__22812),
            .in3(N__22800),
            .lcout(sTrigCounterZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47813),
            .ce(),
            .sr(N__27540));
    defparam sTrigCounter_RNO_0_4_LC_8_9_2.C_ON=1'b0;
    defparam sTrigCounter_RNO_0_4_LC_8_9_2.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_0_4_LC_8_9_2.LUT_INIT=16'b0100110011001100;
    LogicCell40 sTrigCounter_RNO_0_4_LC_8_9_2 (
            .in0(N__24377),
            .in1(N__22809),
            .in2(N__24314),
            .in3(N__24699),
            .lcout(g1_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_2_5_LC_8_9_3.C_ON=1'b0;
    defparam sTrigCounter_RNO_2_5_LC_8_9_3.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_2_5_LC_8_9_3.LUT_INIT=16'b0100010011110000;
    LogicCell40 sTrigCounter_RNO_2_5_LC_8_9_3 (
            .in0(N__24823),
            .in1(N__22794),
            .in2(N__36878),
            .in3(N__36960),
            .lcout(),
            .ltout(g2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_5_LC_8_9_4.C_ON=1'b0;
    defparam sTrigCounter_5_LC_8_9_4.SEQ_MODE=4'b1000;
    defparam sTrigCounter_5_LC_8_9_4.LUT_INIT=16'b1010101010100110;
    LogicCell40 sTrigCounter_5_LC_8_9_4 (
            .in0(N__24651),
            .in1(N__22782),
            .in2(N__22776),
            .in3(N__24390),
            .lcout(sTrigCounterZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47813),
            .ce(),
            .sr(N__27540));
    defparam un4_speriod_cry_0_c_inv_LC_8_10_0.C_ON=1'b1;
    defparam un4_speriod_cry_0_c_inv_LC_8_10_0.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_0_c_inv_LC_8_10_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_0_c_inv_LC_8_10_0 (
            .in0(_gnd_net_),
            .in1(N__34230),
            .in2(N__22767),
            .in3(N__22773),
            .lcout(sEEPeriod_i_0),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(un4_speriod_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_1_c_inv_LC_8_10_1.C_ON=1'b1;
    defparam un4_speriod_cry_1_c_inv_LC_8_10_1.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_1_c_inv_LC_8_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_1_c_inv_LC_8_10_1 (
            .in0(_gnd_net_),
            .in1(N__35058),
            .in2(N__22752),
            .in3(N__22758),
            .lcout(sEEPeriod_i_1),
            .ltout(),
            .carryin(un4_speriod_cry_0),
            .carryout(un4_speriod_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_2_c_inv_LC_8_10_2.C_ON=1'b1;
    defparam un4_speriod_cry_2_c_inv_LC_8_10_2.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_2_c_inv_LC_8_10_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_2_c_inv_LC_8_10_2 (
            .in0(_gnd_net_),
            .in1(N__34957),
            .in2(N__22737),
            .in3(N__22743),
            .lcout(sEEPeriod_i_2),
            .ltout(),
            .carryin(un4_speriod_cry_1),
            .carryout(un4_speriod_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_3_c_inv_LC_8_10_3.C_ON=1'b1;
    defparam un4_speriod_cry_3_c_inv_LC_8_10_3.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_3_c_inv_LC_8_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_3_c_inv_LC_8_10_3 (
            .in0(_gnd_net_),
            .in1(N__34852),
            .in2(N__22722),
            .in3(N__22728),
            .lcout(sEEPeriod_i_3),
            .ltout(),
            .carryin(un4_speriod_cry_2),
            .carryout(un4_speriod_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_4_c_inv_LC_8_10_4.C_ON=1'b1;
    defparam un4_speriod_cry_4_c_inv_LC_8_10_4.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_4_c_inv_LC_8_10_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_4_c_inv_LC_8_10_4 (
            .in0(_gnd_net_),
            .in1(N__36855),
            .in2(N__22902),
            .in3(N__22908),
            .lcout(sEEPeriod_i_4),
            .ltout(),
            .carryin(un4_speriod_cry_3),
            .carryout(un4_speriod_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_5_c_inv_LC_8_10_5.C_ON=1'b1;
    defparam un4_speriod_cry_5_c_inv_LC_8_10_5.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_5_c_inv_LC_8_10_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_5_c_inv_LC_8_10_5 (
            .in0(_gnd_net_),
            .in1(N__34710),
            .in2(N__22887),
            .in3(N__22893),
            .lcout(sEEPeriod_i_5),
            .ltout(),
            .carryin(un4_speriod_cry_4),
            .carryout(un4_speriod_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_6_c_inv_LC_8_10_6.C_ON=1'b1;
    defparam un4_speriod_cry_6_c_inv_LC_8_10_6.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_6_c_inv_LC_8_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_6_c_inv_LC_8_10_6 (
            .in0(_gnd_net_),
            .in1(N__34605),
            .in2(N__22872),
            .in3(N__22878),
            .lcout(sEEPeriod_i_6),
            .ltout(),
            .carryin(un4_speriod_cry_5),
            .carryout(un4_speriod_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_7_c_inv_LC_8_10_7.C_ON=1'b1;
    defparam un4_speriod_cry_7_c_inv_LC_8_10_7.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_7_c_inv_LC_8_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_7_c_inv_LC_8_10_7 (
            .in0(_gnd_net_),
            .in1(N__34479),
            .in2(N__22857),
            .in3(N__22863),
            .lcout(sEEPeriod_i_7),
            .ltout(),
            .carryin(un4_speriod_cry_6),
            .carryout(un4_speriod_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_8_c_inv_LC_8_11_0.C_ON=1'b1;
    defparam un4_speriod_cry_8_c_inv_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_8_c_inv_LC_8_11_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_8_c_inv_LC_8_11_0 (
            .in0(_gnd_net_),
            .in1(N__35877),
            .in2(N__22848),
            .in3(N__24999),
            .lcout(sEEPeriod_i_8),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(un4_speriod_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_9_c_inv_LC_8_11_1.C_ON=1'b1;
    defparam un4_speriod_cry_9_c_inv_LC_8_11_1.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_9_c_inv_LC_8_11_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_9_c_inv_LC_8_11_1 (
            .in0(_gnd_net_),
            .in1(N__35762),
            .in2(N__22839),
            .in3(N__24993),
            .lcout(sEEPeriod_i_9),
            .ltout(),
            .carryin(un4_speriod_cry_8),
            .carryout(un4_speriod_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_10_c_inv_LC_8_11_2.C_ON=1'b1;
    defparam un4_speriod_cry_10_c_inv_LC_8_11_2.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_10_c_inv_LC_8_11_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_10_c_inv_LC_8_11_2 (
            .in0(_gnd_net_),
            .in1(N__35647),
            .in2(N__22830),
            .in3(N__24561),
            .lcout(sEEPeriod_i_10),
            .ltout(),
            .carryin(un4_speriod_cry_9),
            .carryout(un4_speriod_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_11_c_inv_LC_8_11_3.C_ON=1'b1;
    defparam un4_speriod_cry_11_c_inv_LC_8_11_3.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_11_c_inv_LC_8_11_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_11_c_inv_LC_8_11_3 (
            .in0(_gnd_net_),
            .in1(N__35532),
            .in2(N__22821),
            .in3(N__24555),
            .lcout(sEEPeriod_i_11),
            .ltout(),
            .carryin(un4_speriod_cry_10),
            .carryout(un4_speriod_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_12_c_inv_LC_8_11_4.C_ON=1'b1;
    defparam un4_speriod_cry_12_c_inv_LC_8_11_4.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_12_c_inv_LC_8_11_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_12_c_inv_LC_8_11_4 (
            .in0(_gnd_net_),
            .in1(N__35410),
            .in2(N__23004),
            .in3(N__24549),
            .lcout(sEEPeriod_i_12),
            .ltout(),
            .carryin(un4_speriod_cry_11),
            .carryout(un4_speriod_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_13_c_inv_LC_8_11_5.C_ON=1'b1;
    defparam un4_speriod_cry_13_c_inv_LC_8_11_5.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_13_c_inv_LC_8_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_13_c_inv_LC_8_11_5 (
            .in0(_gnd_net_),
            .in1(N__35306),
            .in2(N__22995),
            .in3(N__24543),
            .lcout(sEEPeriod_i_13),
            .ltout(),
            .carryin(un4_speriod_cry_12),
            .carryout(un4_speriod_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_14_c_inv_LC_8_11_6.C_ON=1'b1;
    defparam un4_speriod_cry_14_c_inv_LC_8_11_6.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_14_c_inv_LC_8_11_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_14_c_inv_LC_8_11_6 (
            .in0(_gnd_net_),
            .in1(N__35195),
            .in2(N__22986),
            .in3(N__25011),
            .lcout(sEEPeriod_i_14),
            .ltout(),
            .carryin(un4_speriod_cry_13),
            .carryout(un4_speriod_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_15_c_inv_LC_8_11_7.C_ON=1'b1;
    defparam un4_speriod_cry_15_c_inv_LC_8_11_7.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_15_c_inv_LC_8_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_15_c_inv_LC_8_11_7 (
            .in0(_gnd_net_),
            .in1(N__36637),
            .in2(N__22977),
            .in3(N__25005),
            .lcout(sEEPeriod_i_15),
            .ltout(),
            .carryin(un4_speriod_cry_14),
            .carryout(un4_speriod_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_16_c_inv_LC_8_12_0.C_ON=1'b1;
    defparam un4_speriod_cry_16_c_inv_LC_8_12_0.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_16_c_inv_LC_8_12_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_16_c_inv_LC_8_12_0 (
            .in0(_gnd_net_),
            .in1(N__36531),
            .in2(N__22962),
            .in3(N__22968),
            .lcout(sEEPeriod_i_16),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(un4_speriod_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_17_c_inv_LC_8_12_1.C_ON=1'b1;
    defparam un4_speriod_cry_17_c_inv_LC_8_12_1.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_17_c_inv_LC_8_12_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_17_c_inv_LC_8_12_1 (
            .in0(_gnd_net_),
            .in1(N__36426),
            .in2(N__22947),
            .in3(N__22953),
            .lcout(sEEPeriod_i_17),
            .ltout(),
            .carryin(un4_speriod_cry_16),
            .carryout(un4_speriod_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_18_c_inv_LC_8_12_2.C_ON=1'b1;
    defparam un4_speriod_cry_18_c_inv_LC_8_12_2.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_18_c_inv_LC_8_12_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_18_c_inv_LC_8_12_2 (
            .in0(_gnd_net_),
            .in1(N__36345),
            .in2(N__22932),
            .in3(N__22938),
            .lcout(sEEPeriod_i_18),
            .ltout(),
            .carryin(un4_speriod_cry_17),
            .carryout(un4_speriod_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_19_c_inv_LC_8_12_3.C_ON=1'b1;
    defparam un4_speriod_cry_19_c_inv_LC_8_12_3.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_19_c_inv_LC_8_12_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_19_c_inv_LC_8_12_3 (
            .in0(_gnd_net_),
            .in1(N__36252),
            .in2(N__22917),
            .in3(N__22923),
            .lcout(sEEPeriod_i_19),
            .ltout(),
            .carryin(un4_speriod_cry_18),
            .carryout(un4_speriod_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_20_c_inv_LC_8_12_4.C_ON=1'b1;
    defparam un4_speriod_cry_20_c_inv_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_20_c_inv_LC_8_12_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_20_c_inv_LC_8_12_4 (
            .in0(_gnd_net_),
            .in1(N__36162),
            .in2(N__23082),
            .in3(N__23088),
            .lcout(sEEPeriod_i_20),
            .ltout(),
            .carryin(un4_speriod_cry_19),
            .carryout(un4_speriod_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_21_c_inv_LC_8_12_5.C_ON=1'b1;
    defparam un4_speriod_cry_21_c_inv_LC_8_12_5.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_21_c_inv_LC_8_12_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_21_c_inv_LC_8_12_5 (
            .in0(_gnd_net_),
            .in1(N__23067),
            .in2(N__36080),
            .in3(N__23073),
            .lcout(sEEPeriod_i_21),
            .ltout(),
            .carryin(un4_speriod_cry_20),
            .carryout(un4_speriod_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_22_c_inv_LC_8_12_6.C_ON=1'b1;
    defparam un4_speriod_cry_22_c_inv_LC_8_12_6.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_22_c_inv_LC_8_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_22_c_inv_LC_8_12_6 (
            .in0(_gnd_net_),
            .in1(N__23055),
            .in2(N__35995),
            .in3(N__23061),
            .lcout(sEEPeriod_i_22),
            .ltout(),
            .carryin(un4_speriod_cry_21),
            .carryout(un4_speriod_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_23_c_inv_LC_8_12_7.C_ON=1'b1;
    defparam un4_speriod_cry_23_c_inv_LC_8_12_7.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_23_c_inv_LC_8_12_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_speriod_cry_23_c_inv_LC_8_12_7 (
            .in0(_gnd_net_),
            .in1(N__37074),
            .in2(N__23043),
            .in3(N__23049),
            .lcout(sEEPeriod_i_23),
            .ltout(),
            .carryin(un4_speriod_cry_22),
            .carryout(un4_speriod_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_23_THRU_LUT4_0_LC_8_13_0.C_ON=1'b0;
    defparam un4_speriod_cry_23_THRU_LUT4_0_LC_8_13_0.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_23_THRU_LUT4_0_LC_8_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un4_speriod_cry_23_THRU_LUT4_0_LC_8_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23034),
            .lcout(un4_speriod_cry_23_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNI3GS21_22_LC_8_13_3.C_ON=1'b0;
    defparam sCounter_RNI3GS21_22_LC_8_13_3.SEQ_MODE=4'b0000;
    defparam sCounter_RNI3GS21_22_LC_8_13_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNI3GS21_22_LC_8_13_3 (
            .in0(N__34929),
            .in1(N__34201),
            .in2(N__35979),
            .in3(N__35024),
            .lcout(un1_reset_rpi_inv_2_i_o3_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNI5HE71_8_LC_8_13_4.C_ON=1'b0;
    defparam sCounter_RNI5HE71_8_LC_8_13_4.SEQ_MODE=4'b0000;
    defparam sCounter_RNI5HE71_8_LC_8_13_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNI5HE71_8_LC_8_13_4 (
            .in0(N__35857),
            .in1(N__34695),
            .in2(N__35761),
            .in3(N__34827),
            .lcout(un1_reset_rpi_inv_2_i_o3_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_0_LC_8_13_7.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_0_LC_8_13_7.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_0_LC_8_13_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_0_LC_8_13_7 (
            .in0(N__23415),
            .in1(N__23436),
            .in2(N__23397),
            .in3(N__23454),
            .lcout(sbuttonModeStatus_0_sqmuxa_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_0_LC_8_14_0.C_ON=1'b1;
    defparam sCounter_0_LC_8_14_0.SEQ_MODE=4'b1010;
    defparam sCounter_0_LC_8_14_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_0_LC_8_14_0 (
            .in0(N__23244),
            .in1(N__34207),
            .in2(_gnd_net_),
            .in3(N__23007),
            .lcout(un7_spon_0),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(sCounter_cry_0),
            .clk(N__47822),
            .ce(),
            .sr(N__53016));
    defparam sCounter_1_LC_8_14_1.C_ON=1'b1;
    defparam sCounter_1_LC_8_14_1.SEQ_MODE=4'b1010;
    defparam sCounter_1_LC_8_14_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_1_LC_8_14_1 (
            .in0(N__23223),
            .in1(N__35034),
            .in2(_gnd_net_),
            .in3(N__23115),
            .lcout(un7_spon_1),
            .ltout(),
            .carryin(sCounter_cry_0),
            .carryout(sCounter_cry_1),
            .clk(N__47822),
            .ce(),
            .sr(N__53016));
    defparam sCounter_2_LC_8_14_2.C_ON=1'b1;
    defparam sCounter_2_LC_8_14_2.SEQ_MODE=4'b1010;
    defparam sCounter_2_LC_8_14_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_2_LC_8_14_2 (
            .in0(N__23245),
            .in1(N__34941),
            .in2(_gnd_net_),
            .in3(N__23112),
            .lcout(un7_spon_2),
            .ltout(),
            .carryin(sCounter_cry_1),
            .carryout(sCounter_cry_2),
            .clk(N__47822),
            .ce(),
            .sr(N__53016));
    defparam sCounter_3_LC_8_14_3.C_ON=1'b1;
    defparam sCounter_3_LC_8_14_3.SEQ_MODE=4'b1010;
    defparam sCounter_3_LC_8_14_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_3_LC_8_14_3 (
            .in0(N__23224),
            .in1(N__34833),
            .in2(_gnd_net_),
            .in3(N__23109),
            .lcout(un7_spon_3),
            .ltout(),
            .carryin(sCounter_cry_2),
            .carryout(sCounter_cry_3),
            .clk(N__47822),
            .ce(),
            .sr(N__53016));
    defparam sCounter_4_LC_8_14_4.C_ON=1'b1;
    defparam sCounter_4_LC_8_14_4.SEQ_MODE=4'b1010;
    defparam sCounter_4_LC_8_14_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_4_LC_8_14_4 (
            .in0(N__23246),
            .in1(N__36804),
            .in2(_gnd_net_),
            .in3(N__23106),
            .lcout(un7_spon_4),
            .ltout(),
            .carryin(sCounter_cry_3),
            .carryout(sCounter_cry_4),
            .clk(N__47822),
            .ce(),
            .sr(N__53016));
    defparam sCounter_5_LC_8_14_5.C_ON=1'b1;
    defparam sCounter_5_LC_8_14_5.SEQ_MODE=4'b1010;
    defparam sCounter_5_LC_8_14_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_5_LC_8_14_5 (
            .in0(N__23225),
            .in1(N__34699),
            .in2(_gnd_net_),
            .in3(N__23103),
            .lcout(un7_spon_5),
            .ltout(),
            .carryin(sCounter_cry_4),
            .carryout(sCounter_cry_5),
            .clk(N__47822),
            .ce(),
            .sr(N__53016));
    defparam sCounter_6_LC_8_14_6.C_ON=1'b1;
    defparam sCounter_6_LC_8_14_6.SEQ_MODE=4'b1010;
    defparam sCounter_6_LC_8_14_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_6_LC_8_14_6 (
            .in0(N__23247),
            .in1(N__34575),
            .in2(_gnd_net_),
            .in3(N__23100),
            .lcout(un7_spon_6),
            .ltout(),
            .carryin(sCounter_cry_5),
            .carryout(sCounter_cry_6),
            .clk(N__47822),
            .ce(),
            .sr(N__53016));
    defparam sCounter_7_LC_8_14_7.C_ON=1'b1;
    defparam sCounter_7_LC_8_14_7.SEQ_MODE=4'b1010;
    defparam sCounter_7_LC_8_14_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_7_LC_8_14_7 (
            .in0(N__23226),
            .in1(N__34453),
            .in2(_gnd_net_),
            .in3(N__23097),
            .lcout(un7_spon_7),
            .ltout(),
            .carryin(sCounter_cry_6),
            .carryout(sCounter_cry_7),
            .clk(N__47822),
            .ce(),
            .sr(N__53016));
    defparam sCounter_8_LC_8_15_0.C_ON=1'b1;
    defparam sCounter_8_LC_8_15_0.SEQ_MODE=4'b1010;
    defparam sCounter_8_LC_8_15_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_8_LC_8_15_0 (
            .in0(N__23218),
            .in1(N__35850),
            .in2(_gnd_net_),
            .in3(N__23094),
            .lcout(un7_spon_8),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(sCounter_cry_8),
            .clk(N__47831),
            .ce(),
            .sr(N__53008));
    defparam sCounter_9_LC_8_15_1.C_ON=1'b1;
    defparam sCounter_9_LC_8_15_1.SEQ_MODE=4'b1010;
    defparam sCounter_9_LC_8_15_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_9_LC_8_15_1 (
            .in0(N__23230),
            .in1(N__35739),
            .in2(_gnd_net_),
            .in3(N__23091),
            .lcout(un7_spon_9),
            .ltout(),
            .carryin(sCounter_cry_8),
            .carryout(sCounter_cry_9),
            .clk(N__47831),
            .ce(),
            .sr(N__53008));
    defparam sCounter_10_LC_8_15_2.C_ON=1'b1;
    defparam sCounter_10_LC_8_15_2.SEQ_MODE=4'b1010;
    defparam sCounter_10_LC_8_15_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_10_LC_8_15_2 (
            .in0(N__23215),
            .in1(N__35627),
            .in2(_gnd_net_),
            .in3(N__23142),
            .lcout(un7_spon_10),
            .ltout(),
            .carryin(sCounter_cry_9),
            .carryout(sCounter_cry_10),
            .clk(N__47831),
            .ce(),
            .sr(N__53008));
    defparam sCounter_11_LC_8_15_3.C_ON=1'b1;
    defparam sCounter_11_LC_8_15_3.SEQ_MODE=4'b1010;
    defparam sCounter_11_LC_8_15_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_11_LC_8_15_3 (
            .in0(N__23227),
            .in1(N__35516),
            .in2(_gnd_net_),
            .in3(N__23139),
            .lcout(un7_spon_11),
            .ltout(),
            .carryin(sCounter_cry_10),
            .carryout(sCounter_cry_11),
            .clk(N__47831),
            .ce(),
            .sr(N__53008));
    defparam sCounter_12_LC_8_15_4.C_ON=1'b1;
    defparam sCounter_12_LC_8_15_4.SEQ_MODE=4'b1010;
    defparam sCounter_12_LC_8_15_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_12_LC_8_15_4 (
            .in0(N__23216),
            .in1(N__35379),
            .in2(_gnd_net_),
            .in3(N__23136),
            .lcout(un7_spon_12),
            .ltout(),
            .carryin(sCounter_cry_11),
            .carryout(sCounter_cry_12),
            .clk(N__47831),
            .ce(),
            .sr(N__53008));
    defparam sCounter_13_LC_8_15_5.C_ON=1'b1;
    defparam sCounter_13_LC_8_15_5.SEQ_MODE=4'b1010;
    defparam sCounter_13_LC_8_15_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_13_LC_8_15_5 (
            .in0(N__23228),
            .in1(N__35291),
            .in2(_gnd_net_),
            .in3(N__23133),
            .lcout(un7_spon_13),
            .ltout(),
            .carryin(sCounter_cry_12),
            .carryout(sCounter_cry_13),
            .clk(N__47831),
            .ce(),
            .sr(N__53008));
    defparam sCounter_14_LC_8_15_6.C_ON=1'b1;
    defparam sCounter_14_LC_8_15_6.SEQ_MODE=4'b1010;
    defparam sCounter_14_LC_8_15_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_14_LC_8_15_6 (
            .in0(N__23217),
            .in1(N__35164),
            .in2(_gnd_net_),
            .in3(N__23130),
            .lcout(un7_spon_14),
            .ltout(),
            .carryin(sCounter_cry_13),
            .carryout(sCounter_cry_14),
            .clk(N__47831),
            .ce(),
            .sr(N__53008));
    defparam sCounter_15_LC_8_15_7.C_ON=1'b1;
    defparam sCounter_15_LC_8_15_7.SEQ_MODE=4'b1010;
    defparam sCounter_15_LC_8_15_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_15_LC_8_15_7 (
            .in0(N__23229),
            .in1(N__36633),
            .in2(_gnd_net_),
            .in3(N__23127),
            .lcout(un7_spon_15),
            .ltout(),
            .carryin(sCounter_cry_14),
            .carryout(sCounter_cry_15),
            .clk(N__47831),
            .ce(),
            .sr(N__53008));
    defparam sCounter_16_LC_8_16_0.C_ON=1'b1;
    defparam sCounter_16_LC_8_16_0.SEQ_MODE=4'b1010;
    defparam sCounter_16_LC_8_16_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_16_LC_8_16_0 (
            .in0(N__23240),
            .in1(N__36521),
            .in2(_gnd_net_),
            .in3(N__23124),
            .lcout(un7_spon_16),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(sCounter_cry_16),
            .clk(N__47838),
            .ce(),
            .sr(N__53000));
    defparam sCounter_17_LC_8_16_1.C_ON=1'b1;
    defparam sCounter_17_LC_8_16_1.SEQ_MODE=4'b1010;
    defparam sCounter_17_LC_8_16_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_17_LC_8_16_1 (
            .in0(N__23219),
            .in1(N__36405),
            .in2(_gnd_net_),
            .in3(N__23121),
            .lcout(un7_spon_17),
            .ltout(),
            .carryin(sCounter_cry_16),
            .carryout(sCounter_cry_17),
            .clk(N__47838),
            .ce(),
            .sr(N__53000));
    defparam sCounter_18_LC_8_16_2.C_ON=1'b1;
    defparam sCounter_18_LC_8_16_2.SEQ_MODE=4'b1010;
    defparam sCounter_18_LC_8_16_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_18_LC_8_16_2 (
            .in0(N__23241),
            .in1(N__36327),
            .in2(_gnd_net_),
            .in3(N__23118),
            .lcout(un7_spon_18),
            .ltout(),
            .carryin(sCounter_cry_17),
            .carryout(sCounter_cry_18),
            .clk(N__47838),
            .ce(),
            .sr(N__53000));
    defparam sCounter_19_LC_8_16_3.C_ON=1'b1;
    defparam sCounter_19_LC_8_16_3.SEQ_MODE=4'b1010;
    defparam sCounter_19_LC_8_16_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_19_LC_8_16_3 (
            .in0(N__23220),
            .in1(N__36229),
            .in2(_gnd_net_),
            .in3(N__23259),
            .lcout(un7_spon_19),
            .ltout(),
            .carryin(sCounter_cry_18),
            .carryout(sCounter_cry_19),
            .clk(N__47838),
            .ce(),
            .sr(N__53000));
    defparam sCounter_20_LC_8_16_4.C_ON=1'b1;
    defparam sCounter_20_LC_8_16_4.SEQ_MODE=4'b1010;
    defparam sCounter_20_LC_8_16_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_20_LC_8_16_4 (
            .in0(N__23242),
            .in1(N__36136),
            .in2(_gnd_net_),
            .in3(N__23256),
            .lcout(un7_spon_20),
            .ltout(),
            .carryin(sCounter_cry_19),
            .carryout(sCounter_cry_20),
            .clk(N__47838),
            .ce(),
            .sr(N__53000));
    defparam sCounter_21_LC_8_16_5.C_ON=1'b1;
    defparam sCounter_21_LC_8_16_5.SEQ_MODE=4'b1010;
    defparam sCounter_21_LC_8_16_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_21_LC_8_16_5 (
            .in0(N__23221),
            .in1(N__36064),
            .in2(_gnd_net_),
            .in3(N__23253),
            .lcout(un7_spon_21),
            .ltout(),
            .carryin(sCounter_cry_20),
            .carryout(sCounter_cry_21),
            .clk(N__47838),
            .ce(),
            .sr(N__53000));
    defparam sCounter_22_LC_8_16_6.C_ON=1'b1;
    defparam sCounter_22_LC_8_16_6.SEQ_MODE=4'b1010;
    defparam sCounter_22_LC_8_16_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_22_LC_8_16_6 (
            .in0(N__23243),
            .in1(N__35950),
            .in2(_gnd_net_),
            .in3(N__23250),
            .lcout(un7_spon_22),
            .ltout(),
            .carryin(sCounter_cry_21),
            .carryout(sCounter_cry_22),
            .clk(N__47838),
            .ce(),
            .sr(N__53000));
    defparam sCounter_23_LC_8_16_7.C_ON=1'b0;
    defparam sCounter_23_LC_8_16_7.SEQ_MODE=4'b1010;
    defparam sCounter_23_LC_8_16_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounter_23_LC_8_16_7 (
            .in0(N__23222),
            .in1(N__37053),
            .in2(_gnd_net_),
            .in3(N__23154),
            .lcout(un7_spon_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47838),
            .ce(),
            .sr(N__53000));
    defparam sbuttonModeStatus_RNO_3_LC_8_17_0.C_ON=1'b1;
    defparam sbuttonModeStatus_RNO_3_LC_8_17_0.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_3_LC_8_17_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 sbuttonModeStatus_RNO_3_LC_8_17_0 (
            .in0(_gnd_net_),
            .in1(N__26274),
            .in2(N__26313),
            .in3(N__32500),
            .lcout(sbuttonModeStatus_0_sqmuxa_0),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(un1_button_debounce_counter_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam button_debounce_counter_2_LC_8_17_1.C_ON=1'b1;
    defparam button_debounce_counter_2_LC_8_17_1.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_2_LC_8_17_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_2_LC_8_17_1 (
            .in0(N__32496),
            .in1(N__25197),
            .in2(_gnd_net_),
            .in3(N__23151),
            .lcout(button_debounce_counterZ0Z_2),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_1),
            .carryout(un1_button_debounce_counter_cry_2),
            .clk(N__53280),
            .ce(),
            .sr(N__26240));
    defparam button_debounce_counter_3_LC_8_17_2.C_ON=1'b1;
    defparam button_debounce_counter_3_LC_8_17_2.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_3_LC_8_17_2.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_3_LC_8_17_2 (
            .in0(N__32634),
            .in1(N__25224),
            .in2(_gnd_net_),
            .in3(N__23148),
            .lcout(button_debounce_counterZ0Z_3),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_2),
            .carryout(un1_button_debounce_counter_cry_3),
            .clk(N__53280),
            .ce(),
            .sr(N__26240));
    defparam button_debounce_counter_4_LC_8_17_3.C_ON=1'b1;
    defparam button_debounce_counter_4_LC_8_17_3.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_4_LC_8_17_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_4_LC_8_17_3 (
            .in0(N__32497),
            .in1(N__25236),
            .in2(_gnd_net_),
            .in3(N__23145),
            .lcout(button_debounce_counterZ0Z_4),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_3),
            .carryout(un1_button_debounce_counter_cry_4),
            .clk(N__53280),
            .ce(),
            .sr(N__26240));
    defparam button_debounce_counter_5_LC_8_17_4.C_ON=1'b1;
    defparam button_debounce_counter_5_LC_8_17_4.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_5_LC_8_17_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_5_LC_8_17_4 (
            .in0(N__32635),
            .in1(N__25211),
            .in2(_gnd_net_),
            .in3(N__23370),
            .lcout(button_debounce_counterZ0Z_5),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_4),
            .carryout(un1_button_debounce_counter_cry_5),
            .clk(N__53280),
            .ce(),
            .sr(N__26240));
    defparam button_debounce_counter_6_LC_8_17_5.C_ON=1'b1;
    defparam button_debounce_counter_6_LC_8_17_5.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_6_LC_8_17_5.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_6_LC_8_17_5 (
            .in0(N__32498),
            .in1(N__23367),
            .in2(_gnd_net_),
            .in3(N__23355),
            .lcout(button_debounce_counterZ0Z_6),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_5),
            .carryout(un1_button_debounce_counter_cry_6),
            .clk(N__53280),
            .ce(),
            .sr(N__26240));
    defparam button_debounce_counter_7_LC_8_17_6.C_ON=1'b1;
    defparam button_debounce_counter_7_LC_8_17_6.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_7_LC_8_17_6.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_7_LC_8_17_6 (
            .in0(N__32636),
            .in1(N__23352),
            .in2(_gnd_net_),
            .in3(N__23340),
            .lcout(button_debounce_counterZ0Z_7),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_6),
            .carryout(un1_button_debounce_counter_cry_7),
            .clk(N__53280),
            .ce(),
            .sr(N__26240));
    defparam button_debounce_counter_8_LC_8_17_7.C_ON=1'b1;
    defparam button_debounce_counter_8_LC_8_17_7.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_8_LC_8_17_7.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_8_LC_8_17_7 (
            .in0(N__32499),
            .in1(N__23337),
            .in2(_gnd_net_),
            .in3(N__23325),
            .lcout(button_debounce_counterZ0Z_8),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_7),
            .carryout(un1_button_debounce_counter_cry_8),
            .clk(N__53280),
            .ce(),
            .sr(N__26240));
    defparam button_debounce_counter_9_LC_8_18_0.C_ON=1'b1;
    defparam button_debounce_counter_9_LC_8_18_0.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_9_LC_8_18_0.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_9_LC_8_18_0 (
            .in0(N__32684),
            .in1(N__23321),
            .in2(_gnd_net_),
            .in3(N__23307),
            .lcout(button_debounce_counterZ0Z_9),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(un1_button_debounce_counter_cry_9),
            .clk(N__53281),
            .ce(),
            .sr(N__26241));
    defparam button_debounce_counter_10_LC_8_18_1.C_ON=1'b1;
    defparam button_debounce_counter_10_LC_8_18_1.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_10_LC_8_18_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_10_LC_8_18_1 (
            .in0(N__32677),
            .in1(N__23304),
            .in2(_gnd_net_),
            .in3(N__23292),
            .lcout(button_debounce_counterZ0Z_10),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_9),
            .carryout(un1_button_debounce_counter_cry_10),
            .clk(N__53281),
            .ce(),
            .sr(N__26241));
    defparam button_debounce_counter_11_LC_8_18_2.C_ON=1'b1;
    defparam button_debounce_counter_11_LC_8_18_2.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_11_LC_8_18_2.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_11_LC_8_18_2 (
            .in0(N__32681),
            .in1(N__23289),
            .in2(_gnd_net_),
            .in3(N__23277),
            .lcout(button_debounce_counterZ0Z_11),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_10),
            .carryout(un1_button_debounce_counter_cry_11),
            .clk(N__53281),
            .ce(),
            .sr(N__26241));
    defparam button_debounce_counter_12_LC_8_18_3.C_ON=1'b1;
    defparam button_debounce_counter_12_LC_8_18_3.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_12_LC_8_18_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_12_LC_8_18_3 (
            .in0(N__32678),
            .in1(N__23274),
            .in2(_gnd_net_),
            .in3(N__23262),
            .lcout(button_debounce_counterZ0Z_12),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_11),
            .carryout(un1_button_debounce_counter_cry_12),
            .clk(N__53281),
            .ce(),
            .sr(N__26241));
    defparam button_debounce_counter_13_LC_8_18_4.C_ON=1'b1;
    defparam button_debounce_counter_13_LC_8_18_4.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_13_LC_8_18_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_13_LC_8_18_4 (
            .in0(N__32682),
            .in1(N__23516),
            .in2(_gnd_net_),
            .in3(N__23502),
            .lcout(button_debounce_counterZ0Z_13),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_12),
            .carryout(un1_button_debounce_counter_cry_13),
            .clk(N__53281),
            .ce(),
            .sr(N__26241));
    defparam button_debounce_counter_14_LC_8_18_5.C_ON=1'b1;
    defparam button_debounce_counter_14_LC_8_18_5.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_14_LC_8_18_5.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_14_LC_8_18_5 (
            .in0(N__32679),
            .in1(N__23499),
            .in2(_gnd_net_),
            .in3(N__23487),
            .lcout(button_debounce_counterZ0Z_14),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_13),
            .carryout(un1_button_debounce_counter_cry_14),
            .clk(N__53281),
            .ce(),
            .sr(N__26241));
    defparam button_debounce_counter_15_LC_8_18_6.C_ON=1'b1;
    defparam button_debounce_counter_15_LC_8_18_6.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_15_LC_8_18_6.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_15_LC_8_18_6 (
            .in0(N__32683),
            .in1(N__23484),
            .in2(_gnd_net_),
            .in3(N__23472),
            .lcout(button_debounce_counterZ0Z_15),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_14),
            .carryout(un1_button_debounce_counter_cry_15),
            .clk(N__53281),
            .ce(),
            .sr(N__26241));
    defparam button_debounce_counter_16_LC_8_18_7.C_ON=1'b1;
    defparam button_debounce_counter_16_LC_8_18_7.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_16_LC_8_18_7.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_16_LC_8_18_7 (
            .in0(N__32680),
            .in1(N__23469),
            .in2(_gnd_net_),
            .in3(N__23457),
            .lcout(button_debounce_counterZ0Z_16),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_15),
            .carryout(un1_button_debounce_counter_cry_16),
            .clk(N__53281),
            .ce(),
            .sr(N__26241));
    defparam button_debounce_counter_17_LC_8_19_0.C_ON=1'b1;
    defparam button_debounce_counter_17_LC_8_19_0.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_17_LC_8_19_0.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_17_LC_8_19_0 (
            .in0(N__32685),
            .in1(N__23450),
            .in2(_gnd_net_),
            .in3(N__23439),
            .lcout(button_debounce_counterZ0Z_17),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(un1_button_debounce_counter_cry_17),
            .clk(N__53282),
            .ce(),
            .sr(N__26242));
    defparam button_debounce_counter_18_LC_8_19_1.C_ON=1'b1;
    defparam button_debounce_counter_18_LC_8_19_1.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_18_LC_8_19_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_18_LC_8_19_1 (
            .in0(N__32688),
            .in1(N__23429),
            .in2(_gnd_net_),
            .in3(N__23418),
            .lcout(button_debounce_counterZ0Z_18),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_17),
            .carryout(un1_button_debounce_counter_cry_18),
            .clk(N__53282),
            .ce(),
            .sr(N__26242));
    defparam button_debounce_counter_19_LC_8_19_2.C_ON=1'b1;
    defparam button_debounce_counter_19_LC_8_19_2.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_19_LC_8_19_2.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_19_LC_8_19_2 (
            .in0(N__32686),
            .in1(N__23411),
            .in2(_gnd_net_),
            .in3(N__23400),
            .lcout(button_debounce_counterZ0Z_19),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_18),
            .carryout(un1_button_debounce_counter_cry_19),
            .clk(N__53282),
            .ce(),
            .sr(N__26242));
    defparam button_debounce_counter_20_LC_8_19_3.C_ON=1'b1;
    defparam button_debounce_counter_20_LC_8_19_3.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_20_LC_8_19_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_20_LC_8_19_3 (
            .in0(N__32689),
            .in1(N__23387),
            .in2(_gnd_net_),
            .in3(N__23376),
            .lcout(button_debounce_counterZ0Z_20),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_19),
            .carryout(un1_button_debounce_counter_cry_20),
            .clk(N__53282),
            .ce(),
            .sr(N__26242));
    defparam button_debounce_counter_21_LC_8_19_4.C_ON=1'b1;
    defparam button_debounce_counter_21_LC_8_19_4.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_21_LC_8_19_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_21_LC_8_19_4 (
            .in0(N__32687),
            .in1(N__25286),
            .in2(_gnd_net_),
            .in3(N__23373),
            .lcout(button_debounce_counterZ0Z_21),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_20),
            .carryout(un1_button_debounce_counter_cry_21),
            .clk(N__53282),
            .ce(),
            .sr(N__26242));
    defparam button_debounce_counter_22_LC_8_19_5.C_ON=1'b1;
    defparam button_debounce_counter_22_LC_8_19_5.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_22_LC_8_19_5.LUT_INIT=16'b0110011011001100;
    LogicCell40 button_debounce_counter_22_LC_8_19_5 (
            .in0(N__32690),
            .in1(N__25265),
            .in2(_gnd_net_),
            .in3(N__23553),
            .lcout(button_debounce_counterZ0Z_22),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_21),
            .carryout(un1_button_debounce_counter_cry_22),
            .clk(N__53282),
            .ce(),
            .sr(N__26242));
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_0_LC_8_19_6.C_ON=1'b1;
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_0_LC_8_19_6.SEQ_MODE=4'b0000;
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_0_LC_8_19_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_button_debounce_counter_cry_22_c_THRU_CRY_0_LC_8_19_6 (
            .in0(_gnd_net_),
            .in1(N__38020),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_22),
            .carryout(un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_1_LC_8_19_7.C_ON=1'b1;
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_1_LC_8_19_7.SEQ_MODE=4'b0000;
    defparam un1_button_debounce_counter_cry_22_c_THRU_CRY_1_LC_8_19_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_button_debounce_counter_cry_22_c_THRU_CRY_1_LC_8_19_7 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__38068),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_button_debounce_counter_cry_22_THRU_CRY_0_THRU_CO),
            .carryout(un1_button_debounce_counter_cry_22_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam button_debounce_counter_esr_23_LC_8_20_0.C_ON=1'b0;
    defparam button_debounce_counter_esr_23_LC_8_20_0.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_esr_23_LC_8_20_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 button_debounce_counter_esr_23_LC_8_20_0 (
            .in0(_gnd_net_),
            .in1(N__23543),
            .in2(_gnd_net_),
            .in3(N__23550),
            .lcout(button_debounce_counterZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53283),
            .ce(N__25470),
            .sr(N__26243));
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_c_LC_9_3_0 .C_ON=1'b1;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_c_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_c_LC_9_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_c_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(N__25552),
            .in2(N__25503),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_3_0_),
            .carryout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_LUT4_0_LC_9_3_1 .C_ON=1'b1;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_LUT4_0_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_LUT4_0_LC_9_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_LUT4_0_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(N__25574),
            .in2(_gnd_net_),
            .in3(N__23529),
            .lcout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_0 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_LUT4_0_LC_9_3_2 .C_ON=1'b1;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_LUT4_0_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_LUT4_0_LC_9_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_LUT4_0_LC_9_3_2  (
            .in0(_gnd_net_),
            .in1(N__25774),
            .in2(_gnd_net_),
            .in3(N__23526),
            .lcout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_1 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_3_LC_9_3_3 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_3_LC_9_3_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_3_LC_9_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_3_LC_9_3_3  (
            .in0(_gnd_net_),
            .in1(N__25590),
            .in2(_gnd_net_),
            .in3(N__23523),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_2 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3 ),
            .clk(N__30703),
            .ce(),
            .sr(N__53123));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_4_LC_9_3_4 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_4_LC_9_3_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_4_LC_9_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_4_LC_9_3_4  (
            .in0(_gnd_net_),
            .in1(N__25533),
            .in2(_gnd_net_),
            .in3(N__23520),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_3 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_pos_sclk_i_cry_4 ),
            .clk(N__30703),
            .ce(),
            .sr(N__53123));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_5_LC_9_3_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_5_LC_9_3_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_5_LC_9_3_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_5_LC_9_3_5  (
            .in0(_gnd_net_),
            .in1(N__25796),
            .in2(_gnd_net_),
            .in3(N__23607),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30703),
            .ce(),
            .sr(N__53123));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_1_LC_9_4_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_1_LC_9_4_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_1_LC_9_4_0 .LUT_INIT=16'b0010100000111100;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_1_LC_9_4_0  (
            .in0(N__33222),
            .in1(N__23604),
            .in2(N__25578),
            .in3(N__25517),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30705),
            .ce(),
            .sr(N__53108));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_2_LC_9_4_4 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_2_LC_9_4_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_2_LC_9_4_4 .LUT_INIT=16'b0000101110110000;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_2_LC_9_4_4  (
            .in0(N__33223),
            .in1(N__25518),
            .in2(N__25779),
            .in3(N__23598),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30705),
            .ce(),
            .sr(N__53108));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_0_LC_9_4_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_0_LC_9_4_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_0_LC_9_4_5 .LUT_INIT=16'b0011110000010100;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_0_LC_9_4_5  (
            .in0(N__25516),
            .in1(N__25502),
            .in2(N__25557),
            .in3(N__33221),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30705),
            .ce(),
            .sr(N__53108));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_12_LC_9_5_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_12_LC_9_5_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_12_LC_9_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_12_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25716),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53250),
            .ce(),
            .sr(N__53094));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_2_LC_9_5_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_2_LC_9_5_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_2_LC_9_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_2_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25728),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53250),
            .ce(),
            .sr(N__53094));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_3_LC_9_5_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_3_LC_9_5_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_3_LC_9_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_3_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25710),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53250),
            .ce(),
            .sr(N__53094));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_4_LC_9_5_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_4_LC_9_5_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_4_LC_9_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_4_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28737),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53250),
            .ce(),
            .sr(N__53094));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_5_LC_9_5_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_5_LC_9_5_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_5_LC_9_5_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_5_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__28728),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53250),
            .ce(),
            .sr(N__53094));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_15_LC_9_5_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_15_LC_9_5_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_15_LC_9_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_15_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25986),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53250),
            .ce(),
            .sr(N__53094));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_11_LC_9_5_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_11_LC_9_5_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_11_LC_9_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_11_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25722),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53250),
            .ce(),
            .sr(N__53094));
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_10_LC_9_5_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_10_LC_9_5_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.txdata_reg_i_10_LC_9_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.txdata_reg_i_10_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28761),
            .lcout(\spi_master_inst.spi_data_path_u1.txdata_reg_iZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53250),
            .ce(),
            .sr(N__53094));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNISEQE3_1_LC_9_6_0 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNISEQE3_1_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNISEQE3_1_LC_9_6_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNISEQE3_1_LC_9_6_0  (
            .in0(N__25964),
            .in1(N__24072),
            .in2(N__25947),
            .in3(N__23613),
            .lcout(\spi_master_inst.sclk_gen_u0.N_158_7 ),
            .ltout(\spi_master_inst.sclk_gen_u0.N_158_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNO_0_LC_9_6_1 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNO_0_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNO_0_LC_9_6_1 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNO_0_LC_9_6_1  (
            .in0(N__23735),
            .in1(N__26994),
            .in2(N__23697),
            .in3(N__23678),
            .lcout(\spi_master_inst.sclk_gen_u0.un1_delay_count_start_i_0_sqmuxa_2_0_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNIK09A_LC_9_6_2 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNIK09A_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNIK09A_LC_9_6_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \spi_master_inst.sclk_gen_u0.falling_count_start_i_RNIK09A_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__23641),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_master_inst.sclk_gen_u0.falling_count_start_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_ft_ibuf_RNI4OFN_1_LC_9_6_3.C_ON=1'b0;
    defparam trig_ft_ibuf_RNI4OFN_1_LC_9_6_3.SEQ_MODE=4'b0000;
    defparam trig_ft_ibuf_RNI4OFN_1_LC_9_6_3.LUT_INIT=16'b0000000000010001;
    LogicCell40 trig_ft_ibuf_RNI4OFN_1_LC_9_6_3 (
            .in0(N__24065),
            .in1(N__23978),
            .in2(_gnd_net_),
            .in3(N__23877),
            .lcout(un3_trig_0_0),
            .ltout(un3_trig_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_3_5_LC_9_6_4.C_ON=1'b0;
    defparam sTrigCounter_RNO_3_5_LC_9_6_4.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_3_5_LC_9_6_4.LUT_INIT=16'b1100100011111010;
    LogicCell40 sTrigCounter_RNO_3_5_LC_9_6_4 (
            .in0(N__24506),
            .in1(N__24941),
            .in2(N__23616),
            .in3(N__29093),
            .lcout(g1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNIKGMR_0_LC_9_6_5 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNIKGMR_0_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNIKGMR_0_LC_9_6_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNIKGMR_0_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(N__25913),
            .in2(_gnd_net_),
            .in3(N__25979),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNILEDN1_7_LC_9_6_6 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNILEDN1_7_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNILEDN1_7_LC_9_6_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_RNILEDN1_7_LC_9_6_6  (
            .in0(N__25898),
            .in1(N__25829),
            .in2(N__25884),
            .in3(N__25928),
            .lcout(\spi_master_inst.sclk_gen_u0.spim_clk_state_i_ns_i_a3_0_7_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_ft_ibuf_RNI4OFN_4_LC_9_6_7.C_ON=1'b0;
    defparam trig_ft_ibuf_RNI4OFN_4_LC_9_6_7.SEQ_MODE=4'b0000;
    defparam trig_ft_ibuf_RNI4OFN_4_LC_9_6_7.LUT_INIT=16'b0000000000010001;
    LogicCell40 trig_ft_ibuf_RNI4OFN_4_LC_9_6_7 (
            .in0(N__24066),
            .in1(N__23979),
            .in2(_gnd_net_),
            .in3(N__23878),
            .lcout(un3_trig_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNINQ4B1_2_LC_9_7_0.C_ON=1'b0;
    defparam sEETrigCounter_RNINQ4B1_2_LC_9_7_0.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNINQ4B1_2_LC_9_7_0.LUT_INIT=16'b0000000000000101;
    LogicCell40 sEETrigCounter_RNINQ4B1_2_LC_9_7_0 (
            .in0(N__26013),
            .in1(_gnd_net_),
            .in2(N__26082),
            .in3(N__26111),
            .lcout(),
            .ltout(un8_trig_prev_0_c5_a0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNII5M43_6_LC_9_7_1.C_ON=1'b0;
    defparam sEETrigCounter_RNII5M43_6_LC_9_7_1.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNII5M43_6_LC_9_7_1.LUT_INIT=16'b1100110001101100;
    LogicCell40 sEETrigCounter_RNII5M43_6_LC_9_7_1 (
            .in0(N__24163),
            .in1(N__23808),
            .in2(N__23826),
            .in3(N__23820),
            .lcout(un10_trig_prev_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIHO9M2_5_LC_9_7_2.C_ON=1'b0;
    defparam sEETrigCounter_RNIHO9M2_5_LC_9_7_2.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIHO9M2_5_LC_9_7_2.LUT_INIT=16'b1001101010101010;
    LogicCell40 sEETrigCounter_RNIHO9M2_5_LC_9_7_2 (
            .in0(N__23819),
            .in1(N__26116),
            .in2(N__24165),
            .in3(N__23789),
            .lcout(un10_trig_prev_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIPGOS_2_LC_9_7_3.C_ON=1'b0;
    defparam sEETrigCounter_RNIPGOS_2_LC_9_7_3.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIPGOS_2_LC_9_7_3.LUT_INIT=16'b0000000000110011;
    LogicCell40 sEETrigCounter_RNIPGOS_2_LC_9_7_3 (
            .in0(_gnd_net_),
            .in1(N__26012),
            .in2(_gnd_net_),
            .in3(N__26076),
            .lcout(un8_trig_prev_0_c4_a0_1),
            .ltout(un8_trig_prev_0_c4_a0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIHCT72_4_LC_9_7_4.C_ON=1'b0;
    defparam sEETrigCounter_RNIHCT72_4_LC_9_7_4.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIHCT72_4_LC_9_7_4.LUT_INIT=16'b1110111100010000;
    LogicCell40 sEETrigCounter_RNIHCT72_4_LC_9_7_4 (
            .in0(N__26036),
            .in1(N__26115),
            .in2(N__23823),
            .in3(N__24176),
            .lcout(un10_trig_prev_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIV25B1_6_LC_9_7_5.C_ON=1'b0;
    defparam sEETrigCounter_RNIV25B1_6_LC_9_7_5.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIV25B1_6_LC_9_7_5.LUT_INIT=16'b0000000000000011;
    LogicCell40 sEETrigCounter_RNIV25B1_6_LC_9_7_5 (
            .in0(_gnd_net_),
            .in1(N__23818),
            .in2(N__26120),
            .in3(N__23807),
            .lcout(),
            .ltout(un8_trig_prev_0_c7_a0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIKJ2J3_7_LC_9_7_6.C_ON=1'b0;
    defparam sEETrigCounter_RNIKJ2J3_7_LC_9_7_6.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIKJ2J3_7_LC_9_7_6.LUT_INIT=16'b0110101010101010;
    LogicCell40 sEETrigCounter_RNIKJ2J3_7_LC_9_7_6 (
            .in0(N__23799),
            .in1(N__24164),
            .in2(N__23793),
            .in3(N__23790),
            .lcout(un10_trig_prev_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIQHOS_4_LC_9_7_7.C_ON=1'b0;
    defparam sEETrigCounter_RNIQHOS_4_LC_9_7_7.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIQHOS_4_LC_9_7_7.LUT_INIT=16'b0000000000001111;
    LogicCell40 sEETrigCounter_RNIQHOS_4_LC_9_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24177),
            .in3(N__26035),
            .lcout(un8_trig_prev_0_c5_a0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_0_c_inv_LC_9_8_0.C_ON=1'b1;
    defparam un10_trig_prev_cry_0_c_inv_LC_9_8_0.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_0_c_inv_LC_9_8_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_0_c_inv_LC_9_8_0 (
            .in0(_gnd_net_),
            .in1(N__24147),
            .in2(N__26055),
            .in3(N__31379),
            .lcout(sTrigCounter_i_0),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(un10_trig_prev_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_1_c_inv_LC_9_8_1.C_ON=1'b1;
    defparam un10_trig_prev_cry_1_c_inv_LC_9_8_1.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_1_c_inv_LC_9_8_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_1_c_inv_LC_9_8_1 (
            .in0(_gnd_net_),
            .in1(N__24141),
            .in2(N__25995),
            .in3(N__31298),
            .lcout(sTrigCounter_i_1),
            .ltout(),
            .carryin(un10_trig_prev_cry_0),
            .carryout(un10_trig_prev_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_2_c_inv_LC_9_8_2.C_ON=1'b1;
    defparam un10_trig_prev_cry_2_c_inv_LC_9_8_2.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_2_c_inv_LC_9_8_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_2_c_inv_LC_9_8_2 (
            .in0(_gnd_net_),
            .in1(N__26061),
            .in2(N__24135),
            .in3(N__24612),
            .lcout(sTrigCounter_i_2),
            .ltout(),
            .carryin(un10_trig_prev_cry_1),
            .carryout(un10_trig_prev_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_3_c_inv_LC_9_8_3.C_ON=1'b1;
    defparam un10_trig_prev_cry_3_c_inv_LC_9_8_3.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_3_c_inv_LC_9_8_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 un10_trig_prev_cry_3_c_inv_LC_9_8_3 (
            .in0(N__24200),
            .in1(N__24126),
            .in2(N__26094),
            .in3(_gnd_net_),
            .lcout(sTrigCounter_i_3),
            .ltout(),
            .carryin(un10_trig_prev_cry_2),
            .carryout(un10_trig_prev_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_4_c_inv_LC_9_8_4.C_ON=1'b1;
    defparam un10_trig_prev_cry_4_c_inv_LC_9_8_4.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_4_c_inv_LC_9_8_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 un10_trig_prev_cry_4_c_inv_LC_9_8_4 (
            .in0(N__24231),
            .in1(N__24111),
            .in2(N__24120),
            .in3(_gnd_net_),
            .lcout(sTrigCounter_i_4),
            .ltout(),
            .carryin(un10_trig_prev_cry_3),
            .carryout(un10_trig_prev_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_5_c_inv_LC_9_8_5.C_ON=1'b1;
    defparam un10_trig_prev_cry_5_c_inv_LC_9_8_5.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_5_c_inv_LC_9_8_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_5_c_inv_LC_9_8_5 (
            .in0(_gnd_net_),
            .in1(N__24096),
            .in2(N__24105),
            .in3(N__24645),
            .lcout(sTrigCounter_i_5),
            .ltout(),
            .carryin(un10_trig_prev_cry_4),
            .carryout(un10_trig_prev_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_6_c_inv_LC_9_8_6.C_ON=1'b1;
    defparam un10_trig_prev_cry_6_c_inv_LC_9_8_6.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_6_c_inv_LC_9_8_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un10_trig_prev_cry_6_c_inv_LC_9_8_6 (
            .in0(N__25076),
            .in1(N__24081),
            .in2(N__24090),
            .in3(_gnd_net_),
            .lcout(sTrigCounter_i_6),
            .ltout(),
            .carryin(un10_trig_prev_cry_5),
            .carryout(un10_trig_prev_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_7_c_inv_LC_9_8_7.C_ON=1'b1;
    defparam un10_trig_prev_cry_7_c_inv_LC_9_8_7.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_7_c_inv_LC_9_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un10_trig_prev_cry_7_c_inv_LC_9_8_7 (
            .in0(_gnd_net_),
            .in1(N__24528),
            .in2(N__24537),
            .in3(N__25032),
            .lcout(sTrigCounter_i_7),
            .ltout(),
            .carryin(un10_trig_prev_cry_6),
            .carryout(un10_trig_prev_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un10_trig_prev_cry_7_THRU_LUT4_0_LC_9_9_0.C_ON=1'b0;
    defparam un10_trig_prev_cry_7_THRU_LUT4_0_LC_9_9_0.SEQ_MODE=4'b0000;
    defparam un10_trig_prev_cry_7_THRU_LUT4_0_LC_9_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un10_trig_prev_cry_7_THRU_LUT4_0_LC_9_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24522),
            .lcout(un10_trig_prev_cry_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_1_1_LC_9_9_1.C_ON=1'b0;
    defparam sAddress_RNI9IH12_1_1_LC_9_9_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_1_1_LC_9_9_1.LUT_INIT=16'b0000000100000000;
    LogicCell40 sAddress_RNI9IH12_1_1_LC_9_9_1 (
            .in0(N__46451),
            .in1(N__31106),
            .in2(N__44478),
            .in3(N__44745),
            .lcout(sAddress_RNI9IH12_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_3_2_LC_9_9_2.C_ON=1'b0;
    defparam sTrigCounter_RNO_3_2_LC_9_9_2.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_3_2_LC_9_9_2.LUT_INIT=16'b1100100011111010;
    LogicCell40 sTrigCounter_RNO_3_2_LC_9_9_2 (
            .in0(N__24510),
            .in1(N__24943),
            .in2(N__24428),
            .in3(N__29084),
            .lcout(g1_0_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_0_5_LC_9_9_3.C_ON=1'b0;
    defparam sTrigCounter_RNO_0_5_LC_9_9_3.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_0_5_LC_9_9_3.LUT_INIT=16'b0111111100000000;
    LogicCell40 sTrigCounter_RNO_0_5_LC_9_9_3 (
            .in0(N__24273),
            .in1(N__24378),
            .in2(N__24713),
            .in3(N__24399),
            .lcout(g1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_0_7_LC_9_9_4.C_ON=1'b0;
    defparam sTrigCounter_RNO_0_7_LC_9_9_4.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_0_7_LC_9_9_4.LUT_INIT=16'b0111000011110000;
    LogicCell40 sTrigCounter_RNO_0_7_LC_9_9_4 (
            .in0(N__24379),
            .in1(N__24272),
            .in2(N__27576),
            .in3(N__24694),
            .lcout(N_123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNI9UM4_4_LC_9_9_5.C_ON=1'b0;
    defparam sTrigCounter_RNI9UM4_4_LC_9_9_5.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNI9UM4_4_LC_9_9_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 sTrigCounter_RNI9UM4_4_LC_9_9_5 (
            .in0(_gnd_net_),
            .in1(N__24228),
            .in2(_gnd_net_),
            .in3(N__24201),
            .lcout(un1_sTrigCounter_ac0_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_4_4_LC_9_9_7.C_ON=1'b0;
    defparam sTrigCounter_RNO_4_4_LC_9_9_7.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_4_4_LC_9_9_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 sTrigCounter_RNO_4_4_LC_9_9_7 (
            .in0(N__32562),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24202),
            .lcout(g1_0_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_2_6_LC_9_10_0.C_ON=1'b0;
    defparam sTrigCounter_RNO_2_6_LC_9_10_0.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_2_6_LC_9_10_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 sTrigCounter_RNO_2_6_LC_9_10_0 (
            .in0(_gnd_net_),
            .in1(N__31293),
            .in2(_gnd_net_),
            .in3(N__31390),
            .lcout(),
            .ltout(un1_sTrigCounter_ac0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_1_6_LC_9_10_1.C_ON=1'b0;
    defparam sTrigCounter_RNO_1_6_LC_9_10_1.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_1_6_LC_9_10_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 sTrigCounter_RNO_1_6_LC_9_10_1 (
            .in0(N__24626),
            .in1(N__24646),
            .in2(N__24744),
            .in3(N__24613),
            .lcout(),
            .ltout(un1_sTrigCounter_ac0_0_2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_0_6_LC_9_10_2.C_ON=1'b0;
    defparam sTrigCounter_RNO_0_6_LC_9_10_2.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_0_6_LC_9_10_2.LUT_INIT=16'b0111000001010000;
    LogicCell40 sTrigCounter_RNO_0_6_LC_9_10_2 (
            .in0(N__27568),
            .in1(N__24741),
            .in2(N__24723),
            .in3(N__24698),
            .lcout(un1_sTrigCounter_ac0_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_2_7_LC_9_10_3.C_ON=1'b0;
    defparam sTrigCounter_RNO_2_7_LC_9_10_3.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_2_7_LC_9_10_3.LUT_INIT=16'b1010000000000000;
    LogicCell40 sTrigCounter_RNO_2_7_LC_9_10_3 (
            .in0(N__31391),
            .in1(_gnd_net_),
            .in2(N__31302),
            .in3(N__24614),
            .lcout(),
            .ltout(un1_sTrigCounter_ac0_3_out_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_1_7_LC_9_10_4.C_ON=1'b0;
    defparam sTrigCounter_RNO_1_7_LC_9_10_4.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_1_7_LC_9_10_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 sTrigCounter_RNO_1_7_LC_9_10_4 (
            .in0(N__24647),
            .in1(N__24627),
            .in2(N__24618),
            .in3(N__25077),
            .lcout(un1_sTrigCounter_axbxc7_m7_0_a2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_RNO_1_4_LC_9_10_6.C_ON=1'b0;
    defparam sTrigCounter_RNO_1_4_LC_9_10_6.SEQ_MODE=4'b0000;
    defparam sTrigCounter_RNO_1_4_LC_9_10_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 sTrigCounter_RNO_1_4_LC_9_10_6 (
            .in0(N__24615),
            .in1(N__31297),
            .in2(N__24576),
            .in3(N__31392),
            .lcout(g1_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPeriod_10_LC_9_11_0.C_ON=1'b0;
    defparam sEEPeriod_10_LC_9_11_0.SEQ_MODE=4'b1011;
    defparam sEEPeriod_10_LC_9_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_10_LC_9_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50281),
            .lcout(sEEPeriodZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47776),
            .ce(N__28944),
            .sr(N__53028));
    defparam sEEPeriod_11_LC_9_11_1.C_ON=1'b0;
    defparam sEEPeriod_11_LC_9_11_1.SEQ_MODE=4'b1010;
    defparam sEEPeriod_11_LC_9_11_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 sEEPeriod_11_LC_9_11_1 (
            .in0(_gnd_net_),
            .in1(N__49785),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47776),
            .ce(N__28944),
            .sr(N__53028));
    defparam sEEPeriod_12_LC_9_11_2.C_ON=1'b0;
    defparam sEEPeriod_12_LC_9_11_2.SEQ_MODE=4'b1010;
    defparam sEEPeriod_12_LC_9_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_12_LC_9_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49367),
            .lcout(sEEPeriodZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47776),
            .ce(N__28944),
            .sr(N__53028));
    defparam sEEPeriod_13_LC_9_11_3.C_ON=1'b0;
    defparam sEEPeriod_13_LC_9_11_3.SEQ_MODE=4'b1010;
    defparam sEEPeriod_13_LC_9_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_13_LC_9_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47062),
            .lcout(sEEPeriodZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47776),
            .ce(N__28944),
            .sr(N__53028));
    defparam sEEPeriod_14_LC_9_11_4.C_ON=1'b0;
    defparam sEEPeriod_14_LC_9_11_4.SEQ_MODE=4'b1010;
    defparam sEEPeriod_14_LC_9_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_14_LC_9_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48244),
            .lcout(sEEPeriodZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47776),
            .ce(N__28944),
            .sr(N__53028));
    defparam sEEPeriod_15_LC_9_11_5.C_ON=1'b0;
    defparam sEEPeriod_15_LC_9_11_5.SEQ_MODE=4'b1011;
    defparam sEEPeriod_15_LC_9_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_15_LC_9_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48633),
            .lcout(sEEPeriodZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47776),
            .ce(N__28944),
            .sr(N__53028));
    defparam sEEPeriod_8_LC_9_11_6.C_ON=1'b0;
    defparam sEEPeriod_8_LC_9_11_6.SEQ_MODE=4'b1010;
    defparam sEEPeriod_8_LC_9_11_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPeriod_8_LC_9_11_6 (
            .in0(N__51139),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPeriodZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47776),
            .ce(N__28944),
            .sr(N__53028));
    defparam sEEPeriod_9_LC_9_11_7.C_ON=1'b0;
    defparam sEEPeriod_9_LC_9_11_7.SEQ_MODE=4'b1011;
    defparam sEEPeriod_9_LC_9_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPeriod_9_LC_9_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50665),
            .lcout(sEEPeriodZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47776),
            .ce(N__28944),
            .sr(N__53028));
    defparam sCounter_RNIM34L_0_10_LC_9_12_0.C_ON=1'b0;
    defparam sCounter_RNIM34L_0_10_LC_9_12_0.SEQ_MODE=4'b0000;
    defparam sCounter_RNIM34L_0_10_LC_9_12_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNIM34L_0_10_LC_9_12_0 (
            .in0(N__35522),
            .in1(N__35298),
            .in2(N__35396),
            .in3(N__35632),
            .lcout(op_gt_op_gt_un13_striginternallto23_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIM34L_10_LC_9_12_1.C_ON=1'b0;
    defparam sCounter_RNIM34L_10_LC_9_12_1.SEQ_MODE=4'b0000;
    defparam sCounter_RNIM34L_10_LC_9_12_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounter_RNIM34L_10_LC_9_12_1 (
            .in0(N__35631),
            .in1(N__35380),
            .in2(N__35310),
            .in3(N__35521),
            .lcout(un1_reset_rpi_inv_2_i_o3_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIO6BU_23_LC_9_12_2.C_ON=1'b0;
    defparam sCounter_RNIO6BU_23_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam sCounter_RNIO6BU_23_LC_9_12_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 sCounter_RNIO6BU_23_LC_9_12_2 (
            .in0(N__35981),
            .in1(N__34949),
            .in2(N__37089),
            .in3(N__35050),
            .lcout(op_gt_op_gt_un13_striginternallto23_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_speriod_cry_23_c_RNIHTOK1_LC_9_12_3.C_ON=1'b0;
    defparam un4_speriod_cry_23_c_RNIHTOK1_LC_9_12_3.SEQ_MODE=4'b0000;
    defparam un4_speriod_cry_23_c_RNIHTOK1_LC_9_12_3.LUT_INIT=16'b0000000010110000;
    LogicCell40 un4_speriod_cry_23_c_RNIHTOK1_LC_9_12_3 (
            .in0(N__24944),
            .in1(N__29060),
            .in2(N__24843),
            .in3(N__24790),
            .lcout(),
            .ltout(un1_reset_rpi_inv_2_i_1_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIT8E57_4_LC_9_12_4.C_ON=1'b0;
    defparam sCounter_RNIT8E57_4_LC_9_12_4.SEQ_MODE=4'b0000;
    defparam sCounter_RNIT8E57_4_LC_9_12_4.LUT_INIT=16'b1111011111010101;
    LogicCell40 sCounter_RNIT8E57_4_LC_9_12_4 (
            .in0(N__32547),
            .in1(N__36957),
            .in2(N__24747),
            .in3(N__36844),
            .lcout(un1_reset_rpi_inv_2_i_1),
            .ltout(un1_reset_rpi_inv_2_i_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sTrigCounter_6_LC_9_12_5.C_ON=1'b0;
    defparam sTrigCounter_6_LC_9_12_5.SEQ_MODE=4'b1000;
    defparam sTrigCounter_6_LC_9_12_5.LUT_INIT=16'b1100001111001100;
    LogicCell40 sTrigCounter_6_LC_9_12_5 (
            .in0(_gnd_net_),
            .in1(N__25075),
            .in2(N__25089),
            .in3(N__25086),
            .lcout(sTrigCounterZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47790),
            .ce(),
            .sr(N__27536));
    defparam sTrigCounter_7_LC_9_12_6.C_ON=1'b0;
    defparam sTrigCounter_7_LC_9_12_6.SEQ_MODE=4'b1000;
    defparam sTrigCounter_7_LC_9_12_6.LUT_INIT=16'b1111000011010010;
    LogicCell40 sTrigCounter_7_LC_9_12_6 (
            .in0(N__25056),
            .in1(N__25047),
            .in2(N__25031),
            .in3(N__25041),
            .lcout(sTrigCounterZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47790),
            .ce(),
            .sr(N__27536));
    defparam un1_spoff_cry_0_c_inv_LC_9_13_0.C_ON=1'b1;
    defparam un1_spoff_cry_0_c_inv_LC_9_13_0.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_0_c_inv_LC_9_13_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_0_c_inv_LC_9_13_0 (
            .in0(_gnd_net_),
            .in1(N__29316),
            .in2(N__26169),
            .in3(N__34200),
            .lcout(sCounter_i_0),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(un1_spoff_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_1_c_inv_LC_9_13_1.C_ON=1'b1;
    defparam un1_spoff_cry_1_c_inv_LC_9_13_1.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_1_c_inv_LC_9_13_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_1_c_inv_LC_9_13_1 (
            .in0(_gnd_net_),
            .in1(N__26151),
            .in2(N__29307),
            .in3(N__35023),
            .lcout(sCounter_i_1),
            .ltout(),
            .carryin(un1_spoff_cry_0),
            .carryout(un1_spoff_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_2_c_inv_LC_9_13_2.C_ON=1'b1;
    defparam un1_spoff_cry_2_c_inv_LC_9_13_2.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_2_c_inv_LC_9_13_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_2_c_inv_LC_9_13_2 (
            .in0(_gnd_net_),
            .in1(N__29292),
            .in2(N__26460),
            .in3(N__34925),
            .lcout(sCounter_i_2),
            .ltout(),
            .carryin(un1_spoff_cry_1),
            .carryout(un1_spoff_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_3_c_inv_LC_9_13_3.C_ON=1'b1;
    defparam un1_spoff_cry_3_c_inv_LC_9_13_3.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_3_c_inv_LC_9_13_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_3_c_inv_LC_9_13_3 (
            .in0(_gnd_net_),
            .in1(N__29283),
            .in2(N__26442),
            .in3(N__34817),
            .lcout(sCounter_i_3),
            .ltout(),
            .carryin(un1_spoff_cry_2),
            .carryout(un1_spoff_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_4_c_inv_LC_9_13_4.C_ON=1'b1;
    defparam un1_spoff_cry_4_c_inv_LC_9_13_4.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_4_c_inv_LC_9_13_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_4_c_inv_LC_9_13_4 (
            .in0(_gnd_net_),
            .in1(N__29274),
            .in2(N__26424),
            .in3(N__36782),
            .lcout(sCounter_i_4),
            .ltout(),
            .carryin(un1_spoff_cry_3),
            .carryout(un1_spoff_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_5_c_inv_LC_9_13_5.C_ON=1'b1;
    defparam un1_spoff_cry_5_c_inv_LC_9_13_5.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_5_c_inv_LC_9_13_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_5_c_inv_LC_9_13_5 (
            .in0(_gnd_net_),
            .in1(N__29265),
            .in2(N__26406),
            .in3(N__34691),
            .lcout(sCounter_i_5),
            .ltout(),
            .carryin(un1_spoff_cry_4),
            .carryout(un1_spoff_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_6_c_inv_LC_9_13_6.C_ON=1'b1;
    defparam un1_spoff_cry_6_c_inv_LC_9_13_6.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_6_c_inv_LC_9_13_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_6_c_inv_LC_9_13_6 (
            .in0(_gnd_net_),
            .in1(N__29256),
            .in2(N__26388),
            .in3(N__34567),
            .lcout(sCounter_i_6),
            .ltout(),
            .carryin(un1_spoff_cry_5),
            .carryout(un1_spoff_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_7_c_inv_LC_9_13_7.C_ON=1'b1;
    defparam un1_spoff_cry_7_c_inv_LC_9_13_7.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_7_c_inv_LC_9_13_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_spoff_cry_7_c_inv_LC_9_13_7 (
            .in0(N__34445),
            .in1(N__29247),
            .in2(N__26370),
            .in3(_gnd_net_),
            .lcout(sCounter_i_7),
            .ltout(),
            .carryin(un1_spoff_cry_6),
            .carryout(un1_spoff_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_8_c_inv_LC_9_14_0.C_ON=1'b1;
    defparam un1_spoff_cry_8_c_inv_LC_9_14_0.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_8_c_inv_LC_9_14_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_8_c_inv_LC_9_14_0 (
            .in0(_gnd_net_),
            .in1(N__29355),
            .in2(N__26349),
            .in3(N__35842),
            .lcout(sCounter_i_8),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(un1_spoff_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_9_c_inv_LC_9_14_1.C_ON=1'b1;
    defparam un1_spoff_cry_9_c_inv_LC_9_14_1.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_9_c_inv_LC_9_14_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_9_c_inv_LC_9_14_1 (
            .in0(_gnd_net_),
            .in1(N__29346),
            .in2(N__26331),
            .in3(N__35731),
            .lcout(sCounter_i_9),
            .ltout(),
            .carryin(un1_spoff_cry_8),
            .carryout(un1_spoff_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_10_c_inv_LC_9_14_2.C_ON=1'b1;
    defparam un1_spoff_cry_10_c_inv_LC_9_14_2.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_10_c_inv_LC_9_14_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_10_c_inv_LC_9_14_2 (
            .in0(_gnd_net_),
            .in1(N__29238),
            .in2(N__26583),
            .in3(N__35617),
            .lcout(sCounter_i_10),
            .ltout(),
            .carryin(un1_spoff_cry_9),
            .carryout(un1_spoff_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_11_c_inv_LC_9_14_3.C_ON=1'b1;
    defparam un1_spoff_cry_11_c_inv_LC_9_14_3.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_11_c_inv_LC_9_14_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_11_c_inv_LC_9_14_3 (
            .in0(_gnd_net_),
            .in1(N__29409),
            .in2(N__26565),
            .in3(N__35496),
            .lcout(sCounter_i_11),
            .ltout(),
            .carryin(un1_spoff_cry_10),
            .carryout(un1_spoff_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_12_c_inv_LC_9_14_4.C_ON=1'b1;
    defparam un1_spoff_cry_12_c_inv_LC_9_14_4.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_12_c_inv_LC_9_14_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_12_c_inv_LC_9_14_4 (
            .in0(_gnd_net_),
            .in1(N__29397),
            .in2(N__26547),
            .in3(N__35369),
            .lcout(sCounter_i_12),
            .ltout(),
            .carryin(un1_spoff_cry_11),
            .carryout(un1_spoff_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_13_c_inv_LC_9_14_5.C_ON=1'b1;
    defparam un1_spoff_cry_13_c_inv_LC_9_14_5.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_13_c_inv_LC_9_14_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_13_c_inv_LC_9_14_5 (
            .in0(_gnd_net_),
            .in1(N__29385),
            .in2(N__26529),
            .in3(N__35284),
            .lcout(sCounter_i_13),
            .ltout(),
            .carryin(un1_spoff_cry_12),
            .carryout(un1_spoff_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_14_c_inv_LC_9_14_6.C_ON=1'b1;
    defparam un1_spoff_cry_14_c_inv_LC_9_14_6.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_14_c_inv_LC_9_14_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_14_c_inv_LC_9_14_6 (
            .in0(_gnd_net_),
            .in1(N__29376),
            .in2(N__26511),
            .in3(N__35156),
            .lcout(sCounter_i_14),
            .ltout(),
            .carryin(un1_spoff_cry_13),
            .carryout(un1_spoff_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_15_c_inv_LC_9_14_7.C_ON=1'b1;
    defparam un1_spoff_cry_15_c_inv_LC_9_14_7.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_15_c_inv_LC_9_14_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_15_c_inv_LC_9_14_7 (
            .in0(_gnd_net_),
            .in1(N__26492),
            .in2(N__29367),
            .in3(N__36616),
            .lcout(sCounter_i_15),
            .ltout(),
            .carryin(un1_spoff_cry_14),
            .carryout(un1_spoff_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_16_c_inv_LC_9_15_0.C_ON=1'b1;
    defparam un1_spoff_cry_16_c_inv_LC_9_15_0.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_16_c_inv_LC_9_15_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_16_c_inv_LC_9_15_0 (
            .in0(_gnd_net_),
            .in1(N__25137),
            .in2(_gnd_net_),
            .in3(N__36507),
            .lcout(sCounter_i_16),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(un1_spoff_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_17_c_inv_LC_9_15_1.C_ON=1'b1;
    defparam un1_spoff_cry_17_c_inv_LC_9_15_1.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_17_c_inv_LC_9_15_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_spoff_cry_17_c_inv_LC_9_15_1 (
            .in0(N__36406),
            .in1(N__25131),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sCounter_i_17),
            .ltout(),
            .carryin(un1_spoff_cry_16),
            .carryout(un1_spoff_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_18_c_inv_LC_9_15_2.C_ON=1'b1;
    defparam un1_spoff_cry_18_c_inv_LC_9_15_2.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_18_c_inv_LC_9_15_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_spoff_cry_18_c_inv_LC_9_15_2 (
            .in0(N__36310),
            .in1(N__25125),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sCounter_i_18),
            .ltout(),
            .carryin(un1_spoff_cry_17),
            .carryout(un1_spoff_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_19_c_inv_LC_9_15_3.C_ON=1'b1;
    defparam un1_spoff_cry_19_c_inv_LC_9_15_3.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_19_c_inv_LC_9_15_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_19_c_inv_LC_9_15_3 (
            .in0(_gnd_net_),
            .in1(N__25119),
            .in2(_gnd_net_),
            .in3(N__36230),
            .lcout(sCounter_i_19),
            .ltout(),
            .carryin(un1_spoff_cry_18),
            .carryout(un1_spoff_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_20_c_inv_LC_9_15_4.C_ON=1'b1;
    defparam un1_spoff_cry_20_c_inv_LC_9_15_4.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_20_c_inv_LC_9_15_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_20_c_inv_LC_9_15_4 (
            .in0(_gnd_net_),
            .in1(N__25113),
            .in2(_gnd_net_),
            .in3(N__36137),
            .lcout(sCounter_i_20),
            .ltout(),
            .carryin(un1_spoff_cry_19),
            .carryout(un1_spoff_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_21_c_inv_LC_9_15_5.C_ON=1'b1;
    defparam un1_spoff_cry_21_c_inv_LC_9_15_5.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_21_c_inv_LC_9_15_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_21_c_inv_LC_9_15_5 (
            .in0(_gnd_net_),
            .in1(N__25107),
            .in2(_gnd_net_),
            .in3(N__36053),
            .lcout(sCounter_i_21),
            .ltout(),
            .carryin(un1_spoff_cry_20),
            .carryout(un1_spoff_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_22_c_inv_LC_9_15_6.C_ON=1'b1;
    defparam un1_spoff_cry_22_c_inv_LC_9_15_6.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_22_c_inv_LC_9_15_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_spoff_cry_22_c_inv_LC_9_15_6 (
            .in0(N__35951),
            .in1(N__25101),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sCounter_i_22),
            .ltout(),
            .carryin(un1_spoff_cry_21),
            .carryout(un1_spoff_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_spoff_cry_23_c_inv_LC_9_15_7.C_ON=1'b1;
    defparam un1_spoff_cry_23_c_inv_LC_9_15_7.SEQ_MODE=4'b0000;
    defparam un1_spoff_cry_23_c_inv_LC_9_15_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_spoff_cry_23_c_inv_LC_9_15_7 (
            .in0(_gnd_net_),
            .in1(N__25095),
            .in2(_gnd_net_),
            .in3(N__37054),
            .lcout(sCounter_i_23),
            .ltout(),
            .carryin(un1_spoff_cry_22),
            .carryout(un1_spoff_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam poff_obuf_RNO_LC_9_16_0.C_ON=1'b0;
    defparam poff_obuf_RNO_LC_9_16_0.SEQ_MODE=4'b0000;
    defparam poff_obuf_RNO_LC_9_16_0.LUT_INIT=16'b0011001111111111;
    LogicCell40 poff_obuf_RNO_LC_9_16_0 (
            .in0(_gnd_net_),
            .in1(N__25350),
            .in2(_gnd_net_),
            .in3(N__25338),
            .lcout(N_1612_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sRead_data_RNI74VQ_LC_9_16_1.C_ON=1'b0;
    defparam sRead_data_RNI74VQ_LC_9_16_1.SEQ_MODE=4'b0000;
    defparam sRead_data_RNI74VQ_LC_9_16_1.LUT_INIT=16'b1101110111111111;
    LogicCell40 sRead_data_RNI74VQ_LC_9_16_1 (
            .in0(N__27474),
            .in1(N__25322),
            .in2(_gnd_net_),
            .in3(N__25308),
            .lcout(spi_data_miso_0_sqmuxa_2_i_o2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_1_LC_9_16_3.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_1_LC_9_16_3.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_1_LC_9_16_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_1_LC_9_16_3 (
            .in0(N__26309),
            .in1(N__25293),
            .in2(N__25275),
            .in3(N__25254),
            .lcout(sbuttonModeStatus_0_sqmuxa_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sbuttonModeStatus_RNO_4_LC_9_16_7.C_ON=1'b0;
    defparam sbuttonModeStatus_RNO_4_LC_9_16_7.SEQ_MODE=4'b0000;
    defparam sbuttonModeStatus_RNO_4_LC_9_16_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 sbuttonModeStatus_RNO_4_LC_9_16_7 (
            .in0(N__25235),
            .in1(N__25223),
            .in2(N__25212),
            .in3(N__25196),
            .lcout(sbuttonModeStatus_0_sqmuxa_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_0_c_inv_LC_9_17_0.C_ON=1'b1;
    defparam un4_sacqtime_cry_0_c_inv_LC_9_17_0.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_0_c_inv_LC_9_17_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_0_c_inv_LC_9_17_0 (
            .in0(_gnd_net_),
            .in1(N__34226),
            .in2(N__25173),
            .in3(N__26739),
            .lcout(sEEDelayACQ_i_0),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(un4_sacqtime_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_1_c_inv_LC_9_17_1.C_ON=1'b1;
    defparam un4_sacqtime_cry_1_c_inv_LC_9_17_1.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_1_c_inv_LC_9_17_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_1_c_inv_LC_9_17_1 (
            .in0(_gnd_net_),
            .in1(N__35051),
            .in2(N__25164),
            .in3(N__26733),
            .lcout(sEEDelayACQ_i_1),
            .ltout(),
            .carryin(un4_sacqtime_cry_0),
            .carryout(un4_sacqtime_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_2_c_inv_LC_9_17_2.C_ON=1'b1;
    defparam un4_sacqtime_cry_2_c_inv_LC_9_17_2.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_2_c_inv_LC_9_17_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_2_c_inv_LC_9_17_2 (
            .in0(_gnd_net_),
            .in1(N__34942),
            .in2(N__25155),
            .in3(N__26727),
            .lcout(sEEDelayACQ_i_2),
            .ltout(),
            .carryin(un4_sacqtime_cry_1),
            .carryout(un4_sacqtime_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_3_c_inv_LC_9_17_3.C_ON=1'b1;
    defparam un4_sacqtime_cry_3_c_inv_LC_9_17_3.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_3_c_inv_LC_9_17_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_3_c_inv_LC_9_17_3 (
            .in0(_gnd_net_),
            .in1(N__34835),
            .in2(N__25146),
            .in3(N__26721),
            .lcout(sEEDelayACQ_i_3),
            .ltout(),
            .carryin(un4_sacqtime_cry_2),
            .carryout(un4_sacqtime_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_4_c_inv_LC_9_17_4.C_ON=1'b1;
    defparam un4_sacqtime_cry_4_c_inv_LC_9_17_4.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_4_c_inv_LC_9_17_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_sacqtime_cry_4_c_inv_LC_9_17_4 (
            .in0(N__26715),
            .in1(N__36819),
            .in2(N__25419),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQ_i_4),
            .ltout(),
            .carryin(un4_sacqtime_cry_3),
            .carryout(un4_sacqtime_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_5_c_inv_LC_9_17_5.C_ON=1'b1;
    defparam un4_sacqtime_cry_5_c_inv_LC_9_17_5.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_5_c_inv_LC_9_17_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_5_c_inv_LC_9_17_5 (
            .in0(_gnd_net_),
            .in1(N__34706),
            .in2(N__25410),
            .in3(N__26709),
            .lcout(sEEDelayACQ_i_5),
            .ltout(),
            .carryin(un4_sacqtime_cry_4),
            .carryout(un4_sacqtime_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_6_c_inv_LC_9_17_6.C_ON=1'b1;
    defparam un4_sacqtime_cry_6_c_inv_LC_9_17_6.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_6_c_inv_LC_9_17_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_6_c_inv_LC_9_17_6 (
            .in0(_gnd_net_),
            .in1(N__34601),
            .in2(N__25401),
            .in3(N__26808),
            .lcout(sEEDelayACQ_i_6),
            .ltout(),
            .carryin(un4_sacqtime_cry_5),
            .carryout(un4_sacqtime_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_7_c_inv_LC_9_17_7.C_ON=1'b1;
    defparam un4_sacqtime_cry_7_c_inv_LC_9_17_7.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_7_c_inv_LC_9_17_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un4_sacqtime_cry_7_c_inv_LC_9_17_7 (
            .in0(N__26802),
            .in1(N__25392),
            .in2(N__34475),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQ_i_7),
            .ltout(),
            .carryin(un4_sacqtime_cry_6),
            .carryout(un4_sacqtime_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_8_c_inv_LC_9_18_0.C_ON=1'b1;
    defparam un4_sacqtime_cry_8_c_inv_LC_9_18_0.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_8_c_inv_LC_9_18_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_8_c_inv_LC_9_18_0 (
            .in0(_gnd_net_),
            .in1(N__35870),
            .in2(N__25386),
            .in3(N__26760),
            .lcout(sEEDelayACQ_i_8),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(un4_sacqtime_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_9_c_inv_LC_9_18_1.C_ON=1'b1;
    defparam un4_sacqtime_cry_9_c_inv_LC_9_18_1.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_9_c_inv_LC_9_18_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_9_c_inv_LC_9_18_1 (
            .in0(_gnd_net_),
            .in1(N__35768),
            .in2(N__25377),
            .in3(N__26952),
            .lcout(sEEDelayACQ_i_9),
            .ltout(),
            .carryin(un4_sacqtime_cry_8),
            .carryout(un4_sacqtime_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_10_c_inv_LC_9_18_2.C_ON=1'b1;
    defparam un4_sacqtime_cry_10_c_inv_LC_9_18_2.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_10_c_inv_LC_9_18_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_10_c_inv_LC_9_18_2 (
            .in0(_gnd_net_),
            .in1(N__35633),
            .in2(N__25368),
            .in3(N__26796),
            .lcout(sEEDelayACQ_i_10),
            .ltout(),
            .carryin(un4_sacqtime_cry_9),
            .carryout(un4_sacqtime_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_11_c_inv_LC_9_18_3.C_ON=1'b1;
    defparam un4_sacqtime_cry_11_c_inv_LC_9_18_3.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_11_c_inv_LC_9_18_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_11_c_inv_LC_9_18_3 (
            .in0(_gnd_net_),
            .in1(N__35520),
            .in2(N__25359),
            .in3(N__26790),
            .lcout(sEEDelayACQ_i_11),
            .ltout(),
            .carryin(un4_sacqtime_cry_10),
            .carryout(un4_sacqtime_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_12_c_inv_LC_9_18_4.C_ON=1'b1;
    defparam un4_sacqtime_cry_12_c_inv_LC_9_18_4.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_12_c_inv_LC_9_18_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_12_c_inv_LC_9_18_4 (
            .in0(_gnd_net_),
            .in1(N__35384),
            .in2(N__25452),
            .in3(N__26784),
            .lcout(sEEDelayACQ_i_12),
            .ltout(),
            .carryin(un4_sacqtime_cry_11),
            .carryout(un4_sacqtime_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_13_c_inv_LC_9_18_5.C_ON=1'b1;
    defparam un4_sacqtime_cry_13_c_inv_LC_9_18_5.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_13_c_inv_LC_9_18_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_13_c_inv_LC_9_18_5 (
            .in0(_gnd_net_),
            .in1(N__35302),
            .in2(N__25443),
            .in3(N__26778),
            .lcout(sEEDelayACQ_i_13),
            .ltout(),
            .carryin(un4_sacqtime_cry_12),
            .carryout(un4_sacqtime_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_14_c_inv_LC_9_18_6.C_ON=1'b1;
    defparam un4_sacqtime_cry_14_c_inv_LC_9_18_6.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_14_c_inv_LC_9_18_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_14_c_inv_LC_9_18_6 (
            .in0(_gnd_net_),
            .in1(N__35188),
            .in2(N__25434),
            .in3(N__26772),
            .lcout(sEEDelayACQ_i_14),
            .ltout(),
            .carryin(un4_sacqtime_cry_13),
            .carryout(un4_sacqtime_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_15_c_inv_LC_9_18_7.C_ON=1'b1;
    defparam un4_sacqtime_cry_15_c_inv_LC_9_18_7.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_15_c_inv_LC_9_18_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un4_sacqtime_cry_15_c_inv_LC_9_18_7 (
            .in0(_gnd_net_),
            .in1(N__25425),
            .in2(N__36653),
            .in3(N__26766),
            .lcout(sEEDelayACQ_i_15),
            .ltout(),
            .carryin(un4_sacqtime_cry_14),
            .carryout(un4_sacqtime_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_16_c_LC_9_19_0.C_ON=1'b1;
    defparam un4_sacqtime_cry_16_c_LC_9_19_0.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_16_c_LC_9_19_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_16_c_LC_9_19_0 (
            .in0(_gnd_net_),
            .in1(N__36530),
            .in2(N__38072),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(un4_sacqtime_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_17_c_LC_9_19_1.C_ON=1'b1;
    defparam un4_sacqtime_cry_17_c_LC_9_19_1.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_17_c_LC_9_19_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_17_c_LC_9_19_1 (
            .in0(_gnd_net_),
            .in1(N__36431),
            .in2(N__38070),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_sacqtime_cry_16),
            .carryout(un4_sacqtime_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_18_c_LC_9_19_2.C_ON=1'b1;
    defparam un4_sacqtime_cry_18_c_LC_9_19_2.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_18_c_LC_9_19_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_18_c_LC_9_19_2 (
            .in0(_gnd_net_),
            .in1(N__36328),
            .in2(N__38073),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_sacqtime_cry_17),
            .carryout(un4_sacqtime_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_19_c_LC_9_19_3.C_ON=1'b1;
    defparam un4_sacqtime_cry_19_c_LC_9_19_3.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_19_c_LC_9_19_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_19_c_LC_9_19_3 (
            .in0(_gnd_net_),
            .in1(N__36247),
            .in2(N__38071),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_sacqtime_cry_18),
            .carryout(un4_sacqtime_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_20_c_LC_9_19_4.C_ON=1'b1;
    defparam un4_sacqtime_cry_20_c_LC_9_19_4.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_20_c_LC_9_19_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_20_c_LC_9_19_4 (
            .in0(_gnd_net_),
            .in1(N__36147),
            .in2(N__38074),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_sacqtime_cry_19),
            .carryout(un4_sacqtime_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounter_RNIR3KA_0_20_LC_9_19_5.C_ON=1'b1;
    defparam sCounter_RNIR3KA_0_20_LC_9_19_5.SEQ_MODE=4'b0000;
    defparam sCounter_RNIR3KA_0_20_LC_9_19_5.LUT_INIT=16'b0001000100010001;
    LogicCell40 sCounter_RNIR3KA_0_20_LC_9_19_5 (
            .in0(N__36148),
            .in1(N__36065),
            .in2(N__38069),
            .in3(_gnd_net_),
            .lcout(op_gt_op_gt_un13_striginternallto23_8),
            .ltout(),
            .carryin(un4_sacqtime_cry_20),
            .carryout(un4_sacqtime_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_22_c_LC_9_19_6.C_ON=1'b1;
    defparam un4_sacqtime_cry_22_c_LC_9_19_6.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_22_c_LC_9_19_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_22_c_LC_9_19_6 (
            .in0(_gnd_net_),
            .in1(N__38033),
            .in2(N__35980),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_sacqtime_cry_21),
            .carryout(un4_sacqtime_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_23_c_LC_9_19_7.C_ON=1'b1;
    defparam un4_sacqtime_cry_23_c_LC_9_19_7.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_23_c_LC_9_19_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un4_sacqtime_cry_23_c_LC_9_19_7 (
            .in0(_gnd_net_),
            .in1(N__38043),
            .in2(N__37083),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un4_sacqtime_cry_22),
            .carryout(un4_sacqtime_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_23_THRU_LUT4_0_LC_9_20_0.C_ON=1'b0;
    defparam un4_sacqtime_cry_23_THRU_LUT4_0_LC_9_20_0.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_23_THRU_LUT4_0_LC_9_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un4_sacqtime_cry_23_THRU_LUT4_0_LC_9_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25473),
            .lcout(un4_sacqtime_cry_23_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam button_debounce_counter_esr_RNO_0_23_LC_9_20_1.C_ON=1'b0;
    defparam button_debounce_counter_esr_RNO_0_23_LC_9_20_1.SEQ_MODE=4'b0000;
    defparam button_debounce_counter_esr_RNO_0_23_LC_9_20_1.LUT_INIT=16'b1111111110101010;
    LogicCell40 button_debounce_counter_esr_RNO_0_23_LC_9_20_1 (
            .in0(N__32624),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26250),
            .lcout(LED3_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_0_LC_10_2_0 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_0_LC_10_2_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_0_LC_10_2_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_0_LC_10_2_0  (
            .in0(N__26826),
            .in1(N__25661),
            .in2(N__25605),
            .in3(N__25604),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_2_0_),
            .carryout(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0 ),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53124));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_1_LC_10_2_1 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_1_LC_10_2_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_1_LC_10_2_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_1_LC_10_2_1  (
            .in0(N__26828),
            .in1(N__25674),
            .in2(_gnd_net_),
            .in3(N__25461),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_1 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_0 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1 ),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53124));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_2_LC_10_2_2 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_2_LC_10_2_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_2_LC_10_2_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_2_LC_10_2_2  (
            .in0(N__26827),
            .in1(N__25620),
            .in2(_gnd_net_),
            .in3(N__25458),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_2 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_1 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2 ),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53124));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_3_LC_10_2_3 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_3_LC_10_2_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_3_LC_10_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_3_LC_10_2_3  (
            .in0(_gnd_net_),
            .in1(N__25647),
            .in2(_gnd_net_),
            .in3(N__25455),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_2 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3 ),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53124));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_4_LC_10_2_4 .C_ON=1'b1;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_4_LC_10_2_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_4_LC_10_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_4_LC_10_2_4  (
            .in0(_gnd_net_),
            .in1(N__25686),
            .in2(_gnd_net_),
            .in3(N__25692),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_3 ),
            .carryout(\spi_slave_inst.un1_rx_data_count_neg_sclk_i_cry_4 ),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53124));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_5_LC_10_2_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_5_LC_10_2_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_5_LC_10_2_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_5_LC_10_2_5  (
            .in0(_gnd_net_),
            .in1(N__25635),
            .in2(_gnd_net_),
            .in3(N__25689),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVspi_slave_inst.rx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53124));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNICMDR1_0_LC_10_3_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNICMDR1_0_LC_10_3_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNICMDR1_0_LC_10_3_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_RNICMDR1_0_LC_10_3_0  (
            .in0(N__25685),
            .in1(N__25673),
            .in2(N__25662),
            .in3(N__25646),
            .lcout(),
            .ltout(\spi_slave_inst.rx_data_count_neg_sclk_i6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNILK4P2_5_LC_10_3_1 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNILK4P2_5_LC_10_3_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNILK4P2_5_LC_10_3_1 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_RNILK4P2_5_LC_10_3_1  (
            .in0(N__25634),
            .in1(_gnd_net_),
            .in2(N__25623),
            .in3(N__25619),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_i6 ),
            .ltout(\spi_slave_inst.rx_data_count_neg_sclk_i6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3_5_LC_10_3_2 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3_5_LC_10_3_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3_5_LC_10_3_2 .LUT_INIT=16'b0000010000000111;
    LogicCell40 \spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3_5_LC_10_3_2  (
            .in0(N__52419),
            .in1(N__38525),
            .in2(N__25608),
            .in3(N__33286),
            .lcout(\spi_slave_inst.rx_data_count_neg_sclk_i_RNIKVPI3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNICH5T1_0_LC_10_3_4 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNICH5T1_0_LC_10_3_4 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNICH5T1_0_LC_10_3_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_RNICH5T1_0_LC_10_3_4  (
            .in0(N__25589),
            .in1(N__25573),
            .in2(N__25556),
            .in3(N__25532),
            .lcout(\spi_slave_inst.un23_i_ssn_3 ),
            .ltout(\spi_slave_inst.un23_i_ssn_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI5DOR2_5_LC_10_3_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI5DOR2_5_LC_10_3_5 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI5DOR2_5_LC_10_3_5 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_RNI5DOR2_5_LC_10_3_5  (
            .in0(_gnd_net_),
            .in1(N__25795),
            .in2(N__25521),
            .in3(N__25773),
            .lcout(\spi_slave_inst.un23_i_ssn ),
            .ltout(\spi_slave_inst.un23_i_ssn_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI4ODL3_5_LC_10_3_6 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI4ODL3_5_LC_10_3_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_data_count_pos_sclk_i_RNI4ODL3_5_LC_10_3_6 .LUT_INIT=16'b0000010000000111;
    LogicCell40 \spi_slave_inst.rx_data_count_pos_sclk_i_RNI4ODL3_5_LC_10_3_6  (
            .in0(N__52420),
            .in1(N__38526),
            .in2(N__25506),
            .in3(N__33287),
            .lcout(\spi_slave_inst.rx_data_count_pos_sclk_i_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.spi_cs_i_LC_10_3_7 .C_ON=1'b0;
    defparam \spi_slave_inst.spi_cs_i_LC_10_3_7 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.spi_cs_i_LC_10_3_7 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \spi_slave_inst.spi_cs_i_LC_10_3_7  (
            .in0(N__38527),
            .in1(_gnd_net_),
            .in2(N__33291),
            .in3(N__52421),
            .lcout(\spi_slave_inst.spi_cs_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_done_pos_sclk_i_LC_10_4_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_pos_sclk_i_LC_10_4_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_done_pos_sclk_i_LC_10_4_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \spi_slave_inst.rx_done_pos_sclk_i_LC_10_4_0  (
            .in0(N__25803),
            .in1(N__25797),
            .in2(_gnd_net_),
            .in3(N__25778),
            .lcout(\spi_slave_inst.rx_done_pos_sclk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30704),
            .ce(N__30664),
            .sr(N__53095));
    defparam \spi_master_inst.spi_data_path_u1.data_in_6_LC_10_5_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_6_LC_10_5_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_6_LC_10_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_6_LC_10_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42252),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53247),
            .ce(N__28842),
            .sr(N__53082));
    defparam \spi_master_inst.spi_data_path_u1.data_in_1_LC_10_5_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_1_LC_10_5_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_1_LC_10_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_1_LC_10_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37623),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53247),
            .ce(N__28842),
            .sr(N__53082));
    defparam \spi_master_inst.spi_data_path_u1.data_in_2_LC_10_5_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_2_LC_10_5_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_2_LC_10_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_2_LC_10_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26841),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53247),
            .ce(N__28842),
            .sr(N__53082));
    defparam \spi_master_inst.spi_data_path_u1.data_in_11_LC_10_5_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_11_LC_10_5_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_11_LC_10_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_11_LC_10_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37605),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53247),
            .ce(N__28842),
            .sr(N__53082));
    defparam \spi_master_inst.spi_data_path_u1.data_in_12_LC_10_5_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_12_LC_10_5_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_12_LC_10_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_12_LC_10_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37587),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53247),
            .ce(N__28842),
            .sr(N__53082));
    defparam \spi_master_inst.spi_data_path_u1.data_in_3_LC_10_5_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_3_LC_10_5_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_3_LC_10_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_3_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41370),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53247),
            .ce(N__28842),
            .sr(N__53082));
    defparam \spi_master_inst.spi_data_path_u1.data_in_14_LC_10_5_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_14_LC_10_5_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_14_LC_10_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_14_LC_10_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37719),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53247),
            .ce(N__28842),
            .sr(N__53082));
    defparam \spi_master_inst.spi_data_path_u1.data_in_15_LC_10_5_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_15_LC_10_5_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_15_LC_10_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_15_LC_10_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37701),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53247),
            .ce(N__28842),
            .sr(N__53082));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_0_LC_10_6_0 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_0_LC_10_6_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_0_LC_10_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_0_LC_10_6_0  (
            .in0(N__25864),
            .in1(N__25980),
            .in2(_gnd_net_),
            .in3(N__25968),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_6_0_),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0 ),
            .clk(N__53251),
            .ce(N__25818),
            .sr(N__53070));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_1_LC_10_6_1 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_1_LC_10_6_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_1_LC_10_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_1_LC_10_6_1  (
            .in0(N__25859),
            .in1(N__25965),
            .in2(_gnd_net_),
            .in3(N__25950),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_1 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_0 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1 ),
            .clk(N__53251),
            .ce(N__25818),
            .sr(N__53070));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_2_LC_10_6_2 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_2_LC_10_6_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_2_LC_10_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_2_LC_10_6_2  (
            .in0(N__25865),
            .in1(N__25946),
            .in2(_gnd_net_),
            .in3(N__25932),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_2 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_1 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2 ),
            .clk(N__53251),
            .ce(N__25818),
            .sr(N__53070));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_3_LC_10_6_3 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_3_LC_10_6_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_3_LC_10_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_3_LC_10_6_3  (
            .in0(N__25860),
            .in1(N__25929),
            .in2(_gnd_net_),
            .in3(N__25917),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_2 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3 ),
            .clk(N__53251),
            .ce(N__25818),
            .sr(N__53070));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_4_LC_10_6_4 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_4_LC_10_6_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_4_LC_10_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_4_LC_10_6_4  (
            .in0(N__25866),
            .in1(N__25914),
            .in2(_gnd_net_),
            .in3(N__25902),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_3 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4 ),
            .clk(N__53251),
            .ce(N__25818),
            .sr(N__53070));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_5_LC_10_6_5 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_5_LC_10_6_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_5_LC_10_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_5_LC_10_6_5  (
            .in0(N__25861),
            .in1(N__25899),
            .in2(_gnd_net_),
            .in3(N__25887),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_5 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_4 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5 ),
            .clk(N__53251),
            .ce(N__25818),
            .sr(N__53070));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_6_LC_10_6_6 .C_ON=1'b1;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_6_LC_10_6_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_6_LC_10_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_6_LC_10_6_6  (
            .in0(N__25862),
            .in1(N__25883),
            .in2(_gnd_net_),
            .in3(N__25869),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_6 ),
            .ltout(),
            .carryin(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_5 ),
            .carryout(\spi_master_inst.sclk_gen_u0.clk_falling_count_i_cry_6 ),
            .clk(N__53251),
            .ce(N__25818),
            .sr(N__53070));
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_7_LC_10_6_7 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_7_LC_10_6_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.clk_falling_count_i_7_LC_10_6_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \spi_master_inst.sclk_gen_u0.clk_falling_count_i_7_LC_10_6_7  (
            .in0(N__25830),
            .in1(N__25863),
            .in2(_gnd_net_),
            .in3(N__25833),
            .lcout(\spi_master_inst.sclk_gen_u0.clk_falling_count_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53251),
            .ce(N__25818),
            .sr(N__53070));
    defparam sEETrigCounter_0_LC_10_7_1.C_ON=1'b0;
    defparam sEETrigCounter_0_LC_10_7_1.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_0_LC_10_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_0_LC_10_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51041),
            .lcout(sEETrigCounterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47814),
            .ce(N__31016),
            .sr(N__53059));
    defparam sEETrigCounter_1_LC_10_7_5.C_ON=1'b0;
    defparam sEETrigCounter_1_LC_10_7_5.SEQ_MODE=4'b1011;
    defparam sEETrigCounter_1_LC_10_7_5.LUT_INIT=16'b1100110011001100;
    LogicCell40 sEETrigCounter_1_LC_10_7_5 (
            .in0(_gnd_net_),
            .in1(N__50692),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEETrigCounterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47814),
            .ce(N__31016),
            .sr(N__53059));
    defparam sEETrigCounter_2_LC_10_7_6.C_ON=1'b0;
    defparam sEETrigCounter_2_LC_10_7_6.SEQ_MODE=4'b1010;
    defparam sEETrigCounter_2_LC_10_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_2_LC_10_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50123),
            .lcout(sEETrigCounterZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47814),
            .ce(N__31016),
            .sr(N__53059));
    defparam sEETrigCounter_3_LC_10_7_7.C_ON=1'b0;
    defparam sEETrigCounter_3_LC_10_7_7.SEQ_MODE=4'b1011;
    defparam sEETrigCounter_3_LC_10_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEETrigCounter_3_LC_10_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49651),
            .lcout(sEETrigCounterZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47814),
            .ce(N__31016),
            .sr(N__53059));
    defparam sEETrigCounter_RNII1HP1_2_LC_10_8_0.C_ON=1'b0;
    defparam sEETrigCounter_RNII1HP1_2_LC_10_8_0.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNII1HP1_2_LC_10_8_0.LUT_INIT=16'b1111000011100001;
    LogicCell40 sEETrigCounter_RNII1HP1_2_LC_10_8_0 (
            .in0(N__26081),
            .in1(N__26042),
            .in2(N__26121),
            .in3(N__26014),
            .lcout(un10_trig_prev_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIKN4B1_2_LC_10_8_1.C_ON=1'b0;
    defparam sEETrigCounter_RNIKN4B1_2_LC_10_8_1.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIKN4B1_2_LC_10_8_1.LUT_INIT=16'b1111101000000101;
    LogicCell40 sEETrigCounter_RNIKN4B1_2_LC_10_8_1 (
            .in0(N__26016),
            .in1(_gnd_net_),
            .in2(N__26043),
            .in3(N__26080),
            .lcout(un10_trig_prev_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNIR6CE_0_LC_10_8_4.C_ON=1'b0;
    defparam sEETrigCounter_RNIR6CE_0_LC_10_8_4.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNIR6CE_0_LC_10_8_4.LUT_INIT=16'b0011001100110011;
    LogicCell40 sEETrigCounter_RNIR6CE_0_LC_10_8_4 (
            .in0(_gnd_net_),
            .in1(N__26037),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un10_trig_prev_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigCounter_RNINEOS_1_LC_10_8_6.C_ON=1'b0;
    defparam sEETrigCounter_RNINEOS_1_LC_10_8_6.SEQ_MODE=4'b0000;
    defparam sEETrigCounter_RNINEOS_1_LC_10_8_6.LUT_INIT=16'b1100110000110011;
    LogicCell40 sEETrigCounter_RNINEOS_1_LC_10_8_6 (
            .in0(_gnd_net_),
            .in1(N__26038),
            .in2(_gnd_net_),
            .in3(N__26015),
            .lcout(un10_trig_prev_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_22_0_LC_10_9_0.C_ON=1'b0;
    defparam sDAC_mem_22_0_LC_10_9_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_0_LC_10_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_0_LC_10_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51138),
            .lcout(sDAC_mem_22Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47791),
            .ce(N__39817),
            .sr(N__53039));
    defparam sDAC_mem_22_7_LC_10_9_1.C_ON=1'b0;
    defparam sDAC_mem_22_7_LC_10_9_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_7_LC_10_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_7_LC_10_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48706),
            .lcout(sDAC_mem_22Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47791),
            .ce(N__39817),
            .sr(N__53039));
    defparam \spi_slave_inst.rx_done_reg3_i_LC_10_10_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_reg3_i_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_done_reg3_i_LC_10_10_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.rx_done_reg3_i_LC_10_10_0  (
            .in0(N__28793),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_inst.rx_done_reg3_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47777),
            .ce(),
            .sr(N__53029));
    defparam \spi_slave_inst.rx_ready_i_RNO_0_LC_10_10_1 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_ready_i_RNO_0_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_ready_i_RNO_0_LC_10_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \spi_slave_inst.rx_ready_i_RNO_0_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__26133),
            .in2(_gnd_net_),
            .in3(N__28792),
            .lcout(),
            .ltout(\spi_slave_inst.rx_ready_i_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rx_ready_i_LC_10_10_2 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_ready_i_LC_10_10_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_ready_i_LC_10_10_2 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \spi_slave_inst.rx_ready_i_LC_10_10_2  (
            .in0(N__32466),
            .in1(N__33230),
            .in2(N__26127),
            .in3(N__27314),
            .lcout(spi_mosi_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47777),
            .ce(),
            .sr(N__53029));
    defparam spi_mosi_ready_prev_LC_10_10_3.C_ON=1'b0;
    defparam spi_mosi_ready_prev_LC_10_10_3.SEQ_MODE=4'b1010;
    defparam spi_mosi_ready_prev_LC_10_10_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 spi_mosi_ready_prev_LC_10_10_3 (
            .in0(N__27315),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_mosi_ready_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47777),
            .ce(),
            .sr(N__53029));
    defparam spi_mosi_ready_prev2_LC_10_10_4.C_ON=1'b0;
    defparam spi_mosi_ready_prev2_LC_10_10_4.SEQ_MODE=4'b1010;
    defparam spi_mosi_ready_prev2_LC_10_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 spi_mosi_ready_prev2_LC_10_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26208),
            .lcout(spi_mosi_ready_prevZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47777),
            .ce(),
            .sr(N__53029));
    defparam \spi_slave_inst.tx_ready_i_RNO_0_LC_10_10_5 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_ready_i_RNO_0_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_ready_i_RNO_0_LC_10_10_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \spi_slave_inst.tx_ready_i_RNO_0_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__27090),
            .in2(_gnd_net_),
            .in3(N__27105),
            .lcout(),
            .ltout(\spi_slave_inst.un4_tx_done_reg2_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_ready_i_LC_10_10_6 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_ready_i_LC_10_10_6 .SEQ_MODE=4'b1011;
    defparam \spi_slave_inst.tx_ready_i_LC_10_10_6 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \spi_slave_inst.tx_ready_i_LC_10_10_6  (
            .in0(N__32467),
            .in1(N__33231),
            .in2(N__26124),
            .in3(N__26183),
            .lcout(\spi_slave_inst.tx_ready_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47777),
            .ce(),
            .sr(N__53029));
    defparam spi_mosi_ready_prev3_LC_10_10_7.C_ON=1'b0;
    defparam spi_mosi_ready_prev3_LC_10_10_7.SEQ_MODE=4'b1010;
    defparam spi_mosi_ready_prev3_LC_10_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 spi_mosi_ready_prev3_LC_10_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26220),
            .lcout(spi_mosi_ready_prevZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47777),
            .ce(),
            .sr(N__53029));
    defparam button_debounce_counter_0_LC_10_11_1.C_ON=1'b0;
    defparam button_debounce_counter_0_LC_10_11_1.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_0_LC_10_11_1.LUT_INIT=16'b0101010110101010;
    LogicCell40 button_debounce_counter_0_LC_10_11_1 (
            .in0(N__32468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26298),
            .lcout(button_debounce_counterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53262),
            .ce(),
            .sr(N__26239));
    defparam button_debounce_counter_1_LC_10_11_2.C_ON=1'b0;
    defparam button_debounce_counter_1_LC_10_11_2.SEQ_MODE=4'b1000;
    defparam button_debounce_counter_1_LC_10_11_2.LUT_INIT=16'b0111011110001000;
    LogicCell40 button_debounce_counter_1_LC_10_11_2 (
            .in0(N__26299),
            .in1(N__32469),
            .in2(_gnd_net_),
            .in3(N__26267),
            .lcout(button_debounce_counterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53262),
            .ce(),
            .sr(N__26239));
    defparam spi_mosi_ready_prev3_RNILKER_LC_10_11_4.C_ON=1'b0;
    defparam spi_mosi_ready_prev3_RNILKER_LC_10_11_4.SEQ_MODE=4'b0000;
    defparam spi_mosi_ready_prev3_RNILKER_LC_10_11_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 spi_mosi_ready_prev3_RNILKER_LC_10_11_4 (
            .in0(N__26219),
            .in1(N__26207),
            .in2(N__26196),
            .in3(N__27313),
            .lcout(spi_mosi_ready_prev3_RNILKERZ0),
            .ltout(spi_mosi_ready_prev3_RNILKERZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_rpi_ibuf_RNI7JCV_LC_10_11_5.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNI7JCV_LC_10_11_5.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNI7JCV_LC_10_11_5.LUT_INIT=16'b0101111101011111;
    LogicCell40 reset_rpi_ibuf_RNI7JCV_LC_10_11_5 (
            .in0(N__32470),
            .in1(_gnd_net_),
            .in2(N__26187),
            .in3(_gnd_net_),
            .lcout(reset_rpi_ibuf_RNI7JCVZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_0_LC_10_12_2.C_ON=1'b0;
    defparam sAddress_RNIA6242_0_LC_10_12_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_0_LC_10_12_2.LUT_INIT=16'b0100000000000000;
    LogicCell40 sAddress_RNIA6242_0_LC_10_12_2 (
            .in0(N__31094),
            .in1(N__40395),
            .in2(N__27141),
            .in3(N__44749),
            .lcout(sAddress_RNIA6242Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_ready_i_RNIBLID_LC_10_12_3 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_ready_i_RNIBLID_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_ready_i_RNIBLID_LC_10_12_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \spi_slave_inst.tx_ready_i_RNIBLID_LC_10_12_3  (
            .in0(N__32398),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26184),
            .lcout(\spi_slave_inst.un4_i_wr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sRead_data_RNO_0_LC_10_12_7.C_ON=1'b0;
    defparam sRead_data_RNO_0_LC_10_12_7.SEQ_MODE=4'b0000;
    defparam sRead_data_RNO_0_LC_10_12_7.LUT_INIT=16'b1100110011111111;
    LogicCell40 sRead_data_RNO_0_LC_10_12_7 (
            .in0(_gnd_net_),
            .in1(N__27978),
            .in2(_gnd_net_),
            .in3(N__27882),
            .lcout(N_86),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sADC_clk_prev_LC_10_13_0.C_ON=1'b0;
    defparam sADC_clk_prev_LC_10_13_0.SEQ_MODE=4'b1000;
    defparam sADC_clk_prev_LC_10_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sADC_clk_prev_LC_10_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27621),
            .lcout(sADC_clk_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47792),
            .ce(N__26754),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_0_c_LC_10_14_0.C_ON=1'b1;
    defparam un1_sacqtime_cry_0_c_LC_10_14_0.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_0_c_LC_10_14_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_0_c_LC_10_14_0 (
            .in0(_gnd_net_),
            .in1(N__34154),
            .in2(N__26168),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(un1_sacqtime_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_1_c_LC_10_14_1.C_ON=1'b1;
    defparam un1_sacqtime_cry_1_c_LC_10_14_1.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_1_c_LC_10_14_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_1_c_LC_10_14_1 (
            .in0(_gnd_net_),
            .in1(N__35075),
            .in2(N__26150),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_0),
            .carryout(un1_sacqtime_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_2_c_LC_10_14_2.C_ON=1'b1;
    defparam un1_sacqtime_cry_2_c_LC_10_14_2.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_2_c_LC_10_14_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_2_c_LC_10_14_2 (
            .in0(_gnd_net_),
            .in1(N__34877),
            .in2(N__26459),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_1),
            .carryout(un1_sacqtime_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_3_c_LC_10_14_3.C_ON=1'b1;
    defparam un1_sacqtime_cry_3_c_LC_10_14_3.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_3_c_LC_10_14_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_3_c_LC_10_14_3 (
            .in0(_gnd_net_),
            .in1(N__34772),
            .in2(N__26441),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_2),
            .carryout(un1_sacqtime_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_4_c_LC_10_14_4.C_ON=1'b1;
    defparam un1_sacqtime_cry_4_c_LC_10_14_4.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_4_c_LC_10_14_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_4_c_LC_10_14_4 (
            .in0(_gnd_net_),
            .in1(N__34745),
            .in2(N__26423),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_3),
            .carryout(un1_sacqtime_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_5_c_LC_10_14_5.C_ON=1'b1;
    defparam un1_sacqtime_cry_5_c_LC_10_14_5.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_5_c_LC_10_14_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_5_c_LC_10_14_5 (
            .in0(_gnd_net_),
            .in1(N__34640),
            .in2(N__26405),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_4),
            .carryout(un1_sacqtime_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_6_c_LC_10_14_6.C_ON=1'b1;
    defparam un1_sacqtime_cry_6_c_LC_10_14_6.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_6_c_LC_10_14_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_6_c_LC_10_14_6 (
            .in0(_gnd_net_),
            .in1(N__34514),
            .in2(N__26387),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_5),
            .carryout(un1_sacqtime_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_7_c_LC_10_14_7.C_ON=1'b1;
    defparam un1_sacqtime_cry_7_c_LC_10_14_7.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_7_c_LC_10_14_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_7_c_LC_10_14_7 (
            .in0(_gnd_net_),
            .in1(N__34397),
            .in2(N__26366),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_6),
            .carryout(un1_sacqtime_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_8_c_LC_10_15_0.C_ON=1'b1;
    defparam un1_sacqtime_cry_8_c_LC_10_15_0.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_8_c_LC_10_15_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_8_c_LC_10_15_0 (
            .in0(_gnd_net_),
            .in1(N__35792),
            .in2(N__26348),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(un1_sacqtime_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_9_c_LC_10_15_1.C_ON=1'b1;
    defparam un1_sacqtime_cry_9_c_LC_10_15_1.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_9_c_LC_10_15_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_9_c_LC_10_15_1 (
            .in0(_gnd_net_),
            .in1(N__35681),
            .in2(N__26330),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_8),
            .carryout(un1_sacqtime_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_10_c_LC_10_15_2.C_ON=1'b1;
    defparam un1_sacqtime_cry_10_c_LC_10_15_2.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_10_c_LC_10_15_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_10_c_LC_10_15_2 (
            .in0(_gnd_net_),
            .in1(N__35567),
            .in2(N__26582),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_9),
            .carryout(un1_sacqtime_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_11_c_LC_10_15_3.C_ON=1'b1;
    defparam un1_sacqtime_cry_11_c_LC_10_15_3.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_11_c_LC_10_15_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_11_c_LC_10_15_3 (
            .in0(_gnd_net_),
            .in1(N__35462),
            .in2(N__26564),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_10),
            .carryout(un1_sacqtime_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_12_c_LC_10_15_4.C_ON=1'b1;
    defparam un1_sacqtime_cry_12_c_LC_10_15_4.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_12_c_LC_10_15_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_12_c_LC_10_15_4 (
            .in0(_gnd_net_),
            .in1(N__35435),
            .in2(N__26546),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_11),
            .carryout(un1_sacqtime_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_13_c_LC_10_15_5.C_ON=1'b1;
    defparam un1_sacqtime_cry_13_c_LC_10_15_5.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_13_c_LC_10_15_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_13_c_LC_10_15_5 (
            .in0(_gnd_net_),
            .in1(N__35231),
            .in2(N__26528),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_12),
            .carryout(un1_sacqtime_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_14_c_LC_10_15_6.C_ON=1'b1;
    defparam un1_sacqtime_cry_14_c_LC_10_15_6.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_14_c_LC_10_15_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_14_c_LC_10_15_6 (
            .in0(_gnd_net_),
            .in1(N__35111),
            .in2(N__26510),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_13),
            .carryout(un1_sacqtime_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_15_c_LC_10_15_7.C_ON=1'b1;
    defparam un1_sacqtime_cry_15_c_LC_10_15_7.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_15_c_LC_10_15_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_sacqtime_cry_15_c_LC_10_15_7 (
            .in0(_gnd_net_),
            .in1(N__36569),
            .in2(N__26493),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_sacqtime_cry_14),
            .carryout(un1_sacqtime_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_16_c_inv_LC_10_16_0.C_ON=1'b1;
    defparam un1_sacqtime_cry_16_c_inv_LC_10_16_0.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_16_c_inv_LC_10_16_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_sacqtime_cry_16_c_inv_LC_10_16_0 (
            .in0(N__36517),
            .in1(_gnd_net_),
            .in2(N__26478),
            .in3(_gnd_net_),
            .lcout(un1_sacqtime_cry_16_sf),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(un1_sacqtime_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_17_c_inv_LC_10_16_1.C_ON=1'b1;
    defparam un1_sacqtime_cry_17_c_inv_LC_10_16_1.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_17_c_inv_LC_10_16_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_sacqtime_cry_17_c_inv_LC_10_16_1 (
            .in0(N__36416),
            .in1(_gnd_net_),
            .in2(N__26469),
            .in3(_gnd_net_),
            .lcout(un1_sacqtime_cry_17_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_16),
            .carryout(un1_sacqtime_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_18_c_inv_LC_10_16_2.C_ON=1'b1;
    defparam un1_sacqtime_cry_18_c_inv_LC_10_16_2.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_18_c_inv_LC_10_16_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_sacqtime_cry_18_c_inv_LC_10_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26703),
            .in3(N__36323),
            .lcout(un1_sacqtime_cry_18_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_17),
            .carryout(un1_sacqtime_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_19_c_inv_LC_10_16_3.C_ON=1'b1;
    defparam un1_sacqtime_cry_19_c_inv_LC_10_16_3.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_19_c_inv_LC_10_16_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_sacqtime_cry_19_c_inv_LC_10_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26694),
            .in3(N__36231),
            .lcout(un1_sacqtime_cry_19_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_18),
            .carryout(un1_sacqtime_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_20_c_inv_LC_10_16_4.C_ON=1'b1;
    defparam un1_sacqtime_cry_20_c_inv_LC_10_16_4.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_20_c_inv_LC_10_16_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_sacqtime_cry_20_c_inv_LC_10_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26685),
            .in3(N__36146),
            .lcout(un1_sacqtime_cry_20_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_19),
            .carryout(un1_sacqtime_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_21_c_inv_LC_10_16_5.C_ON=1'b1;
    defparam un1_sacqtime_cry_21_c_inv_LC_10_16_5.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_21_c_inv_LC_10_16_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_sacqtime_cry_21_c_inv_LC_10_16_5 (
            .in0(N__36063),
            .in1(_gnd_net_),
            .in2(N__26676),
            .in3(_gnd_net_),
            .lcout(un1_sacqtime_cry_21_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_20),
            .carryout(un1_sacqtime_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_22_c_inv_LC_10_16_6.C_ON=1'b1;
    defparam un1_sacqtime_cry_22_c_inv_LC_10_16_6.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_22_c_inv_LC_10_16_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_sacqtime_cry_22_c_inv_LC_10_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26667),
            .in3(N__35960),
            .lcout(un1_sacqtime_cry_22_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_21),
            .carryout(un1_sacqtime_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_23_c_inv_LC_10_16_7.C_ON=1'b1;
    defparam un1_sacqtime_cry_23_c_inv_LC_10_16_7.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_23_c_inv_LC_10_16_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_sacqtime_cry_23_c_inv_LC_10_16_7 (
            .in0(N__37058),
            .in1(_gnd_net_),
            .in2(N__26658),
            .in3(_gnd_net_),
            .lcout(un1_sacqtime_cry_23_sf),
            .ltout(),
            .carryin(un1_sacqtime_cry_22),
            .carryout(un1_sacqtime_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_sacqtime_cry_23_THRU_LUT4_0_LC_10_17_0.C_ON=1'b0;
    defparam un1_sacqtime_cry_23_THRU_LUT4_0_LC_10_17_0.SEQ_MODE=4'b0000;
    defparam un1_sacqtime_cry_23_THRU_LUT4_0_LC_10_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_sacqtime_cry_23_THRU_LUT4_0_LC_10_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26649),
            .lcout(un1_sacqtime_cry_23_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_10_RNO_0_15_LC_10_17_1.C_ON=1'b0;
    defparam RAM_DATA_cl_10_RNO_0_15_LC_10_17_1.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_10_RNO_0_15_LC_10_17_1.LUT_INIT=16'b0101010100000000;
    LogicCell40 RAM_DATA_cl_10_RNO_0_15_LC_10_17_1 (
            .in0(N__26627),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31670),
            .lcout(N_106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPointerReset_RNI2CQM_LC_10_17_3.C_ON=1'b0;
    defparam sEEPointerReset_RNI2CQM_LC_10_17_3.SEQ_MODE=4'b0000;
    defparam sEEPointerReset_RNI2CQM_LC_10_17_3.LUT_INIT=16'b1011101010101010;
    LogicCell40 sEEPointerReset_RNI2CQM_LC_10_17_3 (
            .in0(N__33475),
            .in1(N__31669),
            .in2(N__32178),
            .in3(N__31847),
            .lcout(N_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sADC_clk_prev_RNO_LC_10_17_4.C_ON=1'b0;
    defparam sADC_clk_prev_RNO_LC_10_17_4.SEQ_MODE=4'b0000;
    defparam sADC_clk_prev_RNO_LC_10_17_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 sADC_clk_prev_RNO_LC_10_17_4 (
            .in0(N__31848),
            .in1(N__32102),
            .in2(_gnd_net_),
            .in3(N__32413),
            .lcout(N_76_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sADC_clk_prev_RNI4BVG_LC_10_17_5.C_ON=1'b0;
    defparam sADC_clk_prev_RNI4BVG_LC_10_17_5.SEQ_MODE=4'b0000;
    defparam sADC_clk_prev_RNI4BVG_LC_10_17_5.LUT_INIT=16'b1010101011111111;
    LogicCell40 sADC_clk_prev_RNI4BVG_LC_10_17_5 (
            .in0(N__27636),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27606),
            .lcout(N_71),
            .ltout(N_71_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_15_RNO_0_15_LC_10_17_6.C_ON=1'b0;
    defparam RAM_DATA_cl_15_RNO_0_15_LC_10_17_6.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_15_RNO_0_15_LC_10_17_6.LUT_INIT=16'b0000000011110000;
    LogicCell40 RAM_DATA_cl_15_RNO_0_15_LC_10_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26742),
            .in3(N__28352),
            .lcout(N_102),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEDelayACQ_0_LC_10_18_0.C_ON=1'b0;
    defparam sEEDelayACQ_0_LC_10_18_0.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_0_LC_10_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_0_LC_10_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51266),
            .lcout(sEEDelayACQZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__27219),
            .sr(N__52979));
    defparam sEEDelayACQ_1_LC_10_18_1.C_ON=1'b0;
    defparam sEEDelayACQ_1_LC_10_18_1.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_1_LC_10_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_1_LC_10_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50769),
            .lcout(sEEDelayACQZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__27219),
            .sr(N__52979));
    defparam sEEDelayACQ_2_LC_10_18_2.C_ON=1'b0;
    defparam sEEDelayACQ_2_LC_10_18_2.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_2_LC_10_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_2_LC_10_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50305),
            .lcout(sEEDelayACQZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__27219),
            .sr(N__52979));
    defparam sEEDelayACQ_3_LC_10_18_3.C_ON=1'b0;
    defparam sEEDelayACQ_3_LC_10_18_3.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_3_LC_10_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_3_LC_10_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49834),
            .lcout(sEEDelayACQZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__27219),
            .sr(N__52979));
    defparam sEEDelayACQ_4_LC_10_18_4.C_ON=1'b0;
    defparam sEEDelayACQ_4_LC_10_18_4.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_4_LC_10_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_4_LC_10_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49306),
            .lcout(sEEDelayACQZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__27219),
            .sr(N__52979));
    defparam sEEDelayACQ_5_LC_10_18_5.C_ON=1'b0;
    defparam sEEDelayACQ_5_LC_10_18_5.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_5_LC_10_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_5_LC_10_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47130),
            .lcout(sEEDelayACQZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__27219),
            .sr(N__52979));
    defparam sEEDelayACQ_6_LC_10_18_6.C_ON=1'b0;
    defparam sEEDelayACQ_6_LC_10_18_6.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_6_LC_10_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_6_LC_10_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48230),
            .lcout(sEEDelayACQZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__27219),
            .sr(N__52979));
    defparam sEEDelayACQ_7_LC_10_18_7.C_ON=1'b0;
    defparam sEEDelayACQ_7_LC_10_18_7.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_7_LC_10_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_7_LC_10_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48832),
            .lcout(sEEDelayACQZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47839),
            .ce(N__27219),
            .sr(N__52979));
    defparam sEEDelayACQ_10_LC_10_19_0.C_ON=1'b0;
    defparam sEEDelayACQ_10_LC_10_19_0.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_10_LC_10_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_10_LC_10_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50306),
            .lcout(sEEDelayACQZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(N__26946),
            .sr(N__52975));
    defparam sEEDelayACQ_11_LC_10_19_1.C_ON=1'b0;
    defparam sEEDelayACQ_11_LC_10_19_1.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_11_LC_10_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_11_LC_10_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49790),
            .lcout(sEEDelayACQZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(N__26946),
            .sr(N__52975));
    defparam sEEDelayACQ_12_LC_10_19_2.C_ON=1'b0;
    defparam sEEDelayACQ_12_LC_10_19_2.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_12_LC_10_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_12_LC_10_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49189),
            .lcout(sEEDelayACQZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(N__26946),
            .sr(N__52975));
    defparam sEEDelayACQ_13_LC_10_19_3.C_ON=1'b0;
    defparam sEEDelayACQ_13_LC_10_19_3.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_13_LC_10_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_13_LC_10_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47149),
            .lcout(sEEDelayACQZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(N__26946),
            .sr(N__52975));
    defparam sEEDelayACQ_14_LC_10_19_4.C_ON=1'b0;
    defparam sEEDelayACQ_14_LC_10_19_4.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_14_LC_10_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_14_LC_10_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48231),
            .lcout(sEEDelayACQZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(N__26946),
            .sr(N__52975));
    defparam sEEDelayACQ_15_LC_10_19_5.C_ON=1'b0;
    defparam sEEDelayACQ_15_LC_10_19_5.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_15_LC_10_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDelayACQ_15_LC_10_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48768),
            .lcout(sEEDelayACQZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(N__26946),
            .sr(N__52975));
    defparam sEEDelayACQ_8_LC_10_19_6.C_ON=1'b0;
    defparam sEEDelayACQ_8_LC_10_19_6.SEQ_MODE=4'b1010;
    defparam sEEDelayACQ_8_LC_10_19_6.LUT_INIT=16'b1100110011001100;
    LogicCell40 sEEDelayACQ_8_LC_10_19_6 (
            .in0(_gnd_net_),
            .in1(N__51267),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(N__26946),
            .sr(N__52975));
    defparam sEEDelayACQ_9_LC_10_19_7.C_ON=1'b0;
    defparam sEEDelayACQ_9_LC_10_19_7.SEQ_MODE=4'b1011;
    defparam sEEDelayACQ_9_LC_10_19_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 sEEDelayACQ_9_LC_10_19_7 (
            .in0(_gnd_net_),
            .in1(N__50770),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEDelayACQZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47847),
            .ce(N__26946),
            .sr(N__52975));
    defparam RAM_DATA_cl_12_RNO_0_15_LC_10_20_1.C_ON=1'b0;
    defparam RAM_DATA_cl_12_RNO_0_15_LC_10_20_1.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_12_RNO_0_15_LC_10_20_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 RAM_DATA_cl_12_RNO_0_15_LC_10_20_1 (
            .in0(_gnd_net_),
            .in1(N__26912),
            .in2(_gnd_net_),
            .in3(N__31708),
            .lcout(),
            .ltout(N_99_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_12_15_LC_10_20_2.C_ON=1'b0;
    defparam RAM_DATA_cl_12_15_LC_10_20_2.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_12_15_LC_10_20_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 RAM_DATA_cl_12_15_LC_10_20_2 (
            .in0(N__32502),
            .in1(N__32067),
            .in2(N__26934),
            .in3(N__31968),
            .lcout(RAM_DATA_cl_12Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47851),
            .ce(),
            .sr(N__52971));
    defparam RAM_DATA_cl_11_RNO_0_15_LC_10_20_3.C_ON=1'b0;
    defparam RAM_DATA_cl_11_RNO_0_15_LC_10_20_3.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_11_RNO_0_15_LC_10_20_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 RAM_DATA_cl_11_RNO_0_15_LC_10_20_3 (
            .in0(_gnd_net_),
            .in1(N__26879),
            .in2(_gnd_net_),
            .in3(N__31707),
            .lcout(),
            .ltout(N_94_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_11_15_LC_10_20_4.C_ON=1'b0;
    defparam RAM_DATA_cl_11_15_LC_10_20_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_11_15_LC_10_20_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 RAM_DATA_cl_11_15_LC_10_20_4 (
            .in0(N__32501),
            .in1(N__32066),
            .in2(N__26901),
            .in3(N__31967),
            .lcout(RAM_DATA_cl_11Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47851),
            .ce(),
            .sr(N__52971));
    defparam RAM_DATA_cl_14_RNO_0_15_LC_10_20_5.C_ON=1'b0;
    defparam RAM_DATA_cl_14_RNO_0_15_LC_10_20_5.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_14_RNO_0_15_LC_10_20_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 RAM_DATA_cl_14_RNO_0_15_LC_10_20_5 (
            .in0(_gnd_net_),
            .in1(N__26852),
            .in2(_gnd_net_),
            .in3(N__31709),
            .lcout(),
            .ltout(N_104_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_14_15_LC_10_20_6.C_ON=1'b0;
    defparam RAM_DATA_cl_14_15_LC_10_20_6.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_14_15_LC_10_20_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 RAM_DATA_cl_14_15_LC_10_20_6 (
            .in0(N__32503),
            .in1(N__32068),
            .in2(N__26868),
            .in3(N__31969),
            .lcout(RAM_DATA_cl_14Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47851),
            .ce(),
            .sr(N__52971));
    defparam sDAC_data_2_LC_11_2_1.C_ON=1'b0;
    defparam sDAC_data_2_LC_11_2_1.SEQ_MODE=4'b1010;
    defparam sDAC_data_2_LC_11_2_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_2_LC_11_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53243),
            .ce(N__42234),
            .sr(N__53109));
    defparam \spi_slave_inst.rx_done_neg_sclk_i_LC_11_3_7 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_neg_sclk_i_LC_11_3_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_done_neg_sclk_i_LC_11_3_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \spi_slave_inst.rx_done_neg_sclk_i_LC_11_3_7  (
            .in0(N__27065),
            .in1(N__33194),
            .in2(_gnd_net_),
            .in3(N__26829),
            .lcout(\spi_slave_inst.rx_done_neg_sclk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVspi_slave_inst.rx_done_neg_sclk_iC_net ),
            .ce(),
            .sr(N__53096));
    defparam \spi_slave_inst.rx_done_reg1_i_LC_11_4_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_reg1_i_LC_11_4_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_done_reg1_i_LC_11_4_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \spi_slave_inst.rx_done_reg1_i_LC_11_4_0  (
            .in0(N__27066),
            .in1(N__33214),
            .in2(_gnd_net_),
            .in3(N__27054),
            .lcout(\spi_slave_inst.rx_done_reg1_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47832),
            .ce(),
            .sr(N__53083));
    defparam \spi_slave_inst.txdata_reg_i_5_LC_11_4_2 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_5_LC_11_4_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_5_LC_11_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_5_LC_11_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27378),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47832),
            .ce(),
            .sr(N__53083));
    defparam \spi_slave_inst.txdata_reg_i_4_LC_11_4_7 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_4_LC_11_4_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_4_LC_11_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_4_LC_11_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27237),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47832),
            .ce(),
            .sr(N__53083));
    defparam \spi_master_inst.spi_data_path_u1.tx_ready_i_LC_11_5_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_ready_i_LC_11_5_0 .SEQ_MODE=4'b1011;
    defparam \spi_master_inst.spi_data_path_u1.tx_ready_i_LC_11_5_0 .LUT_INIT=16'b0000000011110100;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_ready_i_LC_11_5_0  (
            .in0(N__27048),
            .in1(N__27041),
            .in2(N__28837),
            .in3(N__47306),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_ready_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53245),
            .ce(),
            .sr(N__53071));
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg3_i_LC_11_5_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg3_i_LC_11_5_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg3_i_LC_11_5_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_done_reg3_i_LC_11_5_1  (
            .in0(N__27042),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_done_reg3_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53245),
            .ce(),
            .sr(N__53071));
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg2_i_LC_11_5_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg2_i_LC_11_5_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg2_i_LC_11_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_done_reg2_i_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27009),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_done_reg2_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53245),
            .ce(),
            .sr(N__53071));
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg1_i_LC_11_5_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg1_i_LC_11_5_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.tx_done_reg1_i_LC_11_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.tx_done_reg1_i_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27033),
            .lcout(\spi_master_inst.spi_data_path_u1.tx_done_reg1_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53245),
            .ce(),
            .sr(N__53071));
    defparam \spi_master_inst.sclk_gen_u0.spi_start_i_LC_11_5_4 .C_ON=1'b0;
    defparam \spi_master_inst.sclk_gen_u0.spi_start_i_LC_11_5_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.sclk_gen_u0.spi_start_i_LC_11_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.sclk_gen_u0.spi_start_i_LC_11_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47307),
            .lcout(\spi_master_inst.sclk_gen_u0.spi_start_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53245),
            .ce(),
            .sr(N__53071));
    defparam \spi_slave_inst.txdata_reg_i_RNI1IQC_0_LC_11_5_7 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_RNI1IQC_0_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.txdata_reg_i_RNI1IQC_0_LC_11_5_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi_slave_inst.txdata_reg_i_RNI1IQC_0_LC_11_5_7  (
            .in0(N__37153),
            .in1(N__26958),
            .in2(_gnd_net_),
            .in3(N__27078),
            .lcout(\spi_slave_inst.txdata_reg_i_RNI1IQCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.txdata_reg_i_RNI7OQC_3_LC_11_6_2 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_RNI7OQC_3_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.txdata_reg_i_RNI7OQC_3_LC_11_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi_slave_inst.txdata_reg_i_RNI7OQC_3_LC_11_6_2  (
            .in0(N__27204),
            .in1(N__27195),
            .in2(_gnd_net_),
            .in3(N__37162),
            .lcout(),
            .ltout(\spi_slave_inst.txdata_reg_i_RNI7OQCZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIUCSS_1_LC_11_6_3 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIUCSS_1_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIUCSS_1_LC_11_6_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNIUCSS_1_LC_11_6_3  (
            .in0(N__27177),
            .in1(_gnd_net_),
            .in2(N__27129),
            .in3(N__37221),
            .lcout(\spi_slave_inst.N_1394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ8SS_1_LC_11_6_5 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ8SS_1_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ8SS_1_LC_11_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ8SS_1_LC_11_6_5  (
            .in0(N__27162),
            .in1(N__27126),
            .in2(_gnd_net_),
            .in3(N__37220),
            .lcout(),
            .ltout(\spi_slave_inst.N_1397_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIA0LM2_0_LC_11_6_6 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIA0LM2_0_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIA0LM2_0_LC_11_6_6 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNIA0LM2_0_LC_11_6_6  (
            .in0(N__33224),
            .in1(N__27120),
            .in2(N__27114),
            .in3(N__37251),
            .lcout(\spi_slave_inst.spi_miso ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_23_7_LC_11_7_7.C_ON=1'b0;
    defparam sDAC_mem_23_7_LC_11_7_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_7_LC_11_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_7_LC_11_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48599),
            .lcout(sDAC_mem_23Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47804),
            .ce(N__28989),
            .sr(N__53049));
    defparam sPointer_1_LC_11_8_0.C_ON=1'b0;
    defparam sPointer_1_LC_11_8_0.SEQ_MODE=4'b1010;
    defparam sPointer_1_LC_11_8_0.LUT_INIT=16'b0110011001000100;
    LogicCell40 sPointer_1_LC_11_8_0 (
            .in0(N__29217),
            .in1(N__43832),
            .in2(_gnd_net_),
            .in3(N__29189),
            .lcout(sPointerZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47793),
            .ce(),
            .sr(N__53040));
    defparam \spi_slave_inst.tx_done_reg1_i_LC_11_8_1 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_done_reg1_i_LC_11_8_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_done_reg1_i_LC_11_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.tx_done_reg1_i_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33159),
            .lcout(\spi_slave_inst.tx_done_reg1_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47793),
            .ce(),
            .sr(N__53040));
    defparam \spi_slave_inst.tx_done_reg2_i_LC_11_8_2 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_done_reg2_i_LC_11_8_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_done_reg2_i_LC_11_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.tx_done_reg2_i_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27111),
            .lcout(\spi_slave_inst.tx_done_reg2_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47793),
            .ce(),
            .sr(N__53040));
    defparam \spi_slave_inst.tx_done_reg3_i_LC_11_8_3 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_done_reg3_i_LC_11_8_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_done_reg3_i_LC_11_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.tx_done_reg3_i_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27104),
            .lcout(\spi_slave_inst.tx_done_reg3_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47793),
            .ce(),
            .sr(N__53040));
    defparam \spi_slave_inst.txdata_reg_i_0_LC_11_8_4 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_0_LC_11_8_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_0_LC_11_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_0_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27273),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47793),
            .ce(),
            .sr(N__53040));
    defparam \spi_slave_inst.txdata_reg_i_3_LC_11_8_5 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_3_LC_11_8_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_3_LC_11_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_3_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27246),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47793),
            .ce(),
            .sr(N__53040));
    defparam \spi_slave_inst.txdata_reg_i_7_LC_11_8_7 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_7_LC_11_8_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_7_LC_11_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.txdata_reg_i_7_LC_11_8_7  (
            .in0(N__27357),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47793),
            .ce(),
            .sr(N__53040));
    defparam \spi_slave_inst.txdata_reg_i_RNI3KQC_1_LC_11_9_0 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_RNI3KQC_1_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.txdata_reg_i_RNI3KQC_1_LC_11_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \spi_slave_inst.txdata_reg_i_RNI3KQC_1_LC_11_9_0  (
            .in0(N__27168),
            .in1(N__27186),
            .in2(_gnd_net_),
            .in3(N__37163),
            .lcout(\spi_slave_inst.txdata_reg_i_RNI3KQCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.txdata_reg_i_1_LC_11_9_1 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_1_LC_11_9_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_1_LC_11_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_1_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27264),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47778),
            .ce(),
            .sr(N__53030));
    defparam \spi_slave_inst.txdata_reg_i_RNI5MQC_2_LC_11_9_3 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_RNI5MQC_2_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.txdata_reg_i_RNI5MQC_2_LC_11_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \spi_slave_inst.txdata_reg_i_RNI5MQC_2_LC_11_9_3  (
            .in0(N__37164),
            .in1(N__27147),
            .in2(_gnd_net_),
            .in3(N__27153),
            .lcout(\spi_slave_inst.txdata_reg_i_RNI5MQCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.txdata_reg_i_2_LC_11_9_4 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_2_LC_11_9_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_2_LC_11_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_2_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27255),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47778),
            .ce(),
            .sr(N__53030));
    defparam \spi_slave_inst.txdata_reg_i_6_LC_11_9_5 .C_ON=1'b0;
    defparam \spi_slave_inst.txdata_reg_i_6_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.txdata_reg_i_6_LC_11_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.txdata_reg_i_6_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27366),
            .lcout(\spi_slave_inst.txdata_reg_iZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47778),
            .ce(),
            .sr(N__53030));
    defparam sPointer_0_LC_11_9_7.C_ON=1'b0;
    defparam sPointer_0_LC_11_9_7.SEQ_MODE=4'b1010;
    defparam sPointer_0_LC_11_9_7.LUT_INIT=16'b0001000110101010;
    LogicCell40 sPointer_0_LC_11_9_7 (
            .in0(N__29188),
            .in1(N__43833),
            .in2(_gnd_net_),
            .in3(N__29213),
            .lcout(sPointerZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47778),
            .ce(),
            .sr(N__53030));
    defparam sAddress_RNIAM2A_0_1_LC_11_10_1.C_ON=1'b0;
    defparam sAddress_RNIAM2A_0_1_LC_11_10_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNIAM2A_0_1_LC_11_10_1.LUT_INIT=16'b0000010000000010;
    LogicCell40 sAddress_RNIAM2A_0_1_LC_11_10_1 (
            .in0(N__44952),
            .in1(N__40326),
            .in2(N__40538),
            .in3(N__44869),
            .lcout(N_206),
            .ltout(N_206_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_1_0_LC_11_10_2.C_ON=1'b0;
    defparam sAddress_RNIA6242_1_0_LC_11_10_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_1_0_LC_11_10_2.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNIA6242_1_0_LC_11_10_2 (
            .in0(N__40327),
            .in1(N__31072),
            .in2(N__27222),
            .in3(N__44718),
            .lcout(sAddress_RNIA6242_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIQ63A_6_LC_11_10_3.C_ON=1'b0;
    defparam sAddress_RNIQ63A_6_LC_11_10_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNIQ63A_6_LC_11_10_3.LUT_INIT=16'b1111111101111111;
    LogicCell40 sAddress_RNIQ63A_6_LC_11_10_3 (
            .in0(N__30946),
            .in1(N__46485),
            .in2(N__30926),
            .in3(N__44613),
            .lcout(N_141),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_4_LC_11_10_4.C_ON=1'b0;
    defparam sAddress_4_LC_11_10_4.SEQ_MODE=4'b1010;
    defparam sAddress_4_LC_11_10_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 sAddress_4_LC_11_10_4 (
            .in0(_gnd_net_),
            .in1(N__49230),
            .in2(_gnd_net_),
            .in3(N__43843),
            .lcout(sAddressZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47764),
            .ce(N__43775),
            .sr(N__53020));
    defparam sAddress_6_LC_11_10_5.C_ON=1'b0;
    defparam sAddress_6_LC_11_10_5.SEQ_MODE=4'b1010;
    defparam sAddress_6_LC_11_10_5.LUT_INIT=16'b0101010100000000;
    LogicCell40 sAddress_6_LC_11_10_5 (
            .in0(N__43844),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48159),
            .lcout(sAddressZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47764),
            .ce(N__43775),
            .sr(N__53020));
    defparam sAddress_RNIFL15_6_LC_11_10_6.C_ON=1'b0;
    defparam sAddress_RNIFL15_6_LC_11_10_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNIFL15_6_LC_11_10_6.LUT_INIT=16'b0000000000110011;
    LogicCell40 sAddress_RNIFL15_6_LC_11_10_6 (
            .in0(_gnd_net_),
            .in1(N__30922),
            .in2(_gnd_net_),
            .in3(N__30947),
            .lcout(sDAC_mem_30_1_sqmuxa_0_a2_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_7_LC_11_10_7.C_ON=1'b0;
    defparam sAddress_7_LC_11_10_7.SEQ_MODE=4'b1010;
    defparam sAddress_7_LC_11_10_7.LUT_INIT=16'b0101010100000000;
    LogicCell40 sAddress_7_LC_11_10_7 (
            .in0(N__43845),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48592),
            .lcout(sAddressZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47764),
            .ce(N__43775),
            .sr(N__53020));
    defparam sEEPointerReset_RNO_1_LC_11_11_0.C_ON=1'b0;
    defparam sEEPointerReset_RNO_1_LC_11_11_0.SEQ_MODE=4'b0000;
    defparam sEEPointerReset_RNO_1_LC_11_11_0.LUT_INIT=16'b0100000000000000;
    LogicCell40 sEEPointerReset_RNO_1_LC_11_11_0 (
            .in0(N__43846),
            .in1(N__29191),
            .in2(N__32554),
            .in3(N__29128),
            .lcout(N_269),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sPointer_RNIPU81_0_LC_11_11_1.C_ON=1'b0;
    defparam sPointer_RNIPU81_0_LC_11_11_1.SEQ_MODE=4'b0000;
    defparam sPointer_RNIPU81_0_LC_11_11_1.LUT_INIT=16'b1111111111001100;
    LogicCell40 sPointer_RNIPU81_0_LC_11_11_1 (
            .in0(_gnd_net_),
            .in1(N__29190),
            .in2(_gnd_net_),
            .in3(N__43847),
            .lcout(N_159),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam spi_mosi_ready64_prev_e_0_LC_11_11_2.C_ON=1'b0;
    defparam spi_mosi_ready64_prev_e_0_LC_11_11_2.SEQ_MODE=4'b1000;
    defparam spi_mosi_ready64_prev_e_0_LC_11_11_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 spi_mosi_ready64_prev_e_0_LC_11_11_2 (
            .in0(N__27312),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_mosi_ready64_prevZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47754),
            .ce(N__32515),
            .sr(_gnd_net_));
    defparam spi_mosi_ready64_prev3_e_0_LC_11_11_3.C_ON=1'b0;
    defparam spi_mosi_ready64_prev3_e_0_LC_11_11_3.SEQ_MODE=4'b1000;
    defparam spi_mosi_ready64_prev3_e_0_LC_11_11_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 spi_mosi_ready64_prev3_e_0_LC_11_11_3 (
            .in0(N__27342),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_mosi_ready64_prevZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47754),
            .ce(N__32515),
            .sr(_gnd_net_));
    defparam spi_mosi_ready64_prev2_e_0_LC_11_11_4.C_ON=1'b0;
    defparam spi_mosi_ready64_prev2_e_0_LC_11_11_4.SEQ_MODE=4'b1000;
    defparam spi_mosi_ready64_prev2_e_0_LC_11_11_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 spi_mosi_ready64_prev2_e_0_LC_11_11_4 (
            .in0(N__27333),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_mosi_ready64_prevZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47754),
            .ce(N__32515),
            .sr(_gnd_net_));
    defparam spi_mosi_ready64_prev3_e_0_RNICM2C1_LC_11_11_5.C_ON=1'b0;
    defparam spi_mosi_ready64_prev3_e_0_RNICM2C1_LC_11_11_5.SEQ_MODE=4'b0000;
    defparam spi_mosi_ready64_prev3_e_0_RNICM2C1_LC_11_11_5.LUT_INIT=16'b0000100000000000;
    LogicCell40 spi_mosi_ready64_prev3_e_0_RNICM2C1_LC_11_11_5 (
            .in0(N__27341),
            .in1(N__27332),
            .in2(N__27324),
            .in3(N__27311),
            .lcout(spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1),
            .ltout(spi_mosi_ready64_prev3_e_0_RNICM2CZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sPointer_RNI85NC1_0_LC_11_11_6.C_ON=1'b0;
    defparam sPointer_RNI85NC1_0_LC_11_11_6.SEQ_MODE=4'b0000;
    defparam sPointer_RNI85NC1_0_LC_11_11_6.LUT_INIT=16'b1111000000000000;
    LogicCell40 sPointer_RNI85NC1_0_LC_11_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27291),
            .in3(N__29192),
            .lcout(un1_spointer11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_rpi_ibuf_RNIIUT3_LC_11_11_7.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNIIUT3_LC_11_11_7.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNIIUT3_LC_11_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 reset_rpi_ibuf_RNIIUT3_LC_11_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32516),
            .lcout(LED3_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.data_in_reg_i_0_LC_11_12_0 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_0_LC_11_12_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_0_LC_11_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_0_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29526),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47765),
            .ce(N__27348),
            .sr(N__53009));
    defparam \spi_slave_inst.data_in_reg_i_1_LC_11_12_1 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_1_LC_11_12_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_1_LC_11_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_1_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29481),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47765),
            .ce(N__27348),
            .sr(N__53009));
    defparam \spi_slave_inst.data_in_reg_i_2_LC_11_12_2 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_2_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_2_LC_11_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_2_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29421),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47765),
            .ce(N__27348),
            .sr(N__53009));
    defparam \spi_slave_inst.data_in_reg_i_3_LC_11_12_3 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_3_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_3_LC_11_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_3_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30009),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47765),
            .ce(N__27348),
            .sr(N__53009));
    defparam \spi_slave_inst.data_in_reg_i_4_LC_11_12_4 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_4_LC_11_12_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_4_LC_11_12_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.data_in_reg_i_4_LC_11_12_4  (
            .in0(N__29952),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47765),
            .ce(N__27348),
            .sr(N__53009));
    defparam \spi_slave_inst.data_in_reg_i_5_LC_11_12_5 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_5_LC_11_12_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_5_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_5_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29799),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47765),
            .ce(N__27348),
            .sr(N__53009));
    defparam \spi_slave_inst.data_in_reg_i_6_LC_11_12_6 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_6_LC_11_12_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_6_LC_11_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_6_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27720),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47765),
            .ce(N__27348),
            .sr(N__53009));
    defparam \spi_slave_inst.data_in_reg_i_7_LC_11_12_7 .C_ON=1'b0;
    defparam \spi_slave_inst.data_in_reg_i_7_LC_11_12_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.data_in_reg_i_7_LC_11_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.data_in_reg_i_7_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27669),
            .lcout(\spi_slave_inst.data_in_reg_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47765),
            .ce(N__27348),
            .sr(N__53009));
    defparam sEEACQ_0_LC_11_13_0.C_ON=1'b0;
    defparam sEEACQ_0_LC_11_13_0.SEQ_MODE=4'b1010;
    defparam sEEACQ_0_LC_11_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_0_LC_11_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51080),
            .lcout(sEEACQZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47779),
            .ce(N__28911),
            .sr(N__53001));
    defparam sEEACQ_1_LC_11_13_1.C_ON=1'b0;
    defparam sEEACQ_1_LC_11_13_1.SEQ_MODE=4'b1010;
    defparam sEEACQ_1_LC_11_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_1_LC_11_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50664),
            .lcout(sEEACQZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47779),
            .ce(N__28911),
            .sr(N__53001));
    defparam sEEACQ_2_LC_11_13_2.C_ON=1'b0;
    defparam sEEACQ_2_LC_11_13_2.SEQ_MODE=4'b1010;
    defparam sEEACQ_2_LC_11_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_2_LC_11_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50274),
            .lcout(sEEACQZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47779),
            .ce(N__28911),
            .sr(N__53001));
    defparam sEEACQ_3_LC_11_13_3.C_ON=1'b0;
    defparam sEEACQ_3_LC_11_13_3.SEQ_MODE=4'b1011;
    defparam sEEACQ_3_LC_11_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_3_LC_11_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49689),
            .lcout(sEEACQZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47779),
            .ce(N__28911),
            .sr(N__53001));
    defparam sEEACQ_4_LC_11_13_4.C_ON=1'b0;
    defparam sEEACQ_4_LC_11_13_4.SEQ_MODE=4'b1010;
    defparam sEEACQ_4_LC_11_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_4_LC_11_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49368),
            .lcout(sEEACQZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47779),
            .ce(N__28911),
            .sr(N__53001));
    defparam sEEACQ_5_LC_11_13_5.C_ON=1'b0;
    defparam sEEACQ_5_LC_11_13_5.SEQ_MODE=4'b1010;
    defparam sEEACQ_5_LC_11_13_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEACQ_5_LC_11_13_5 (
            .in0(N__47046),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEACQZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47779),
            .ce(N__28911),
            .sr(N__53001));
    defparam sEEACQ_6_LC_11_13_6.C_ON=1'b0;
    defparam sEEACQ_6_LC_11_13_6.SEQ_MODE=4'b1011;
    defparam sEEACQ_6_LC_11_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_6_LC_11_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48274),
            .lcout(sEEACQZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47779),
            .ce(N__28911),
            .sr(N__53001));
    defparam sEEACQ_7_LC_11_13_7.C_ON=1'b0;
    defparam sEEACQ_7_LC_11_13_7.SEQ_MODE=4'b1011;
    defparam sEEACQ_7_LC_11_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_7_LC_11_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48705),
            .lcout(sEEACQZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47779),
            .ce(N__28911),
            .sr(N__53001));
    defparam spi_data_miso_6_LC_11_14_0.C_ON=1'b0;
    defparam spi_data_miso_6_LC_11_14_0.SEQ_MODE=4'b1010;
    defparam spi_data_miso_6_LC_11_14_0.LUT_INIT=16'b0000000010111000;
    LogicCell40 spi_data_miso_6_LC_11_14_0 (
            .in0(N__27765),
            .in1(N__29852),
            .in2(N__27741),
            .in3(N__29937),
            .lcout(spi_data_misoZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47794),
            .ce(N__29780),
            .sr(N__52992));
    defparam spi_data_miso_7_LC_11_14_1.C_ON=1'b0;
    defparam spi_data_miso_7_LC_11_14_1.SEQ_MODE=4'b1010;
    defparam spi_data_miso_7_LC_11_14_1.LUT_INIT=16'b1110111111101010;
    LogicCell40 spi_data_miso_7_LC_11_14_1 (
            .in0(N__29938),
            .in1(N__27711),
            .in2(N__29868),
            .in3(N__27687),
            .lcout(spi_data_misoZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47794),
            .ce(N__29780),
            .sr(N__52992));
    defparam RAM_nWE_obuf_RNO_LC_11_14_2.C_ON=1'b0;
    defparam RAM_nWE_obuf_RNO_LC_11_14_2.SEQ_MODE=4'b0000;
    defparam RAM_nWE_obuf_RNO_LC_11_14_2.LUT_INIT=16'b1010101011111111;
    LogicCell40 RAM_nWE_obuf_RNO_LC_11_14_2 (
            .in0(N__27617),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29939),
            .lcout(RAM_nWE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sADC_clk_prev_RNIM9TK_LC_11_14_3.C_ON=1'b0;
    defparam sADC_clk_prev_RNIM9TK_LC_11_14_3.SEQ_MODE=4'b0000;
    defparam sADC_clk_prev_RNIM9TK_LC_11_14_3.LUT_INIT=16'b1101110111111111;
    LogicCell40 sADC_clk_prev_RNIM9TK_LC_11_14_3 (
            .in0(N__32351),
            .in1(N__27635),
            .in2(_gnd_net_),
            .in3(N__27616),
            .lcout(sRAM_ADD_0_sqmuxa_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_rpi_ibuf_RNI4GQD1_LC_11_14_4.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNI4GQD1_LC_11_14_4.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNI4GQD1_LC_11_14_4.LUT_INIT=16'b0000000010101010;
    LogicCell40 reset_rpi_ibuf_RNI4GQD1_LC_11_14_4 (
            .in0(N__32350),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27575),
            .lcout(N_1470_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sRead_data_LC_11_15_0.C_ON=1'b0;
    defparam sRead_data_LC_11_15_0.SEQ_MODE=4'b1010;
    defparam sRead_data_LC_11_15_0.LUT_INIT=16'b1110111000000100;
    LogicCell40 sRead_data_LC_11_15_0 (
            .in0(N__29933),
            .in1(N__29851),
            .in2(N__27486),
            .in3(N__27470),
            .lcout(sRead_dataZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47805),
            .ce(),
            .sr(N__52987));
    defparam sCounterRAM_RNISREI1_7_LC_11_15_2.C_ON=1'b0;
    defparam sCounterRAM_RNISREI1_7_LC_11_15_2.SEQ_MODE=4'b0000;
    defparam sCounterRAM_RNISREI1_7_LC_11_15_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounterRAM_RNISREI1_7_LC_11_15_2 (
            .in0(N__27456),
            .in1(N__27438),
            .in2(N__27417),
            .in3(N__27396),
            .lcout(),
            .ltout(spi_data_miso_0_sqmuxa_2_i_o2_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterRAM_RNIS8L63_1_LC_11_15_3.C_ON=1'b0;
    defparam sCounterRAM_RNIS8L63_1_LC_11_15_3.SEQ_MODE=4'b0000;
    defparam sCounterRAM_RNIS8L63_1_LC_11_15_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 sCounterRAM_RNIS8L63_1_LC_11_15_3 (
            .in0(N__28038),
            .in1(N__28020),
            .in2(N__27999),
            .in3(N__27996),
            .lcout(N_75),
            .ltout(N_75_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_23_c_RNIGRPG4_LC_11_15_4.C_ON=1'b0;
    defparam un4_sacqtime_cry_23_c_RNIGRPG4_LC_11_15_4.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_23_c_RNIGRPG4_LC_11_15_4.LUT_INIT=16'b1110111110101111;
    LogicCell40 un4_sacqtime_cry_23_c_RNIGRPG4_LC_11_15_4 (
            .in0(N__27858),
            .in1(N__32217),
            .in2(N__27984),
            .in3(N__31916),
            .lcout(N_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sSPI_MSB0LSB1_RNINK761_LC_11_15_5.C_ON=1'b0;
    defparam sSPI_MSB0LSB1_RNINK761_LC_11_15_5.SEQ_MODE=4'b0000;
    defparam sSPI_MSB0LSB1_RNINK761_LC_11_15_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 sSPI_MSB0LSB1_RNINK761_LC_11_15_5 (
            .in0(_gnd_net_),
            .in1(N__27979),
            .in2(_gnd_net_),
            .in3(N__27897),
            .lcout(N_88),
            .ltout(N_88_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPointerReset_RNILL2C1_LC_11_15_6.C_ON=1'b0;
    defparam sEEPointerReset_RNILL2C1_LC_11_15_6.SEQ_MODE=4'b0000;
    defparam sEEPointerReset_RNILL2C1_LC_11_15_6.LUT_INIT=16'b1011101011111010;
    LogicCell40 sEEPointerReset_RNILL2C1_LC_11_15_6 (
            .in0(N__33434),
            .in1(N__31915),
            .in2(N__27852),
            .in3(N__32216),
            .lcout(N_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_9_RNO_0_15_LC_11_16_1.C_ON=1'b0;
    defparam RAM_DATA_cl_9_RNO_0_15_LC_11_16_1.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_9_RNO_0_15_LC_11_16_1.LUT_INIT=16'b0000000010101010;
    LogicCell40 RAM_DATA_cl_9_RNO_0_15_LC_11_16_1 (
            .in0(N__31684),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27806),
            .lcout(),
            .ltout(N_93_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_9_15_LC_11_16_2.C_ON=1'b0;
    defparam RAM_DATA_cl_9_15_LC_11_16_2.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_9_15_LC_11_16_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 RAM_DATA_cl_9_15_LC_11_16_2 (
            .in0(N__31885),
            .in1(N__32214),
            .in2(N__27825),
            .in3(N__32354),
            .lcout(RAM_DATA_cl_9Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47815),
            .ce(),
            .sr(N__52982));
    defparam RAM_DATA_cl_RNO_0_15_LC_11_16_3.C_ON=1'b0;
    defparam RAM_DATA_cl_RNO_0_15_LC_11_16_3.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_RNO_0_15_LC_11_16_3.LUT_INIT=16'b0000000010101010;
    LogicCell40 RAM_DATA_cl_RNO_0_15_LC_11_16_3 (
            .in0(N__31685),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27776),
            .lcout(),
            .ltout(N_98_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_15_LC_11_16_4.C_ON=1'b0;
    defparam RAM_DATA_cl_15_LC_11_16_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_15_LC_11_16_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 RAM_DATA_cl_15_LC_11_16_4 (
            .in0(N__31883),
            .in1(N__32212),
            .in2(N__27795),
            .in3(N__32352),
            .lcout(RAM_DATA_clZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47815),
            .ce(),
            .sr(N__52982));
    defparam RAM_DATA_cl_8_RNO_0_15_LC_11_16_5.C_ON=1'b0;
    defparam RAM_DATA_cl_8_RNO_0_15_LC_11_16_5.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_8_RNO_0_15_LC_11_16_5.LUT_INIT=16'b0000000010101010;
    LogicCell40 RAM_DATA_cl_8_RNO_0_15_LC_11_16_5 (
            .in0(N__31683),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28310),
            .lcout(),
            .ltout(N_96_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_8_15_LC_11_16_6.C_ON=1'b0;
    defparam RAM_DATA_cl_8_15_LC_11_16_6.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_8_15_LC_11_16_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 RAM_DATA_cl_8_15_LC_11_16_6 (
            .in0(N__31884),
            .in1(N__32213),
            .in2(N__28329),
            .in3(N__32353),
            .lcout(RAM_DATA_cl_8Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47815),
            .ce(),
            .sr(N__52982));
    defparam un4_sacqtime_cry_23_c_RNITTS3_LC_11_16_7.C_ON=1'b0;
    defparam un4_sacqtime_cry_23_c_RNITTS3_LC_11_16_7.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_23_c_RNITTS3_LC_11_16_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 un4_sacqtime_cry_23_c_RNITTS3_LC_11_16_7 (
            .in0(_gnd_net_),
            .in1(N__32211),
            .in2(_gnd_net_),
            .in3(N__31882),
            .lcout(un4_sacqtime_cry_23_c_RNITTSZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sRAM_ADD_14_LC_11_17_0.C_ON=1'b0;
    defparam sRAM_ADD_14_LC_11_17_0.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_14_LC_11_17_0.LUT_INIT=16'b1011100011110000;
    LogicCell40 sRAM_ADD_14_LC_11_17_0 (
            .in0(N__33015),
            .in1(N__32196),
            .in2(N__28299),
            .in3(N__31960),
            .lcout(RAM_ADD_c_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47823),
            .ce(N__30267),
            .sr(_gnd_net_));
    defparam sRAM_ADD_15_LC_11_17_1.C_ON=1'b0;
    defparam sRAM_ADD_15_LC_11_17_1.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_15_LC_11_17_1.LUT_INIT=16'b1101111110000000;
    LogicCell40 sRAM_ADD_15_LC_11_17_1 (
            .in0(N__31957),
            .in1(N__32994),
            .in2(N__32226),
            .in3(N__28248),
            .lcout(RAM_ADD_c_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47823),
            .ce(N__30267),
            .sr(_gnd_net_));
    defparam sRAM_ADD_16_LC_11_17_2.C_ON=1'b0;
    defparam sRAM_ADD_16_LC_11_17_2.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_16_LC_11_17_2.LUT_INIT=16'b1100101010101010;
    LogicCell40 sRAM_ADD_16_LC_11_17_2 (
            .in0(N__28209),
            .in1(N__32973),
            .in2(N__32221),
            .in3(N__31961),
            .lcout(RAM_ADD_c_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47823),
            .ce(N__30267),
            .sr(_gnd_net_));
    defparam sRAM_ADD_17_LC_11_17_3.C_ON=1'b0;
    defparam sRAM_ADD_17_LC_11_17_3.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_17_LC_11_17_3.LUT_INIT=16'b1110110001001100;
    LogicCell40 sRAM_ADD_17_LC_11_17_3 (
            .in0(N__31958),
            .in1(N__28164),
            .in2(N__32227),
            .in3(N__32952),
            .lcout(RAM_ADD_c_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47823),
            .ce(N__30267),
            .sr(_gnd_net_));
    defparam sRAM_ADD_18_LC_11_17_4.C_ON=1'b0;
    defparam sRAM_ADD_18_LC_11_17_4.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_18_LC_11_17_4.LUT_INIT=16'b1011100011110000;
    LogicCell40 sRAM_ADD_18_LC_11_17_4 (
            .in0(N__33327),
            .in1(N__32197),
            .in2(N__28125),
            .in3(N__31962),
            .lcout(RAM_ADD_c_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47823),
            .ce(N__30267),
            .sr(_gnd_net_));
    defparam sRAM_ADD_2_LC_11_17_5.C_ON=1'b0;
    defparam sRAM_ADD_2_LC_11_17_5.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_2_LC_11_17_5.LUT_INIT=16'b1110110001001100;
    LogicCell40 sRAM_ADD_2_LC_11_17_5 (
            .in0(N__31959),
            .in1(N__28080),
            .in2(N__32228),
            .in3(N__32925),
            .lcout(RAM_ADD_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47823),
            .ce(N__30267),
            .sr(_gnd_net_));
    defparam sRAM_ADD_3_LC_11_17_6.C_ON=1'b0;
    defparam sRAM_ADD_3_LC_11_17_6.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_3_LC_11_17_6.LUT_INIT=16'b1111100001110000;
    LogicCell40 sRAM_ADD_3_LC_11_17_6 (
            .in0(N__31956),
            .in1(N__32198),
            .in2(N__28689),
            .in3(N__32904),
            .lcout(RAM_ADD_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47823),
            .ce(N__30267),
            .sr(_gnd_net_));
    defparam sRAM_ADD_4_LC_11_17_7.C_ON=1'b0;
    defparam sRAM_ADD_4_LC_11_17_7.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_4_LC_11_17_7.LUT_INIT=16'b1011111110000000;
    LogicCell40 sRAM_ADD_4_LC_11_17_7 (
            .in0(N__32883),
            .in1(N__31955),
            .in2(N__32229),
            .in3(N__28650),
            .lcout(RAM_ADD_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47823),
            .ce(N__30267),
            .sr(_gnd_net_));
    defparam sRAM_ADD_5_LC_11_18_0.C_ON=1'b0;
    defparam sRAM_ADD_5_LC_11_18_0.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_5_LC_11_18_0.LUT_INIT=16'b1110001010101010;
    LogicCell40 sRAM_ADD_5_LC_11_18_0 (
            .in0(N__28605),
            .in1(N__32163),
            .in2(N__32859),
            .in3(N__31912),
            .lcout(RAM_ADD_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(N__30263),
            .sr(_gnd_net_));
    defparam sRAM_ADD_6_LC_11_18_1.C_ON=1'b0;
    defparam sRAM_ADD_6_LC_11_18_1.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_6_LC_11_18_1.LUT_INIT=16'b1110110001001100;
    LogicCell40 sRAM_ADD_6_LC_11_18_1 (
            .in0(N__31910),
            .in1(N__28560),
            .in2(N__32219),
            .in3(N__32838),
            .lcout(RAM_ADD_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(N__30263),
            .sr(_gnd_net_));
    defparam sRAM_ADD_7_LC_11_18_2.C_ON=1'b0;
    defparam sRAM_ADD_7_LC_11_18_2.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_7_LC_11_18_2.LUT_INIT=16'b1011100011110000;
    LogicCell40 sRAM_ADD_7_LC_11_18_2 (
            .in0(N__32820),
            .in1(N__32164),
            .in2(N__28512),
            .in3(N__31913),
            .lcout(RAM_ADD_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(N__30263),
            .sr(_gnd_net_));
    defparam sRAM_ADD_8_LC_11_18_3.C_ON=1'b0;
    defparam sRAM_ADD_8_LC_11_18_3.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_8_LC_11_18_3.LUT_INIT=16'b1110110001001100;
    LogicCell40 sRAM_ADD_8_LC_11_18_3 (
            .in0(N__31911),
            .in1(N__28464),
            .in2(N__32220),
            .in3(N__32802),
            .lcout(RAM_ADD_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(N__30263),
            .sr(_gnd_net_));
    defparam sRAM_ADD_9_LC_11_18_6.C_ON=1'b0;
    defparam sRAM_ADD_9_LC_11_18_6.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_9_LC_11_18_6.LUT_INIT=16'b1011100011110000;
    LogicCell40 sRAM_ADD_9_LC_11_18_6 (
            .in0(N__32781),
            .in1(N__32165),
            .in2(N__28419),
            .in3(N__31914),
            .lcout(RAM_ADD_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47833),
            .ce(N__30263),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_15_15_LC_11_19_6.C_ON=1'b0;
    defparam RAM_DATA_cl_15_15_LC_11_19_6.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_15_15_LC_11_19_6.LUT_INIT=16'b0000000010000000;
    LogicCell40 RAM_DATA_cl_15_15_LC_11_19_6 (
            .in0(N__31963),
            .in1(N__32444),
            .in2(N__32218),
            .in3(N__28371),
            .lcout(RAM_DATA_cl_15Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47840),
            .ce(),
            .sr(N__52972));
    defparam RAM_DATA_cl_13_15_LC_11_19_7.C_ON=1'b0;
    defparam RAM_DATA_cl_13_15_LC_11_19_7.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_13_15_LC_11_19_7.LUT_INIT=16'b0100000000000000;
    LogicCell40 RAM_DATA_cl_13_15_LC_11_19_7 (
            .in0(N__30492),
            .in1(N__32159),
            .in2(N__32504),
            .in3(N__31964),
            .lcout(RAM_DATA_cl_13Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47840),
            .ce(),
            .sr(N__52972));
    defparam RAM_DATA_cl_1_15_LC_11_20_0.C_ON=1'b0;
    defparam RAM_DATA_cl_1_15_LC_11_20_0.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_1_15_LC_11_20_0.LUT_INIT=16'b0100000000000000;
    LogicCell40 RAM_DATA_cl_1_15_LC_11_20_0 (
            .in0(N__30528),
            .in1(N__32151),
            .in2(N__32505),
            .in3(N__31965),
            .lcout(RAM_DATA_cl_1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47848),
            .ce(),
            .sr(N__52968));
    defparam RAM_DATA_cl_2_15_LC_11_20_6.C_ON=1'b0;
    defparam RAM_DATA_cl_2_15_LC_11_20_6.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_2_15_LC_11_20_6.LUT_INIT=16'b0100000000000000;
    LogicCell40 RAM_DATA_cl_2_15_LC_11_20_6 (
            .in0(N__30459),
            .in1(N__32152),
            .in2(N__32506),
            .in3(N__31966),
            .lcout(RAM_DATA_cl_2Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47848),
            .ce(),
            .sr(N__52968));
    defparam \spi_slave_inst.spi_cs_LC_12_1_0 .C_ON=1'b0;
    defparam \spi_slave_inst.spi_cs_LC_12_1_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.spi_cs_LC_12_1_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \spi_slave_inst.spi_cs_LC_12_1_0  (
            .in0(N__33285),
            .in1(N__38564),
            .in2(_gnd_net_),
            .in3(N__52425),
            .lcout(\spi_slave_inst.spi_csZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.spi_sclk_LC_12_1_6 .C_ON=1'b0;
    defparam \spi_slave_inst.spi_sclk_LC_12_1_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.spi_sclk_LC_12_1_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \spi_slave_inst.spi_sclk_LC_12_1_6  (
            .in0(N__28719),
            .in1(N__38565),
            .in2(_gnd_net_),
            .in3(N__52343),
            .lcout(spi_sclk),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_0_LC_12_2_4.C_ON=1'b0;
    defparam sDAC_data_0_LC_12_2_4.SEQ_MODE=4'b1010;
    defparam sDAC_data_0_LC_12_2_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_0_LC_12_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53241),
            .ce(N__42233),
            .sr(N__53090));
    defparam \spi_slave_inst.rxdata_reg_i_0_LC_12_3_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_0_LC_12_3_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_0_LC_12_3_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_0_LC_12_3_0  (
            .in0(N__30795),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_data_mosi_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(N__28767),
            .sr(N__53079));
    defparam \spi_slave_inst.rxdata_reg_i_1_LC_12_3_1 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_1_LC_12_3_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_1_LC_12_3_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_1_LC_12_3_1  (
            .in0(N__30783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_data_mosi_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(N__28767),
            .sr(N__53079));
    defparam \spi_slave_inst.rxdata_reg_i_2_LC_12_3_2 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_2_LC_12_3_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_2_LC_12_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_2_LC_12_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30771),
            .lcout(spi_data_mosi_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(N__28767),
            .sr(N__53079));
    defparam \spi_slave_inst.rxdata_reg_i_3_LC_12_3_3 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_3_LC_12_3_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_3_LC_12_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_3_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30759),
            .lcout(spi_data_mosi_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(N__28767),
            .sr(N__53079));
    defparam \spi_slave_inst.rxdata_reg_i_4_LC_12_3_4 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_4_LC_12_3_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_4_LC_12_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_4_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30747),
            .lcout(spi_data_mosi_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(N__28767),
            .sr(N__53079));
    defparam \spi_slave_inst.rxdata_reg_i_5_LC_12_3_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_5_LC_12_3_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_5_LC_12_3_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_5_LC_12_3_5  (
            .in0(N__30735),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(spi_data_mosi_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(N__28767),
            .sr(N__53079));
    defparam \spi_slave_inst.rxdata_reg_i_6_LC_12_3_6 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_6_LC_12_3_6 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_6_LC_12_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_6_LC_12_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30723),
            .lcout(spi_data_mosi_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(N__28767),
            .sr(N__53079));
    defparam \spi_slave_inst.rxdata_reg_i_7_LC_12_3_7 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_7_LC_12_3_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rxdata_reg_i_7_LC_12_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_7_LC_12_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30711),
            .lcout(spi_data_mosi_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47834),
            .ce(N__28767),
            .sr(N__53079));
    defparam \spi_slave_inst.rx_done_reg1_i_RNID541_LC_12_4_2 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_done_reg1_i_RNID541_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rx_done_reg1_i_RNID541_LC_12_4_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \spi_slave_inst.rx_done_reg1_i_RNID541_LC_12_4_2  (
            .in0(_gnd_net_),
            .in1(N__28805),
            .in2(_gnd_net_),
            .in3(N__28794),
            .lcout(\spi_slave_inst.rx_done_reg1_i_RNIDZ0Z541 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rxdata_reg_i_RNINNBS_2_LC_12_4_3 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_RNINNBS_2_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rxdata_reg_i_RNINNBS_2_LC_12_4_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_RNINNBS_2_LC_12_4_3  (
            .in0(N__48910),
            .in1(N__49415),
            .in2(N__47948),
            .in3(N__49906),
            .lcout(\spi_slave_inst.un1_spointer11_2_0_a2_0_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_master_inst.spi_data_path_u1.data_in_10_LC_12_5_0 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_10_LC_12_5_0 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_10_LC_12_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_10_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39468),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53244),
            .ce(N__28841),
            .sr(N__53057));
    defparam \spi_master_inst.spi_data_path_u1.data_in_13_LC_12_5_1 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_13_LC_12_5_1 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_13_LC_12_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_13_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37731),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53244),
            .ce(N__28841),
            .sr(N__53057));
    defparam \spi_master_inst.spi_data_path_u1.data_in_4_LC_12_5_2 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_4_LC_12_5_2 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_4_LC_12_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_4_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41202),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53244),
            .ce(N__28841),
            .sr(N__53057));
    defparam \spi_master_inst.spi_data_path_u1.data_in_5_LC_12_5_3 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_5_LC_12_5_3 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_5_LC_12_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_5_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33768),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53244),
            .ce(N__28841),
            .sr(N__53057));
    defparam \spi_master_inst.spi_data_path_u1.data_in_0_LC_12_5_4 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_0_LC_12_5_4 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_0_LC_12_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_0_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28899),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53244),
            .ce(N__28841),
            .sr(N__53057));
    defparam \spi_master_inst.spi_data_path_u1.data_in_7_LC_12_5_5 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_7_LC_12_5_5 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_7_LC_12_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_7_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37425),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53244),
            .ce(N__28841),
            .sr(N__53057));
    defparam \spi_master_inst.spi_data_path_u1.data_in_8_LC_12_5_6 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_8_LC_12_5_6 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_8_LC_12_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_8_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40917),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53244),
            .ce(N__28841),
            .sr(N__53057));
    defparam \spi_master_inst.spi_data_path_u1.data_in_9_LC_12_5_7 .C_ON=1'b0;
    defparam \spi_master_inst.spi_data_path_u1.data_in_9_LC_12_5_7 .SEQ_MODE=4'b1010;
    defparam \spi_master_inst.spi_data_path_u1.data_in_9_LC_12_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_master_inst.spi_data_path_u1.data_in_9_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39171),
            .lcout(\spi_master_inst.spi_data_path_u1.data_inZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53244),
            .ce(N__28841),
            .sr(N__53057));
    defparam sDAC_mem_4_1_LC_12_6_0.C_ON=1'b0;
    defparam sDAC_mem_4_1_LC_12_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_1_LC_12_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_1_LC_12_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50454),
            .lcout(sDAC_mem_4Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47806),
            .ce(N__39635),
            .sr(N__53047));
    defparam sDAC_mem_4_4_LC_12_6_1.C_ON=1'b0;
    defparam sDAC_mem_4_4_LC_12_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_4_LC_12_6_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_4_4_LC_12_6_1 (
            .in0(N__48988),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_4Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47806),
            .ce(N__39635),
            .sr(N__53047));
    defparam sDAC_mem_23_0_LC_12_7_0.C_ON=1'b0;
    defparam sDAC_mem_23_0_LC_12_7_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_0_LC_12_7_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_23_0_LC_12_7_0 (
            .in0(N__50881),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_23Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47795),
            .ce(N__28988),
            .sr(N__53038));
    defparam sDAC_mem_23_1_LC_12_7_1.C_ON=1'b0;
    defparam sDAC_mem_23_1_LC_12_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_1_LC_12_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_1_LC_12_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50455),
            .lcout(sDAC_mem_23Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47795),
            .ce(N__28988),
            .sr(N__53038));
    defparam sDAC_mem_23_2_LC_12_7_2.C_ON=1'b0;
    defparam sDAC_mem_23_2_LC_12_7_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_2_LC_12_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_2_LC_12_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50023),
            .lcout(sDAC_mem_23Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47795),
            .ce(N__28988),
            .sr(N__53038));
    defparam sDAC_mem_23_3_LC_12_7_3.C_ON=1'b0;
    defparam sDAC_mem_23_3_LC_12_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_3_LC_12_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_3_LC_12_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49572),
            .lcout(sDAC_mem_23Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47795),
            .ce(N__28988),
            .sr(N__53038));
    defparam sDAC_mem_23_4_LC_12_7_4.C_ON=1'b0;
    defparam sDAC_mem_23_4_LC_12_7_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_4_LC_12_7_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_23_4_LC_12_7_4 (
            .in0(N__49076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_23Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47795),
            .ce(N__28988),
            .sr(N__53038));
    defparam sDAC_mem_23_5_LC_12_7_5.C_ON=1'b0;
    defparam sDAC_mem_23_5_LC_12_7_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_5_LC_12_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_5_LC_12_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46861),
            .lcout(sDAC_mem_23Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47795),
            .ce(N__28988),
            .sr(N__53038));
    defparam sDAC_mem_23_6_LC_12_7_6.C_ON=1'b0;
    defparam sDAC_mem_23_6_LC_12_7_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_23_6_LC_12_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_23_6_LC_12_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48160),
            .lcout(sDAC_mem_23Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47795),
            .ce(N__28988),
            .sr(N__53038));
    defparam sDAC_mem_33_0_LC_12_8_0.C_ON=1'b0;
    defparam sDAC_mem_33_0_LC_12_8_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_0_LC_12_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_0_LC_12_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51025),
            .lcout(sDAC_mem_33Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47780),
            .ce(N__30858),
            .sr(N__53027));
    defparam sDAC_mem_33_1_LC_12_8_1.C_ON=1'b0;
    defparam sDAC_mem_33_1_LC_12_8_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_1_LC_12_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_1_LC_12_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50456),
            .lcout(sDAC_mem_33Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47780),
            .ce(N__30858),
            .sr(N__53027));
    defparam sDAC_mem_33_2_LC_12_8_2.C_ON=1'b0;
    defparam sDAC_mem_33_2_LC_12_8_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_2_LC_12_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_2_LC_12_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50024),
            .lcout(sDAC_mem_33Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47780),
            .ce(N__30858),
            .sr(N__53027));
    defparam sDAC_mem_33_3_LC_12_8_3.C_ON=1'b0;
    defparam sDAC_mem_33_3_LC_12_8_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_3_LC_12_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_3_LC_12_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49573),
            .lcout(sDAC_mem_33Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47780),
            .ce(N__30858),
            .sr(N__53027));
    defparam sDAC_mem_33_4_LC_12_8_4.C_ON=1'b0;
    defparam sDAC_mem_33_4_LC_12_8_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_4_LC_12_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_4_LC_12_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49131),
            .lcout(sDAC_mem_33Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47780),
            .ce(N__30858),
            .sr(N__53027));
    defparam sDAC_mem_33_5_LC_12_8_5.C_ON=1'b0;
    defparam sDAC_mem_33_5_LC_12_8_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_5_LC_12_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_5_LC_12_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46958),
            .lcout(sDAC_mem_33Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47780),
            .ce(N__30858),
            .sr(N__53027));
    defparam sDAC_mem_33_6_LC_12_8_6.C_ON=1'b0;
    defparam sDAC_mem_33_6_LC_12_8_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_6_LC_12_8_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_33_6_LC_12_8_6 (
            .in0(N__48161),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_33Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47780),
            .ce(N__30858),
            .sr(N__53027));
    defparam sDAC_mem_33_7_LC_12_8_7.C_ON=1'b0;
    defparam sDAC_mem_33_7_LC_12_8_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_33_7_LC_12_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_33_7_LC_12_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48597),
            .lcout(sDAC_mem_33Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47780),
            .ce(N__30858),
            .sr(N__53027));
    defparam sDAC_mem_1_0_LC_12_9_0.C_ON=1'b0;
    defparam sDAC_mem_1_0_LC_12_9_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_0_LC_12_9_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_1_0_LC_12_9_0 (
            .in0(N__51026),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47766),
            .ce(N__42031),
            .sr(N__53019));
    defparam sDAC_mem_1_1_LC_12_9_1.C_ON=1'b0;
    defparam sDAC_mem_1_1_LC_12_9_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_1_LC_12_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_1_LC_12_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50457),
            .lcout(sDAC_mem_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47766),
            .ce(N__42031),
            .sr(N__53019));
    defparam sDAC_mem_1_2_LC_12_9_2.C_ON=1'b0;
    defparam sDAC_mem_1_2_LC_12_9_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_2_LC_12_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_2_LC_12_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50025),
            .lcout(sDAC_mem_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47766),
            .ce(N__42031),
            .sr(N__53019));
    defparam sDAC_mem_1_7_LC_12_9_3.C_ON=1'b0;
    defparam sDAC_mem_1_7_LC_12_9_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_7_LC_12_9_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_1_7_LC_12_9_3 (
            .in0(N__48598),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47766),
            .ce(N__42031),
            .sr(N__53019));
    defparam sAddress_RNI25GS1_1_LC_12_10_0.C_ON=1'b0;
    defparam sAddress_RNI25GS1_1_LC_12_10_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI25GS1_1_LC_12_10_0.LUT_INIT=16'b0001001000000000;
    LogicCell40 sAddress_RNI25GS1_1_LC_12_10_0 (
            .in0(N__44871),
            .in1(N__31071),
            .in2(N__40355),
            .in3(N__44723),
            .lcout(un1_spointer11_5_0_2),
            .ltout(un1_spointer11_5_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_0_2_LC_12_10_1.C_ON=1'b0;
    defparam sAddress_RNIA6242_0_2_LC_12_10_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_0_2_LC_12_10_1.LUT_INIT=16'b0000000001000000;
    LogicCell40 sAddress_RNIA6242_0_2_LC_12_10_1 (
            .in0(N__40518),
            .in1(N__44953),
            .in2(N__28914),
            .in3(N__40325),
            .lcout(sAddress_RNIA6242_0Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_1_2_LC_12_10_2.C_ON=1'b0;
    defparam sAddress_RNIA6242_1_2_LC_12_10_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_1_2_LC_12_10_2.LUT_INIT=16'b0000001000000000;
    LogicCell40 sAddress_RNIA6242_1_2_LC_12_10_2 (
            .in0(N__40323),
            .in1(N__40516),
            .in2(N__44961),
            .in3(N__30991),
            .lcout(sAddress_RNIA6242_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_6_1_LC_12_10_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_6_1_LC_12_10_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_6_1_LC_12_10_3.LUT_INIT=16'b0000000010001000;
    LogicCell40 sAddress_RNI9IH12_6_1_LC_12_10_3 (
            .in0(N__43142),
            .in1(N__44553),
            .in2(_gnd_net_),
            .in3(N__44444),
            .lcout(sDAC_mem_32_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_16_3_LC_12_10_4.C_ON=1'b0;
    defparam sAddress_RNI9IH12_16_3_LC_12_10_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_16_3_LC_12_10_4.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNI9IH12_16_3_LC_12_10_4 (
            .in0(N__40324),
            .in1(N__40517),
            .in2(N__44571),
            .in3(N__43141),
            .lcout(sDAC_mem_23_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sPointer_RNI5LBD1_0_LC_12_10_5.C_ON=1'b0;
    defparam sPointer_RNI5LBD1_0_LC_12_10_5.SEQ_MODE=4'b0000;
    defparam sPointer_RNI5LBD1_0_LC_12_10_5.LUT_INIT=16'b0100010000000000;
    LogicCell40 sPointer_RNI5LBD1_0_LC_12_10_5 (
            .in0(N__29176),
            .in1(N__43856),
            .in2(_gnd_net_),
            .in3(N__29127),
            .lcout(N_275),
            .ltout(N_275_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_rpi_ibuf_RNIHQCR1_LC_12_10_6.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNIHQCR1_LC_12_10_6.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNIHQCR1_LC_12_10_6.LUT_INIT=16'b0000000011000000;
    LogicCell40 reset_rpi_ibuf_RNIHQCR1_LC_12_10_6 (
            .in0(_gnd_net_),
            .in1(N__32558),
            .in2(N__28971),
            .in3(N__31070),
            .lcout(N_360),
            .ltout(N_360_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEPointerReset_RNO_0_LC_12_10_7.C_ON=1'b0;
    defparam sEEPointerReset_RNO_0_LC_12_10_7.SEQ_MODE=4'b0000;
    defparam sEEPointerReset_RNO_0_LC_12_10_7.LUT_INIT=16'b1111111100100000;
    LogicCell40 sEEPointerReset_RNO_0_LC_12_10_7 (
            .in0(N__44549),
            .in1(N__44443),
            .in2(N__28968),
            .in3(N__28965),
            .lcout(N_132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_0_0_LC_12_11_0.C_ON=1'b0;
    defparam sAddress_RNIA6242_0_0_LC_12_11_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_0_0_LC_12_11_0.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNIA6242_0_0_LC_12_11_0 (
            .in0(N__40329),
            .in1(N__31073),
            .in2(N__28935),
            .in3(N__44716),
            .lcout(sAddress_RNIA6242_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIAM2A_1_LC_12_11_1.C_ON=1'b0;
    defparam sAddress_RNIAM2A_1_LC_12_11_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNIAM2A_1_LC_12_11_1.LUT_INIT=16'b0000100001010000;
    LogicCell40 sAddress_RNIAM2A_1_LC_12_11_1 (
            .in0(N__44959),
            .in1(N__40328),
            .in2(N__40539),
            .in3(N__44870),
            .lcout(un1_spointer11_7_0_tz),
            .ltout(un1_spointer11_7_0_tz_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNID9242_3_LC_12_11_2.C_ON=1'b0;
    defparam sAddress_RNID9242_3_LC_12_11_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNID9242_3_LC_12_11_2.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNID9242_3_LC_12_11_2 (
            .in0(N__40519),
            .in1(N__31074),
            .in2(N__28926),
            .in3(N__44717),
            .lcout(sAddress_RNID9242Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_0_LC_12_11_3.C_ON=1'b0;
    defparam sAddress_0_LC_12_11_3.SEQ_MODE=4'b1010;
    defparam sAddress_0_LC_12_11_3.LUT_INIT=16'b0000000010101010;
    LogicCell40 sAddress_0_LC_12_11_3 (
            .in0(N__50873),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43860),
            .lcout(sAddressZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47741),
            .ce(N__43771),
            .sr(N__53006));
    defparam sAddress_3_LC_12_11_4.C_ON=1'b0;
    defparam sAddress_3_LC_12_11_4.SEQ_MODE=4'b1010;
    defparam sAddress_3_LC_12_11_4.LUT_INIT=16'b0101010100000000;
    LogicCell40 sAddress_3_LC_12_11_4 (
            .in0(N__43861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49571),
            .lcout(sAddressZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47741),
            .ce(N__43771),
            .sr(N__53006));
    defparam sAddress_5_LC_12_11_5.C_ON=1'b0;
    defparam sAddress_5_LC_12_11_5.SEQ_MODE=4'b1010;
    defparam sAddress_5_LC_12_11_5.LUT_INIT=16'b0000000011001100;
    LogicCell40 sAddress_5_LC_12_11_5 (
            .in0(_gnd_net_),
            .in1(N__46957),
            .in2(_gnd_net_),
            .in3(N__43862),
            .lcout(sAddressZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47741),
            .ce(N__43771),
            .sr(N__53006));
    defparam \spi_slave_inst.rxdata_reg_i_RNILLBS_1_LC_12_11_6 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_RNILLBS_1_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rxdata_reg_i_RNILLBS_1_LC_12_11_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_RNILLBS_1_LC_12_11_6  (
            .in0(N__46956),
            .in1(N__50560),
            .in2(N__48672),
            .in3(N__50872),
            .lcout(),
            .ltout(\spi_slave_inst.un1_spointer11_2_0_a2_0_6_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.rxdata_reg_i_RNIH2363_1_LC_12_11_7 .C_ON=1'b0;
    defparam \spi_slave_inst.rxdata_reg_i_RNIH2363_1_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.rxdata_reg_i_RNIH2363_1_LC_12_11_7 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \spi_slave_inst.rxdata_reg_i_RNIH2363_1_LC_12_11_7  (
            .in0(N__29229),
            .in1(N__29144),
            .in2(N__29220),
            .in3(N__29129),
            .lcout(un1_spointer11_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_5_3_LC_12_12_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_5_3_LC_12_12_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_5_3_LC_12_12_0.LUT_INIT=16'b0100000000000000;
    LogicCell40 sAddress_RNI9IH12_5_3_LC_12_12_0 (
            .in0(N__40532),
            .in1(N__40334),
            .in2(N__46207),
            .in3(N__43145),
            .lcout(sDAC_mem_22_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI5B15_1_1_LC_12_12_1.C_ON=1'b0;
    defparam sAddress_RNI5B15_1_1_LC_12_12_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI5B15_1_1_LC_12_12_1.LUT_INIT=16'b0000000011001100;
    LogicCell40 sAddress_RNI5B15_1_1_LC_12_12_1 (
            .in0(_gnd_net_),
            .in1(N__44958),
            .in2(_gnd_net_),
            .in3(N__44868),
            .lcout(N_285),
            .ltout(N_285_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_18_3_LC_12_12_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_18_3_LC_12_12_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_18_3_LC_12_12_2.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNI9IH12_18_3_LC_12_12_2 (
            .in0(N__40531),
            .in1(N__40333),
            .in2(N__29199),
            .in3(N__43143),
            .lcout(sDAC_mem_21_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_5_1_LC_12_12_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_5_1_LC_12_12_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_5_1_LC_12_12_3.LUT_INIT=16'b0000000010001000;
    LogicCell40 sAddress_RNI9IH12_5_1_LC_12_12_3 (
            .in0(N__43144),
            .in1(N__46184),
            .in2(_gnd_net_),
            .in3(N__46068),
            .lcout(sDAC_mem_29_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigInternal_RNO_1_LC_12_12_5.C_ON=1'b0;
    defparam sEETrigInternal_RNO_1_LC_12_12_5.SEQ_MODE=4'b0000;
    defparam sEETrigInternal_RNO_1_LC_12_12_5.LUT_INIT=16'b1111111111111011;
    LogicCell40 sEETrigInternal_RNO_1_LC_12_12_5 (
            .in0(N__46067),
            .in1(N__43260),
            .in2(N__29196),
            .in3(N__31090),
            .lcout(),
            .ltout(N_116_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigInternal_RNO_0_LC_12_12_6.C_ON=1'b0;
    defparam sEETrigInternal_RNO_0_LC_12_12_6.SEQ_MODE=4'b0000;
    defparam sEETrigInternal_RNO_0_LC_12_12_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 sEETrigInternal_RNO_0_LC_12_12_6 (
            .in0(_gnd_net_),
            .in1(N__51078),
            .in2(N__29148),
            .in3(N__29040),
            .lcout(),
            .ltout(N_117_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEETrigInternal_LC_12_12_7.C_ON=1'b0;
    defparam sEETrigInternal_LC_12_12_7.SEQ_MODE=4'b1010;
    defparam sEETrigInternal_LC_12_12_7.LUT_INIT=16'b1100000010101010;
    LogicCell40 sEETrigInternal_LC_12_12_7 (
            .in0(N__29041),
            .in1(N__29145),
            .in2(N__29133),
            .in3(N__29130),
            .lcout(sEETrigInternalZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47755),
            .ce(),
            .sr(N__52998));
    defparam sEEPoff_0_LC_12_13_0.C_ON=1'b0;
    defparam sEEPoff_0_LC_12_13_0.SEQ_MODE=4'b1010;
    defparam sEEPoff_0_LC_12_13_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPoff_0_LC_12_13_0 (
            .in0(N__51133),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPoffZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47767),
            .ce(N__30975),
            .sr(N__52991));
    defparam sEEPoff_1_LC_12_13_1.C_ON=1'b0;
    defparam sEEPoff_1_LC_12_13_1.SEQ_MODE=4'b1010;
    defparam sEEPoff_1_LC_12_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_1_LC_12_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50572),
            .lcout(sEEPoffZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47767),
            .ce(N__30975),
            .sr(N__52991));
    defparam sEEPoff_2_LC_12_13_2.C_ON=1'b0;
    defparam sEEPoff_2_LC_12_13_2.SEQ_MODE=4'b1010;
    defparam sEEPoff_2_LC_12_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_2_LC_12_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50026),
            .lcout(sEEPoffZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47767),
            .ce(N__30975),
            .sr(N__52991));
    defparam sEEPoff_3_LC_12_13_3.C_ON=1'b0;
    defparam sEEPoff_3_LC_12_13_3.SEQ_MODE=4'b1011;
    defparam sEEPoff_3_LC_12_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_3_LC_12_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49574),
            .lcout(sEEPoffZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47767),
            .ce(N__30975),
            .sr(N__52991));
    defparam sEEPoff_4_LC_12_13_4.C_ON=1'b0;
    defparam sEEPoff_4_LC_12_13_4.SEQ_MODE=4'b1010;
    defparam sEEPoff_4_LC_12_13_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_4_LC_12_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49130),
            .lcout(sEEPoffZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47767),
            .ce(N__30975),
            .sr(N__52991));
    defparam sEEPoff_5_LC_12_13_5.C_ON=1'b0;
    defparam sEEPoff_5_LC_12_13_5.SEQ_MODE=4'b1010;
    defparam sEEPoff_5_LC_12_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_5_LC_12_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47045),
            .lcout(sEEPoffZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47767),
            .ce(N__30975),
            .sr(N__52991));
    defparam sEEPoff_6_LC_12_13_6.C_ON=1'b0;
    defparam sEEPoff_6_LC_12_13_6.SEQ_MODE=4'b1011;
    defparam sEEPoff_6_LC_12_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_6_LC_12_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48272),
            .lcout(sEEPoffZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47767),
            .ce(N__30975),
            .sr(N__52991));
    defparam sEEPoff_7_LC_12_13_7.C_ON=1'b0;
    defparam sEEPoff_7_LC_12_13_7.SEQ_MODE=4'b1011;
    defparam sEEPoff_7_LC_12_13_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPoff_7_LC_12_13_7 (
            .in0(N__48575),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPoffZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47767),
            .ce(N__30975),
            .sr(N__52991));
    defparam sEEPoff_10_LC_12_14_0.C_ON=1'b0;
    defparam sEEPoff_10_LC_12_14_0.SEQ_MODE=4'b1010;
    defparam sEEPoff_10_LC_12_14_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPoff_10_LC_12_14_0 (
            .in0(N__50180),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPoffZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47781),
            .ce(N__29337),
            .sr(N__52986));
    defparam sEEPoff_11_LC_12_14_1.C_ON=1'b0;
    defparam sEEPoff_11_LC_12_14_1.SEQ_MODE=4'b1010;
    defparam sEEPoff_11_LC_12_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_11_LC_12_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49575),
            .lcout(sEEPoffZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47781),
            .ce(N__29337),
            .sr(N__52986));
    defparam sEEPoff_12_LC_12_14_2.C_ON=1'b0;
    defparam sEEPoff_12_LC_12_14_2.SEQ_MODE=4'b1010;
    defparam sEEPoff_12_LC_12_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_12_LC_12_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49129),
            .lcout(sEEPoffZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47781),
            .ce(N__29337),
            .sr(N__52986));
    defparam sEEPoff_13_LC_12_14_3.C_ON=1'b0;
    defparam sEEPoff_13_LC_12_14_3.SEQ_MODE=4'b1010;
    defparam sEEPoff_13_LC_12_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_13_LC_12_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47053),
            .lcout(sEEPoffZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47781),
            .ce(N__29337),
            .sr(N__52986));
    defparam sEEPoff_14_LC_12_14_4.C_ON=1'b0;
    defparam sEEPoff_14_LC_12_14_4.SEQ_MODE=4'b1010;
    defparam sEEPoff_14_LC_12_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_14_LC_12_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48273),
            .lcout(sEEPoffZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47781),
            .ce(N__29337),
            .sr(N__52986));
    defparam sEEPoff_15_LC_12_14_5.C_ON=1'b0;
    defparam sEEPoff_15_LC_12_14_5.SEQ_MODE=4'b1010;
    defparam sEEPoff_15_LC_12_14_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEPoff_15_LC_12_14_5 (
            .in0(N__48576),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEPoffZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47781),
            .ce(N__29337),
            .sr(N__52986));
    defparam sEEPoff_8_LC_12_14_6.C_ON=1'b0;
    defparam sEEPoff_8_LC_12_14_6.SEQ_MODE=4'b1010;
    defparam sEEPoff_8_LC_12_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_8_LC_12_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51079),
            .lcout(sEEPoffZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47781),
            .ce(N__29337),
            .sr(N__52986));
    defparam sEEPoff_9_LC_12_14_7.C_ON=1'b0;
    defparam sEEPoff_9_LC_12_14_7.SEQ_MODE=4'b1010;
    defparam sEEPoff_9_LC_12_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEPoff_9_LC_12_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50573),
            .lcout(sEEPoffZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47781),
            .ce(N__29337),
            .sr(N__52986));
    defparam sCounterADC_0_LC_12_15_0.C_ON=1'b1;
    defparam sCounterADC_0_LC_12_15_0.SEQ_MODE=4'b1010;
    defparam sCounterADC_0_LC_12_15_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_0_LC_12_15_0 (
            .in0(N__38225),
            .in1(N__38267),
            .in2(_gnd_net_),
            .in3(N__29322),
            .lcout(sCounterADCZ0Z_0),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(sCounterADC_cry_0),
            .clk(N__47796),
            .ce(N__29940),
            .sr(N__52981));
    defparam sCounterADC_1_LC_12_15_1.C_ON=1'b1;
    defparam sCounterADC_1_LC_12_15_1.SEQ_MODE=4'b1010;
    defparam sCounterADC_1_LC_12_15_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_1_LC_12_15_1 (
            .in0(N__38203),
            .in1(N__38282),
            .in2(_gnd_net_),
            .in3(N__29319),
            .lcout(sCounterADCZ0Z_1),
            .ltout(),
            .carryin(sCounterADC_cry_0),
            .carryout(sCounterADC_cry_1),
            .clk(N__47796),
            .ce(N__29940),
            .sr(N__52981));
    defparam sCounterADC_2_LC_12_15_2.C_ON=1'b1;
    defparam sCounterADC_2_LC_12_15_2.SEQ_MODE=4'b1010;
    defparam sCounterADC_2_LC_12_15_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_2_LC_12_15_2 (
            .in0(N__38226),
            .in1(N__34350),
            .in2(_gnd_net_),
            .in3(N__29589),
            .lcout(sCounterADCZ0Z_2),
            .ltout(),
            .carryin(sCounterADC_cry_1),
            .carryout(sCounterADC_cry_2),
            .clk(N__47796),
            .ce(N__29940),
            .sr(N__52981));
    defparam sCounterADC_3_LC_12_15_3.C_ON=1'b1;
    defparam sCounterADC_3_LC_12_15_3.SEQ_MODE=4'b1010;
    defparam sCounterADC_3_LC_12_15_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_3_LC_12_15_3 (
            .in0(N__38204),
            .in1(N__34364),
            .in2(_gnd_net_),
            .in3(N__29586),
            .lcout(sCounterADCZ0Z_3),
            .ltout(),
            .carryin(sCounterADC_cry_2),
            .carryout(sCounterADC_cry_3),
            .clk(N__47796),
            .ce(N__29940),
            .sr(N__52981));
    defparam sCounterADC_4_LC_12_15_4.C_ON=1'b1;
    defparam sCounterADC_4_LC_12_15_4.SEQ_MODE=4'b1010;
    defparam sCounterADC_4_LC_12_15_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_4_LC_12_15_4 (
            .in0(N__38227),
            .in1(N__34304),
            .in2(_gnd_net_),
            .in3(N__29583),
            .lcout(sCounterADCZ0Z_4),
            .ltout(),
            .carryin(sCounterADC_cry_3),
            .carryout(sCounterADC_cry_4),
            .clk(N__47796),
            .ce(N__29940),
            .sr(N__52981));
    defparam sCounterADC_5_LC_12_15_5.C_ON=1'b1;
    defparam sCounterADC_5_LC_12_15_5.SEQ_MODE=4'b1010;
    defparam sCounterADC_5_LC_12_15_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_5_LC_12_15_5 (
            .in0(N__38205),
            .in1(N__34320),
            .in2(_gnd_net_),
            .in3(N__29580),
            .lcout(sCounterADCZ0Z_5),
            .ltout(),
            .carryin(sCounterADC_cry_4),
            .carryout(sCounterADC_cry_5),
            .clk(N__47796),
            .ce(N__29940),
            .sr(N__52981));
    defparam sCounterADC_6_LC_12_15_6.C_ON=1'b1;
    defparam sCounterADC_6_LC_12_15_6.SEQ_MODE=4'b1010;
    defparam sCounterADC_6_LC_12_15_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_6_LC_12_15_6 (
            .in0(N__38228),
            .in1(N__34274),
            .in2(_gnd_net_),
            .in3(N__29577),
            .lcout(sCounterADCZ0Z_6),
            .ltout(),
            .carryin(sCounterADC_cry_5),
            .carryout(sCounterADC_cry_6),
            .clk(N__47796),
            .ce(N__29940),
            .sr(N__52981));
    defparam sCounterADC_7_LC_12_15_7.C_ON=1'b0;
    defparam sCounterADC_7_LC_12_15_7.SEQ_MODE=4'b1010;
    defparam sCounterADC_7_LC_12_15_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sCounterADC_7_LC_12_15_7 (
            .in0(N__38206),
            .in1(N__34259),
            .in2(_gnd_net_),
            .in3(N__29574),
            .lcout(sCounterADCZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47796),
            .ce(N__29940),
            .sr(N__52981));
    defparam spi_data_miso_0_LC_12_16_2.C_ON=1'b0;
    defparam spi_data_miso_0_LC_12_16_2.SEQ_MODE=4'b1010;
    defparam spi_data_miso_0_LC_12_16_2.LUT_INIT=16'b1111111111100010;
    LogicCell40 spi_data_miso_0_LC_12_16_2 (
            .in0(N__29571),
            .in1(N__29856),
            .in2(N__29547),
            .in3(N__29920),
            .lcout(spi_data_misoZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47807),
            .ce(N__29787),
            .sr(N__52978));
    defparam spi_data_miso_1_LC_12_16_3.C_ON=1'b0;
    defparam spi_data_miso_1_LC_12_16_3.SEQ_MODE=4'b1011;
    defparam spi_data_miso_1_LC_12_16_3.LUT_INIT=16'b0101010000000100;
    LogicCell40 spi_data_miso_1_LC_12_16_3 (
            .in0(N__29921),
            .in1(N__29514),
            .in2(N__29869),
            .in3(N__29499),
            .lcout(spi_data_misoZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47807),
            .ce(N__29787),
            .sr(N__52978));
    defparam spi_data_miso_2_LC_12_16_4.C_ON=1'b0;
    defparam spi_data_miso_2_LC_12_16_4.SEQ_MODE=4'b1011;
    defparam spi_data_miso_2_LC_12_16_4.LUT_INIT=16'b0000000011100010;
    LogicCell40 spi_data_miso_2_LC_12_16_4 (
            .in0(N__29469),
            .in1(N__29860),
            .in2(N__29445),
            .in3(N__29922),
            .lcout(spi_data_misoZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47807),
            .ce(N__29787),
            .sr(N__52978));
    defparam spi_data_miso_3_LC_12_16_5.C_ON=1'b0;
    defparam spi_data_miso_3_LC_12_16_5.SEQ_MODE=4'b1010;
    defparam spi_data_miso_3_LC_12_16_5.LUT_INIT=16'b0101010000000100;
    LogicCell40 spi_data_miso_3_LC_12_16_5 (
            .in0(N__29923),
            .in1(N__30051),
            .in2(N__29870),
            .in3(N__30030),
            .lcout(spi_data_misoZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47807),
            .ce(N__29787),
            .sr(N__52978));
    defparam spi_data_miso_4_LC_12_16_6.C_ON=1'b0;
    defparam spi_data_miso_4_LC_12_16_6.SEQ_MODE=4'b1011;
    defparam spi_data_miso_4_LC_12_16_6.LUT_INIT=16'b0000000011100010;
    LogicCell40 spi_data_miso_4_LC_12_16_6 (
            .in0(N__29997),
            .in1(N__29864),
            .in2(N__29976),
            .in3(N__29924),
            .lcout(spi_data_misoZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47807),
            .ce(N__29787),
            .sr(N__52978));
    defparam spi_data_miso_5_LC_12_16_7.C_ON=1'b0;
    defparam spi_data_miso_5_LC_12_16_7.SEQ_MODE=4'b1011;
    defparam spi_data_miso_5_LC_12_16_7.LUT_INIT=16'b0100010101000000;
    LogicCell40 spi_data_miso_5_LC_12_16_7 (
            .in0(N__29925),
            .in1(N__29889),
            .in2(N__29871),
            .in3(N__29823),
            .lcout(spi_data_misoZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47807),
            .ce(N__29787),
            .sr(N__52978));
    defparam sRAM_ADD_0_LC_12_17_0.C_ON=1'b0;
    defparam sRAM_ADD_0_LC_12_17_0.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_0_LC_12_17_0.LUT_INIT=16'b1110010011001100;
    LogicCell40 sRAM_ADD_0_LC_12_17_0 (
            .in0(N__31936),
            .in1(N__29763),
            .in2(N__31623),
            .in3(N__32184),
            .lcout(RAM_ADD_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47816),
            .ce(N__30262),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_23_c_RNIQQ6O1_LC_12_17_1.C_ON=1'b0;
    defparam un4_sacqtime_cry_23_c_RNIQQ6O1_LC_12_17_1.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_23_c_RNIQQ6O1_LC_12_17_1.LUT_INIT=16'b0001101100110011;
    LogicCell40 un4_sacqtime_cry_23_c_RNIQQ6O1_LC_12_17_1 (
            .in0(N__32179),
            .in1(N__29718),
            .in2(N__29703),
            .in3(N__31934),
            .lcout(N_67_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un4_sacqtime_cry_23_c_RNIJ7QO_LC_12_17_2.C_ON=1'b0;
    defparam un4_sacqtime_cry_23_c_RNIJ7QO_LC_12_17_2.SEQ_MODE=4'b0000;
    defparam un4_sacqtime_cry_23_c_RNIJ7QO_LC_12_17_2.LUT_INIT=16'b0010001000000000;
    LogicCell40 un4_sacqtime_cry_23_c_RNIJ7QO_LC_12_17_2 (
            .in0(N__31935),
            .in1(N__29699),
            .in2(_gnd_net_),
            .in3(N__32180),
            .lcout(N_31_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sRAM_ADD_1_LC_12_17_3.C_ON=1'b0;
    defparam sRAM_ADD_1_LC_12_17_3.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_1_LC_12_17_3.LUT_INIT=16'b1110010011001100;
    LogicCell40 sRAM_ADD_1_LC_12_17_3 (
            .in0(N__32183),
            .in1(N__29688),
            .in2(N__31605),
            .in3(N__31941),
            .lcout(RAM_ADD_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47816),
            .ce(N__30262),
            .sr(_gnd_net_));
    defparam sRAM_ADD_10_LC_12_17_4.C_ON=1'b0;
    defparam sRAM_ADD_10_LC_12_17_4.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_10_LC_12_17_4.LUT_INIT=16'b1101100011110000;
    LogicCell40 sRAM_ADD_10_LC_12_17_4 (
            .in0(N__31937),
            .in1(N__33096),
            .in2(N__29646),
            .in3(N__32185),
            .lcout(RAM_ADD_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47816),
            .ce(N__30262),
            .sr(_gnd_net_));
    defparam sRAM_ADD_11_LC_12_17_5.C_ON=1'b0;
    defparam sRAM_ADD_11_LC_12_17_5.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_11_LC_12_17_5.LUT_INIT=16'b1110010011001100;
    LogicCell40 sRAM_ADD_11_LC_12_17_5 (
            .in0(N__32181),
            .in1(N__30405),
            .in2(N__33078),
            .in3(N__31939),
            .lcout(RAM_ADD_c_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47816),
            .ce(N__30262),
            .sr(_gnd_net_));
    defparam sRAM_ADD_12_LC_12_17_6.C_ON=1'b0;
    defparam sRAM_ADD_12_LC_12_17_6.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_12_LC_12_17_6.LUT_INIT=16'b1101100011110000;
    LogicCell40 sRAM_ADD_12_LC_12_17_6 (
            .in0(N__31938),
            .in1(N__33057),
            .in2(N__30354),
            .in3(N__32186),
            .lcout(RAM_ADD_c_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47816),
            .ce(N__30262),
            .sr(_gnd_net_));
    defparam sRAM_ADD_13_LC_12_17_7.C_ON=1'b0;
    defparam sRAM_ADD_13_LC_12_17_7.SEQ_MODE=4'b1000;
    defparam sRAM_ADD_13_LC_12_17_7.LUT_INIT=16'b1110010011001100;
    LogicCell40 sRAM_ADD_13_LC_12_17_7 (
            .in0(N__32182),
            .in1(N__30309),
            .in2(N__33036),
            .in3(N__31940),
            .lcout(RAM_ADD_c_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47816),
            .ce(N__30262),
            .sr(_gnd_net_));
    defparam RAM_DATA_1_3_LC_12_18_0.C_ON=1'b0;
    defparam RAM_DATA_1_3_LC_12_18_0.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_3_LC_12_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_3_LC_12_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30240),
            .lcout(RAM_DATA_1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(N__31181),
            .sr(N__52970));
    defparam RAM_DATA_1_0_LC_12_18_1.C_ON=1'b0;
    defparam RAM_DATA_1_0_LC_12_18_1.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_0_LC_12_18_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 RAM_DATA_1_0_LC_12_18_1 (
            .in0(N__30204),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RAM_DATA_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(N__31181),
            .sr(N__52970));
    defparam RAM_DATA_1_5_LC_12_18_2.C_ON=1'b0;
    defparam RAM_DATA_1_5_LC_12_18_2.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_5_LC_12_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_5_LC_12_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30165),
            .lcout(RAM_DATA_1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(N__31181),
            .sr(N__52970));
    defparam RAM_DATA_1_1_LC_12_18_3.C_ON=1'b0;
    defparam RAM_DATA_1_1_LC_12_18_3.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_1_LC_12_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_1_LC_12_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30123),
            .lcout(RAM_DATA_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(N__31181),
            .sr(N__52970));
    defparam RAM_DATA_1_8_LC_12_18_4.C_ON=1'b0;
    defparam RAM_DATA_1_8_LC_12_18_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_8_LC_12_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_8_LC_12_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30090),
            .lcout(RAM_DATA_1Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(N__31181),
            .sr(N__52970));
    defparam RAM_DATA_1_9_LC_12_18_5.C_ON=1'b0;
    defparam RAM_DATA_1_9_LC_12_18_5.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_9_LC_12_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_9_LC_12_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30639),
            .lcout(RAM_DATA_1Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(N__31181),
            .sr(N__52970));
    defparam RAM_DATA_1_15_LC_12_18_6.C_ON=1'b0;
    defparam RAM_DATA_1_15_LC_12_18_6.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_15_LC_12_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_15_LC_12_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37903),
            .lcout(RAM_DATA_1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(N__31181),
            .sr(N__52970));
    defparam RAM_DATA_1_7_LC_12_18_7.C_ON=1'b0;
    defparam RAM_DATA_1_7_LC_12_18_7.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_7_LC_12_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_7_LC_12_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(RAM_DATA_1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47824),
            .ce(N__31181),
            .sr(N__52970));
    defparam RAM_DATA_cl_1_RNO_0_15_LC_12_19_1.C_ON=1'b0;
    defparam RAM_DATA_cl_1_RNO_0_15_LC_12_19_1.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_1_RNO_0_15_LC_12_19_1.LUT_INIT=16'b0101010100000000;
    LogicCell40 RAM_DATA_cl_1_RNO_0_15_LC_12_19_1 (
            .in0(N__30539),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31711),
            .lcout(N_100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_13_RNO_0_15_LC_12_19_3.C_ON=1'b0;
    defparam RAM_DATA_cl_13_RNO_0_15_LC_12_19_3.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_13_RNO_0_15_LC_12_19_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 RAM_DATA_cl_13_RNO_0_15_LC_12_19_3 (
            .in0(_gnd_net_),
            .in1(N__30503),
            .in2(_gnd_net_),
            .in3(N__31710),
            .lcout(N_97),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_3_RNO_0_15_LC_12_19_5.C_ON=1'b0;
    defparam RAM_DATA_cl_3_RNO_0_15_LC_12_19_5.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_3_RNO_0_15_LC_12_19_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 RAM_DATA_cl_3_RNO_0_15_LC_12_19_5 (
            .in0(_gnd_net_),
            .in1(N__30431),
            .in2(_gnd_net_),
            .in3(N__31713),
            .lcout(N_103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_2_RNO_0_15_LC_12_19_7.C_ON=1'b0;
    defparam RAM_DATA_cl_2_RNO_0_15_LC_12_19_7.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_2_RNO_0_15_LC_12_19_7.LUT_INIT=16'b0011001100000000;
    LogicCell40 RAM_DATA_cl_2_RNO_0_15_LC_12_19_7 (
            .in0(_gnd_net_),
            .in1(N__30470),
            .in2(_gnd_net_),
            .in3(N__31712),
            .lcout(N_101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_3_15_LC_12_20_2.C_ON=1'b0;
    defparam RAM_DATA_cl_3_15_LC_12_20_2.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_3_15_LC_12_20_2.LUT_INIT=16'b0100000000000000;
    LogicCell40 RAM_DATA_cl_3_15_LC_12_20_2 (
            .in0(N__30453),
            .in1(N__32153),
            .in2(N__32675),
            .in3(N__31973),
            .lcout(RAM_DATA_cl_3Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47841),
            .ce(),
            .sr(N__52967));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_0_LC_13_2_3 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_0_LC_13_2_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_0_LC_13_2_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_0_LC_13_2_3  (
            .in0(N__38552),
            .in1(N__52592),
            .in2(_gnd_net_),
            .in3(N__30420),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30697),
            .ce(N__30672),
            .sr(N__53110));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_5_LC_13_3_0 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_5_LC_13_3_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_5_LC_13_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_5_LC_13_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30746),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30700),
            .ce(N__30671),
            .sr(N__53097));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_1_LC_13_3_1 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_1_LC_13_3_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_1_LC_13_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_1_LC_13_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30794),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30700),
            .ce(N__30671),
            .sr(N__53097));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_2_LC_13_3_2 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_2_LC_13_3_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_2_LC_13_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_2_LC_13_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30782),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30700),
            .ce(N__30671),
            .sr(N__53097));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_3_LC_13_3_3 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_3_LC_13_3_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_3_LC_13_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_3_LC_13_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30770),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30700),
            .ce(N__30671),
            .sr(N__53097));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_4_LC_13_3_4 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_4_LC_13_3_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_4_LC_13_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_4_LC_13_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30758),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30700),
            .ce(N__30671),
            .sr(N__53097));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_6_LC_13_3_5 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_6_LC_13_3_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_6_LC_13_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_6_LC_13_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30734),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30700),
            .ce(N__30671),
            .sr(N__53097));
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_7_LC_13_3_7 .C_ON=1'b0;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_7_LC_13_3_7 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.rx_shift_data_pos_sclk_i_7_LC_13_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \spi_slave_inst.rx_shift_data_pos_sclk_i_7_LC_13_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30722),
            .lcout(\spi_slave_inst.rx_shift_data_pos_sclk_iZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30700),
            .ce(N__30671),
            .sr(N__53097));
    defparam sDAC_mem_38_1_LC_13_4_0.C_ON=1'b0;
    defparam sDAC_mem_38_1_LC_13_4_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_1_LC_13_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_1_LC_13_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50422),
            .lcout(sDAC_mem_38Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47817),
            .ce(N__41868),
            .sr(N__53084));
    defparam sDAC_mem_6_2_LC_13_5_0.C_ON=1'b0;
    defparam sDAC_mem_6_2_LC_13_5_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_2_LC_13_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_2_LC_13_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50005),
            .lcout(sDAC_mem_6Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47808),
            .ce(N__43078),
            .sr(N__53072));
    defparam sDAC_mem_6_5_LC_13_5_1.C_ON=1'b0;
    defparam sDAC_mem_6_5_LC_13_5_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_5_LC_13_5_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_6_5_LC_13_5_1 (
            .in0(N__46793),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_6Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47808),
            .ce(N__43078),
            .sr(N__53072));
    defparam sDAC_mem_6_7_LC_13_5_2.C_ON=1'b0;
    defparam sDAC_mem_6_7_LC_13_5_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_7_LC_13_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_7_LC_13_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48671),
            .lcout(sDAC_mem_6Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47808),
            .ce(N__43078),
            .sr(N__53072));
    defparam sDAC_mem_2_0_LC_13_6_0.C_ON=1'b0;
    defparam sDAC_mem_2_0_LC_13_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_0_LC_13_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_0_LC_13_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51024),
            .lcout(sDAC_mem_2Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47797),
            .ce(N__37407),
            .sr(N__53060));
    defparam sDAC_mem_2_1_LC_13_6_1.C_ON=1'b0;
    defparam sDAC_mem_2_1_LC_13_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_1_LC_13_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_1_LC_13_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50625),
            .lcout(sDAC_mem_2Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47797),
            .ce(N__37407),
            .sr(N__53060));
    defparam sDAC_mem_2_2_LC_13_6_2.C_ON=1'b0;
    defparam sDAC_mem_2_2_LC_13_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_2_LC_13_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_2_LC_13_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50006),
            .lcout(sDAC_mem_2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47797),
            .ce(N__37407),
            .sr(N__53060));
    defparam sDAC_mem_2_3_LC_13_6_3.C_ON=1'b0;
    defparam sDAC_mem_2_3_LC_13_6_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_3_LC_13_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_3_LC_13_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49496),
            .lcout(sDAC_mem_2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47797),
            .ce(N__37407),
            .sr(N__53060));
    defparam sDAC_mem_2_4_LC_13_6_4.C_ON=1'b0;
    defparam sDAC_mem_2_4_LC_13_6_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_4_LC_13_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_4_LC_13_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48989),
            .lcout(sDAC_mem_2Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47797),
            .ce(N__37407),
            .sr(N__53060));
    defparam sDAC_mem_2_5_LC_13_6_5.C_ON=1'b0;
    defparam sDAC_mem_2_5_LC_13_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_5_LC_13_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_5_LC_13_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46794),
            .lcout(sDAC_mem_2Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47797),
            .ce(N__37407),
            .sr(N__53060));
    defparam sDAC_mem_2_6_LC_13_6_6.C_ON=1'b0;
    defparam sDAC_mem_2_6_LC_13_6_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_6_LC_13_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_6_LC_13_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48062),
            .lcout(sDAC_mem_2Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47797),
            .ce(N__37407),
            .sr(N__53060));
    defparam sDAC_mem_2_7_LC_13_6_7.C_ON=1'b0;
    defparam sDAC_mem_2_7_LC_13_6_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_2_7_LC_13_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_2_7_LC_13_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48670),
            .lcout(sDAC_mem_2Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47797),
            .ce(N__37407),
            .sr(N__53060));
    defparam sDAC_mem_22_1_LC_13_7_1.C_ON=1'b0;
    defparam sDAC_mem_22_1_LC_13_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_1_LC_13_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_1_LC_13_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50691),
            .lcout(sDAC_mem_22Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47782),
            .ce(N__39824),
            .sr(N__53050));
    defparam sDAC_data_RNO_21_5_LC_13_7_2.C_ON=1'b0;
    defparam sDAC_data_RNO_21_5_LC_13_7_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_5_LC_13_7_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_5_LC_13_7_2 (
            .in0(N__52007),
            .in1(N__30849),
            .in2(_gnd_net_),
            .in3(N__30843),
            .lcout(sDAC_data_RNO_21Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_22_2_LC_13_7_3.C_ON=1'b0;
    defparam sDAC_mem_22_2_LC_13_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_2_LC_13_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_2_LC_13_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50091),
            .lcout(sDAC_mem_22Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47782),
            .ce(N__39824),
            .sr(N__53050));
    defparam sDAC_data_RNO_21_6_LC_13_7_4.C_ON=1'b0;
    defparam sDAC_data_RNO_21_6_LC_13_7_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_6_LC_13_7_4.LUT_INIT=16'b1010111110100000;
    LogicCell40 sDAC_data_RNO_21_6_LC_13_7_4 (
            .in0(N__30837),
            .in1(_gnd_net_),
            .in2(N__52118),
            .in3(N__30831),
            .lcout(sDAC_data_RNO_21Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_22_3_LC_13_7_5.C_ON=1'b0;
    defparam sDAC_mem_22_3_LC_13_7_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_3_LC_13_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_3_LC_13_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49590),
            .lcout(sDAC_mem_22Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47782),
            .ce(N__39824),
            .sr(N__53050));
    defparam sDAC_data_RNO_21_7_LC_13_7_6.C_ON=1'b0;
    defparam sDAC_data_RNO_21_7_LC_13_7_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_7_LC_13_7_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_7_LC_13_7_6 (
            .in0(N__52008),
            .in1(N__30825),
            .in2(_gnd_net_),
            .in3(N__30819),
            .lcout(sDAC_data_RNO_21Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_22_4_LC_13_7_7.C_ON=1'b0;
    defparam sDAC_mem_22_4_LC_13_7_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_4_LC_13_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_4_LC_13_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49077),
            .lcout(sDAC_mem_22Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47782),
            .ce(N__39824),
            .sr(N__53050));
    defparam sAddress_RNIAM2A_3_LC_13_8_0.C_ON=1'b0;
    defparam sAddress_RNIAM2A_3_LC_13_8_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNIAM2A_3_LC_13_8_0.LUT_INIT=16'b0000000000010001;
    LogicCell40 sAddress_RNIAM2A_3_LC_13_8_0 (
            .in0(N__46438),
            .in1(N__40534),
            .in2(_gnd_net_),
            .in3(N__40347),
            .lcout(N_291),
            .ltout(N_291_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_6_LC_13_8_1.C_ON=1'b0;
    defparam sAddress_RNI9IH12_6_LC_13_8_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_6_LC_13_8_1.LUT_INIT=16'b1100000000000000;
    LogicCell40 sAddress_RNI9IH12_6_LC_13_8_1 (
            .in0(_gnd_net_),
            .in1(N__30906),
            .in2(N__30813),
            .in3(N__44730),
            .lcout(sEEPonPoff_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_20_3_LC_13_8_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_20_3_LC_13_8_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_20_3_LC_13_8_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 sAddress_RNI9IH12_20_3_LC_13_8_2 (
            .in0(_gnd_net_),
            .in1(N__30871),
            .in2(_gnd_net_),
            .in3(N__43160),
            .lcout(sDAC_mem_17_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_0_5_LC_13_8_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_0_5_LC_13_8_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_0_5_LC_13_8_3.LUT_INIT=16'b0010001000000000;
    LogicCell40 sAddress_RNI9IH12_0_5_LC_13_8_3 (
            .in0(N__30870),
            .in1(N__46512),
            .in2(_gnd_net_),
            .in3(N__46328),
            .lcout(sDAC_mem_1_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_2_LC_13_8_4.C_ON=1'b0;
    defparam sAddress_RNIA6242_2_LC_13_8_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_2_LC_13_8_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 sAddress_RNIA6242_2_LC_13_8_4 (
            .in0(N__44957),
            .in1(N__40348),
            .in2(N__40555),
            .in3(N__30996),
            .lcout(sAddress_RNIA6242Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIQ63A_0_6_LC_13_8_5.C_ON=1'b0;
    defparam sAddress_RNIQ63A_0_6_LC_13_8_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNIQ63A_0_6_LC_13_8_5.LUT_INIT=16'b0010000000000000;
    LogicCell40 sAddress_RNIQ63A_0_6_LC_13_8_5 (
            .in0(N__30954),
            .in1(N__46511),
            .in2(N__30933),
            .in3(N__44644),
            .lcout(sEEPonPoff_1_sqmuxa_0_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_21_3_LC_13_8_6.C_ON=1'b0;
    defparam sAddress_RNI9IH12_21_3_LC_13_8_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_21_3_LC_13_8_6.LUT_INIT=16'b0000000010001000;
    LogicCell40 sAddress_RNI9IH12_21_3_LC_13_8_6 (
            .in0(N__44731),
            .in1(N__30873),
            .in2(_gnd_net_),
            .in3(N__31105),
            .lcout(sEEPon_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_5_LC_13_8_7.C_ON=1'b0;
    defparam sAddress_RNI9IH12_5_LC_13_8_7.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_5_LC_13_8_7.LUT_INIT=16'b1000100000000000;
    LogicCell40 sAddress_RNI9IH12_5_LC_13_8_7 (
            .in0(N__30872),
            .in1(N__46513),
            .in2(_gnd_net_),
            .in3(N__46329),
            .lcout(sDAC_mem_33_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_17_0_LC_13_9_0.C_ON=1'b0;
    defparam sDAC_mem_17_0_LC_13_9_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_0_LC_13_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_0_LC_13_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51027),
            .lcout(sDAC_mem_17Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47756),
            .ce(N__30960),
            .sr(N__53031));
    defparam sDAC_mem_17_1_LC_13_9_1.C_ON=1'b0;
    defparam sDAC_mem_17_1_LC_13_9_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_1_LC_13_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_1_LC_13_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50693),
            .lcout(sDAC_mem_17Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47756),
            .ce(N__30960),
            .sr(N__53031));
    defparam sDAC_mem_17_2_LC_13_9_2.C_ON=1'b0;
    defparam sDAC_mem_17_2_LC_13_9_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_2_LC_13_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_2_LC_13_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50092),
            .lcout(sDAC_mem_17Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47756),
            .ce(N__30960),
            .sr(N__53031));
    defparam sDAC_mem_17_3_LC_13_9_3.C_ON=1'b0;
    defparam sDAC_mem_17_3_LC_13_9_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_3_LC_13_9_3.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_17_3_LC_13_9_3 (
            .in0(_gnd_net_),
            .in1(N__49591),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_17Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47756),
            .ce(N__30960),
            .sr(N__53031));
    defparam sDAC_mem_17_4_LC_13_9_4.C_ON=1'b0;
    defparam sDAC_mem_17_4_LC_13_9_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_4_LC_13_9_4.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_17_4_LC_13_9_4 (
            .in0(_gnd_net_),
            .in1(N__49075),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_17Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47756),
            .ce(N__30960),
            .sr(N__53031));
    defparam sDAC_mem_17_5_LC_13_9_5.C_ON=1'b0;
    defparam sDAC_mem_17_5_LC_13_9_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_5_LC_13_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_5_LC_13_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46897),
            .lcout(sDAC_mem_17Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47756),
            .ce(N__30960),
            .sr(N__53031));
    defparam sDAC_mem_17_6_LC_13_9_6.C_ON=1'b0;
    defparam sDAC_mem_17_6_LC_13_9_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_6_LC_13_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_6_LC_13_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48124),
            .lcout(sDAC_mem_17Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47756),
            .ce(N__30960),
            .sr(N__53031));
    defparam sDAC_mem_17_7_LC_13_9_7.C_ON=1'b0;
    defparam sDAC_mem_17_7_LC_13_9_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_17_7_LC_13_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_17_7_LC_13_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48668),
            .lcout(sDAC_mem_17Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47756),
            .ce(N__30960),
            .sr(N__53031));
    defparam sDAC_mem_32_0_LC_13_10_0.C_ON=1'b0;
    defparam sDAC_mem_32_0_LC_13_10_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_0_LC_13_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_0_LC_13_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51132),
            .lcout(sDAC_mem_32Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47742),
            .ce(N__31113),
            .sr(N__53021));
    defparam sDAC_mem_32_1_LC_13_10_1.C_ON=1'b0;
    defparam sDAC_mem_32_1_LC_13_10_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_1_LC_13_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_1_LC_13_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50694),
            .lcout(sDAC_mem_32Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47742),
            .ce(N__31113),
            .sr(N__53021));
    defparam sDAC_mem_32_2_LC_13_10_2.C_ON=1'b0;
    defparam sDAC_mem_32_2_LC_13_10_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_2_LC_13_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_2_LC_13_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50093),
            .lcout(sDAC_mem_32Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47742),
            .ce(N__31113),
            .sr(N__53021));
    defparam sDAC_mem_32_3_LC_13_10_3.C_ON=1'b0;
    defparam sDAC_mem_32_3_LC_13_10_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_3_LC_13_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_3_LC_13_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49592),
            .lcout(sDAC_mem_32Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47742),
            .ce(N__31113),
            .sr(N__53021));
    defparam sDAC_mem_32_4_LC_13_10_4.C_ON=1'b0;
    defparam sDAC_mem_32_4_LC_13_10_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_4_LC_13_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_4_LC_13_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49078),
            .lcout(sDAC_mem_32Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47742),
            .ce(N__31113),
            .sr(N__53021));
    defparam sDAC_mem_32_5_LC_13_10_5.C_ON=1'b0;
    defparam sDAC_mem_32_5_LC_13_10_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_5_LC_13_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_5_LC_13_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46898),
            .lcout(sDAC_mem_32Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47742),
            .ce(N__31113),
            .sr(N__53021));
    defparam sDAC_mem_32_6_LC_13_10_6.C_ON=1'b0;
    defparam sDAC_mem_32_6_LC_13_10_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_6_LC_13_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_6_LC_13_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48254),
            .lcout(sDAC_mem_32Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47742),
            .ce(N__31113),
            .sr(N__53021));
    defparam sDAC_mem_32_7_LC_13_10_7.C_ON=1'b0;
    defparam sDAC_mem_32_7_LC_13_10_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_32_7_LC_13_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_32_7_LC_13_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48669),
            .lcout(sDAC_mem_32Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47742),
            .ce(N__31113),
            .sr(N__53021));
    defparam sAddress_RNI9IH12_0_6_LC_13_11_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_0_6_LC_13_11_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_0_6_LC_13_11_0.LUT_INIT=16'b0000000000100000;
    LogicCell40 sAddress_RNI9IH12_0_6_LC_13_11_0 (
            .in0(N__44694),
            .in1(N__46096),
            .in2(N__44595),
            .in3(N__31104),
            .lcout(sEETrigCounter_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI5B15_3_LC_13_11_1.C_ON=1'b0;
    defparam sAddress_RNI5B15_3_LC_13_11_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI5B15_3_LC_13_11_1.LUT_INIT=16'b1111111100110011;
    LogicCell40 sAddress_RNI5B15_3_LC_13_11_1 (
            .in0(_gnd_net_),
            .in1(N__40495),
            .in2(_gnd_net_),
            .in3(N__40304),
            .lcout(N_1480),
            .ltout(N_1480_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_7_1_LC_13_11_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_7_1_LC_13_11_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_7_1_LC_13_11_2.LUT_INIT=16'b0000100000001000;
    LogicCell40 sAddress_RNI9IH12_7_1_LC_13_11_2 (
            .in0(N__43139),
            .in1(N__44592),
            .in2(N__30999),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_31_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_9_3_LC_13_11_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_9_3_LC_13_11_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_9_3_LC_13_11_3.LUT_INIT=16'b0000010000000000;
    LogicCell40 sAddress_RNI9IH12_9_3_LC_13_11_3 (
            .in0(N__40512),
            .in1(N__40306),
            .in2(N__46450),
            .in3(N__43140),
            .lcout(sDAC_mem_18_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIA6242_2_2_LC_13_11_4.C_ON=1'b0;
    defparam sAddress_RNIA6242_2_2_LC_13_11_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNIA6242_2_2_LC_13_11_4.LUT_INIT=16'b0000000100000000;
    LogicCell40 sAddress_RNIA6242_2_2_LC_13_11_4 (
            .in0(N__40305),
            .in1(N__44960),
            .in2(N__40533),
            .in3(N__30992),
            .lcout(sAddress_RNIA6242_2Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIVREN1_0_4_LC_13_11_5.C_ON=1'b0;
    defparam sAddress_RNIVREN1_0_4_LC_13_11_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNIVREN1_0_4_LC_13_11_5.LUT_INIT=16'b0010000000000000;
    LogicCell40 sAddress_RNIVREN1_0_4_LC_13_11_5 (
            .in0(N__46486),
            .in1(N__44637),
            .in2(N__44797),
            .in3(N__44693),
            .lcout(N_280),
            .ltout(N_280_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_3_3_LC_13_11_6.C_ON=1'b0;
    defparam sAddress_RNI9IH12_3_3_LC_13_11_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_3_3_LC_13_11_6.LUT_INIT=16'b0010000000000000;
    LogicCell40 sAddress_RNI9IH12_3_3_LC_13_11_6 (
            .in0(N__44588),
            .in1(N__40511),
            .in2(N__30963),
            .in3(N__40335),
            .lcout(sDAC_mem_24_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_14_3_LC_13_11_7.C_ON=1'b0;
    defparam sAddress_RNI9IH12_14_3_LC_13_11_7.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_14_3_LC_13_11_7.LUT_INIT=16'b0000010000000000;
    LogicCell40 sAddress_RNI9IH12_14_3_LC_13_11_7 (
            .in0(N__40336),
            .in1(N__43269),
            .in2(N__40540),
            .in3(N__43138),
            .lcout(sDAC_mem_19_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_19_0_LC_13_12_0.C_ON=1'b0;
    defparam sDAC_mem_19_0_LC_13_12_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_0_LC_13_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_0_LC_13_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51134),
            .lcout(sDAC_mem_19Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47743),
            .ce(N__31122),
            .sr(N__53010));
    defparam sDAC_mem_19_1_LC_13_12_1.C_ON=1'b0;
    defparam sDAC_mem_19_1_LC_13_12_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_1_LC_13_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_1_LC_13_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50574),
            .lcout(sDAC_mem_19Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47743),
            .ce(N__31122),
            .sr(N__53010));
    defparam sDAC_mem_19_2_LC_13_12_2.C_ON=1'b0;
    defparam sDAC_mem_19_2_LC_13_12_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_2_LC_13_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_2_LC_13_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50179),
            .lcout(sDAC_mem_19Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47743),
            .ce(N__31122),
            .sr(N__53010));
    defparam sDAC_mem_19_3_LC_13_12_3.C_ON=1'b0;
    defparam sDAC_mem_19_3_LC_13_12_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_3_LC_13_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_3_LC_13_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49702),
            .lcout(sDAC_mem_19Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47743),
            .ce(N__31122),
            .sr(N__53010));
    defparam sDAC_mem_19_4_LC_13_12_4.C_ON=1'b0;
    defparam sDAC_mem_19_4_LC_13_12_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_4_LC_13_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_4_LC_13_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49145),
            .lcout(sDAC_mem_19Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47743),
            .ce(N__31122),
            .sr(N__53010));
    defparam sDAC_mem_19_5_LC_13_12_5.C_ON=1'b0;
    defparam sDAC_mem_19_5_LC_13_12_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_5_LC_13_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_5_LC_13_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46993),
            .lcout(sDAC_mem_19Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47743),
            .ce(N__31122),
            .sr(N__53010));
    defparam sDAC_mem_19_6_LC_13_12_6.C_ON=1'b0;
    defparam sDAC_mem_19_6_LC_13_12_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_6_LC_13_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_6_LC_13_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48236),
            .lcout(sDAC_mem_19Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47743),
            .ce(N__31122),
            .sr(N__53010));
    defparam sDAC_mem_19_7_LC_13_12_7.C_ON=1'b0;
    defparam sDAC_mem_19_7_LC_13_12_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_19_7_LC_13_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_19_7_LC_13_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48817),
            .lcout(sDAC_mem_19Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47743),
            .ce(N__31122),
            .sr(N__53010));
    defparam sDAC_mem_18_3_LC_13_13_1.C_ON=1'b0;
    defparam sDAC_mem_18_3_LC_13_13_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_3_LC_13_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_3_LC_13_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49703),
            .lcout(sDAC_mem_18Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47757),
            .ce(N__34089),
            .sr(N__53002));
    defparam sDAC_data_RNO_30_7_LC_13_13_2.C_ON=1'b0;
    defparam sDAC_data_RNO_30_7_LC_13_13_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_7_LC_13_13_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_30_7_LC_13_13_2 (
            .in0(N__52150),
            .in1(N__31152),
            .in2(_gnd_net_),
            .in3(N__31158),
            .lcout(sDAC_data_RNO_30Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_18_4_LC_13_13_3.C_ON=1'b0;
    defparam sDAC_mem_18_4_LC_13_13_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_4_LC_13_13_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_18_4_LC_13_13_3 (
            .in0(N__49307),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_18Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47757),
            .ce(N__34089),
            .sr(N__53002));
    defparam sDAC_data_RNO_30_8_LC_13_13_4.C_ON=1'b0;
    defparam sDAC_data_RNO_30_8_LC_13_13_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_8_LC_13_13_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_30_8_LC_13_13_4 (
            .in0(N__52151),
            .in1(N__31140),
            .in2(_gnd_net_),
            .in3(N__31146),
            .lcout(sDAC_data_RNO_30Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_18_5_LC_13_13_5.C_ON=1'b0;
    defparam sDAC_mem_18_5_LC_13_13_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_5_LC_13_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_5_LC_13_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46994),
            .lcout(sDAC_mem_18Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47757),
            .ce(N__34089),
            .sr(N__53002));
    defparam sDAC_data_RNO_30_9_LC_13_13_6.C_ON=1'b0;
    defparam sDAC_data_RNO_30_9_LC_13_13_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_9_LC_13_13_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_30_9_LC_13_13_6 (
            .in0(N__52152),
            .in1(N__31128),
            .in2(_gnd_net_),
            .in3(N__31134),
            .lcout(sDAC_data_RNO_30Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_18_6_LC_13_13_7.C_ON=1'b0;
    defparam sDAC_mem_18_6_LC_13_13_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_6_LC_13_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_6_LC_13_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48237),
            .lcout(sDAC_mem_18Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47757),
            .ce(N__34089),
            .sr(N__53002));
    defparam sDAC_mem_24_0_LC_13_14_0.C_ON=1'b0;
    defparam sDAC_mem_24_0_LC_13_14_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_0_LC_13_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_0_LC_13_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51216),
            .lcout(sDAC_mem_24Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47768),
            .ce(N__39954),
            .sr(N__52993));
    defparam sDAC_mem_24_1_LC_13_14_1.C_ON=1'b0;
    defparam sDAC_mem_24_1_LC_13_14_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_1_LC_13_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_1_LC_13_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50732),
            .lcout(sDAC_mem_24Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47768),
            .ce(N__39954),
            .sr(N__52993));
    defparam sDAC_mem_24_3_LC_13_14_2.C_ON=1'b0;
    defparam sDAC_mem_24_3_LC_13_14_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_3_LC_13_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_3_LC_13_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49704),
            .lcout(sDAC_mem_24Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47768),
            .ce(N__39954),
            .sr(N__52993));
    defparam sDAC_mem_24_4_LC_13_14_3.C_ON=1'b0;
    defparam sDAC_mem_24_4_LC_13_14_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_4_LC_13_14_3.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_24_4_LC_13_14_3 (
            .in0(_gnd_net_),
            .in1(N__49144),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_24Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47768),
            .ce(N__39954),
            .sr(N__52993));
    defparam sDAC_mem_24_6_LC_13_14_4.C_ON=1'b0;
    defparam sDAC_mem_24_6_LC_13_14_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_6_LC_13_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_6_LC_13_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48303),
            .lcout(sDAC_mem_24Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47768),
            .ce(N__39954),
            .sr(N__52993));
    defparam sEEACQ_10_LC_13_15_0.C_ON=1'b0;
    defparam sEEACQ_10_LC_13_15_0.SEQ_MODE=4'b1010;
    defparam sEEACQ_10_LC_13_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_10_LC_13_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50257),
            .lcout(sEEACQZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47783),
            .ce(N__31170),
            .sr(N__52988));
    defparam sEEACQ_11_LC_13_15_1.C_ON=1'b0;
    defparam sEEACQ_11_LC_13_15_1.SEQ_MODE=4'b1010;
    defparam sEEACQ_11_LC_13_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_11_LC_13_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49786),
            .lcout(sEEACQZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47783),
            .ce(N__31170),
            .sr(N__52988));
    defparam sEEACQ_12_LC_13_15_2.C_ON=1'b0;
    defparam sEEACQ_12_LC_13_15_2.SEQ_MODE=4'b1011;
    defparam sEEACQ_12_LC_13_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_12_LC_13_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49226),
            .lcout(sEEACQZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47783),
            .ce(N__31170),
            .sr(N__52988));
    defparam sEEACQ_13_LC_13_15_3.C_ON=1'b0;
    defparam sEEACQ_13_LC_13_15_3.SEQ_MODE=4'b1011;
    defparam sEEACQ_13_LC_13_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_13_LC_13_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47119),
            .lcout(sEEACQZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47783),
            .ce(N__31170),
            .sr(N__52988));
    defparam sEEACQ_14_LC_13_15_4.C_ON=1'b0;
    defparam sEEACQ_14_LC_13_15_4.SEQ_MODE=4'b1010;
    defparam sEEACQ_14_LC_13_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_14_LC_13_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48304),
            .lcout(sEEACQZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47783),
            .ce(N__31170),
            .sr(N__52988));
    defparam sEEACQ_15_LC_13_15_5.C_ON=1'b0;
    defparam sEEACQ_15_LC_13_15_5.SEQ_MODE=4'b1010;
    defparam sEEACQ_15_LC_13_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_15_LC_13_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48667),
            .lcout(sEEACQZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47783),
            .ce(N__31170),
            .sr(N__52988));
    defparam sEEACQ_8_LC_13_15_6.C_ON=1'b0;
    defparam sEEACQ_8_LC_13_15_6.SEQ_MODE=4'b1010;
    defparam sEEACQ_8_LC_13_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_8_LC_13_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51262),
            .lcout(sEEACQZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47783),
            .ce(N__31170),
            .sr(N__52988));
    defparam sEEACQ_9_LC_13_15_7.C_ON=1'b0;
    defparam sEEACQ_9_LC_13_15_7.SEQ_MODE=4'b1011;
    defparam sEEACQ_9_LC_13_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEACQ_9_LC_13_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50734),
            .lcout(sEEACQZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47783),
            .ce(N__31170),
            .sr(N__52988));
    defparam RAM_DATA_1_4_LC_13_16_0.C_ON=1'b0;
    defparam RAM_DATA_1_4_LC_13_16_0.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_4_LC_13_16_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 RAM_DATA_1_4_LC_13_16_0 (
            .in0(N__31590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RAM_DATA_1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47798),
            .ce(N__31182),
            .sr(N__52983));
    defparam RAM_DATA_1_6_LC_13_16_1.C_ON=1'b0;
    defparam RAM_DATA_1_6_LC_13_16_1.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_6_LC_13_16_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 RAM_DATA_1_6_LC_13_16_1 (
            .in0(N__31554),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RAM_DATA_1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47798),
            .ce(N__31182),
            .sr(N__52983));
    defparam RAM_DATA_1_10_LC_13_16_2.C_ON=1'b0;
    defparam RAM_DATA_1_10_LC_13_16_2.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_10_LC_13_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_10_LC_13_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31521),
            .lcout(RAM_DATA_1Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47798),
            .ce(N__31182),
            .sr(N__52983));
    defparam RAM_DATA_1_11_LC_13_16_3.C_ON=1'b0;
    defparam RAM_DATA_1_11_LC_13_16_3.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_11_LC_13_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_11_LC_13_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31476),
            .lcout(RAM_DATA_1Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47798),
            .ce(N__31182),
            .sr(N__52983));
    defparam RAM_DATA_1_12_LC_13_16_4.C_ON=1'b0;
    defparam RAM_DATA_1_12_LC_13_16_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_12_LC_13_16_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 RAM_DATA_1_12_LC_13_16_4 (
            .in0(N__31434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RAM_DATA_1Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47798),
            .ce(N__31182),
            .sr(N__52983));
    defparam RAM_DATA_1_13_LC_13_16_5.C_ON=1'b0;
    defparam RAM_DATA_1_13_LC_13_16_5.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_13_LC_13_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_13_LC_13_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31389),
            .lcout(RAM_DATA_1Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47798),
            .ce(N__31182),
            .sr(N__52983));
    defparam RAM_DATA_1_14_LC_13_16_6.C_ON=1'b0;
    defparam RAM_DATA_1_14_LC_13_16_6.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_14_LC_13_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_14_LC_13_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31301),
            .lcout(RAM_DATA_1Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47798),
            .ce(N__31182),
            .sr(N__52983));
    defparam RAM_DATA_1_2_LC_13_16_7.C_ON=1'b0;
    defparam RAM_DATA_1_2_LC_13_16_7.SEQ_MODE=4'b1010;
    defparam RAM_DATA_1_2_LC_13_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 RAM_DATA_1_2_LC_13_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31215),
            .lcout(RAM_DATA_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47798),
            .ce(N__31182),
            .sr(N__52983));
    defparam RAM_DATA_cl_4_15_LC_13_17_0.C_ON=1'b0;
    defparam RAM_DATA_cl_4_15_LC_13_17_0.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_4_15_LC_13_17_0.LUT_INIT=16'b0100000000000000;
    LogicCell40 RAM_DATA_cl_4_15_LC_13_17_0 (
            .in0(N__31629),
            .in1(N__32222),
            .in2(N__32546),
            .in3(N__31945),
            .lcout(RAM_DATA_cl_4Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47809),
            .ce(),
            .sr(N__52980));
    defparam RAM_DATA_cl_5_RNO_0_15_LC_13_17_1.C_ON=1'b0;
    defparam RAM_DATA_cl_5_RNO_0_15_LC_13_17_1.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_5_RNO_0_15_LC_13_17_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 RAM_DATA_cl_5_RNO_0_15_LC_13_17_1 (
            .in0(_gnd_net_),
            .in1(N__32735),
            .in2(_gnd_net_),
            .in3(N__31695),
            .lcout(),
            .ltout(N_107_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_5_15_LC_13_17_2.C_ON=1'b0;
    defparam RAM_DATA_cl_5_15_LC_13_17_2.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_5_15_LC_13_17_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 RAM_DATA_cl_5_15_LC_13_17_2 (
            .in0(N__32493),
            .in1(N__32223),
            .in2(N__32757),
            .in3(N__31946),
            .lcout(RAM_DATA_cl_5Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47809),
            .ce(),
            .sr(N__52980));
    defparam RAM_DATA_cl_6_RNO_0_15_LC_13_17_3.C_ON=1'b0;
    defparam RAM_DATA_cl_6_RNO_0_15_LC_13_17_3.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_6_RNO_0_15_LC_13_17_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 RAM_DATA_cl_6_RNO_0_15_LC_13_17_3 (
            .in0(_gnd_net_),
            .in1(N__32702),
            .in2(_gnd_net_),
            .in3(N__31696),
            .lcout(),
            .ltout(N_108_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_6_15_LC_13_17_4.C_ON=1'b0;
    defparam RAM_DATA_cl_6_15_LC_13_17_4.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_6_15_LC_13_17_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 RAM_DATA_cl_6_15_LC_13_17_4 (
            .in0(N__32494),
            .in1(N__32224),
            .in2(N__32724),
            .in3(N__31947),
            .lcout(RAM_DATA_cl_6Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47809),
            .ce(),
            .sr(N__52980));
    defparam RAM_DATA_cl_7_RNO_0_15_LC_13_17_5.C_ON=1'b0;
    defparam RAM_DATA_cl_7_RNO_0_15_LC_13_17_5.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_7_RNO_0_15_LC_13_17_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 RAM_DATA_cl_7_RNO_0_15_LC_13_17_5 (
            .in0(_gnd_net_),
            .in1(N__31757),
            .in2(_gnd_net_),
            .in3(N__31697),
            .lcout(),
            .ltout(N_95_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RAM_DATA_cl_7_15_LC_13_17_6.C_ON=1'b0;
    defparam RAM_DATA_cl_7_15_LC_13_17_6.SEQ_MODE=4'b1010;
    defparam RAM_DATA_cl_7_15_LC_13_17_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 RAM_DATA_cl_7_15_LC_13_17_6 (
            .in0(N__32495),
            .in1(N__32225),
            .in2(N__31980),
            .in3(N__31948),
            .lcout(RAM_DATA_cl_7Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47809),
            .ce(),
            .sr(N__52980));
    defparam RAM_DATA_cl_4_RNO_0_15_LC_13_17_7.C_ON=1'b0;
    defparam RAM_DATA_cl_4_RNO_0_15_LC_13_17_7.SEQ_MODE=4'b0000;
    defparam RAM_DATA_cl_4_RNO_0_15_LC_13_17_7.LUT_INIT=16'b0011001100000000;
    LogicCell40 RAM_DATA_cl_4_RNO_0_15_LC_13_17_7 (
            .in0(_gnd_net_),
            .in1(N__31724),
            .in2(_gnd_net_),
            .in3(N__31694),
            .lcout(N_105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sRAM_pointer_write_0_LC_13_18_0.C_ON=1'b1;
    defparam sRAM_pointer_write_0_LC_13_18_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_0_LC_13_18_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_0_LC_13_18_0 (
            .in0(N__33556),
            .in1(N__31619),
            .in2(_gnd_net_),
            .in3(N__31608),
            .lcout(sRAM_pointer_writeZ0Z_0),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(sRAM_pointer_write_cry_0),
            .clk(N__47818),
            .ce(N__33306),
            .sr(N__52976));
    defparam sRAM_pointer_write_1_LC_13_18_1.C_ON=1'b1;
    defparam sRAM_pointer_write_1_LC_13_18_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_1_LC_13_18_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_1_LC_13_18_1 (
            .in0(N__33552),
            .in1(N__31601),
            .in2(_gnd_net_),
            .in3(N__32928),
            .lcout(sRAM_pointer_writeZ0Z_1),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_0),
            .carryout(sRAM_pointer_write_cry_1),
            .clk(N__47818),
            .ce(N__33306),
            .sr(N__52976));
    defparam sRAM_pointer_write_2_LC_13_18_2.C_ON=1'b1;
    defparam sRAM_pointer_write_2_LC_13_18_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_2_LC_13_18_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_2_LC_13_18_2 (
            .in0(N__33557),
            .in1(N__32918),
            .in2(_gnd_net_),
            .in3(N__32907),
            .lcout(sRAM_pointer_writeZ0Z_2),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_1),
            .carryout(sRAM_pointer_write_cry_2),
            .clk(N__47818),
            .ce(N__33306),
            .sr(N__52976));
    defparam sRAM_pointer_write_3_LC_13_18_3.C_ON=1'b1;
    defparam sRAM_pointer_write_3_LC_13_18_3.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_3_LC_13_18_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_3_LC_13_18_3 (
            .in0(N__33553),
            .in1(N__32897),
            .in2(_gnd_net_),
            .in3(N__32886),
            .lcout(sRAM_pointer_writeZ0Z_3),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_2),
            .carryout(sRAM_pointer_write_cry_3),
            .clk(N__47818),
            .ce(N__33306),
            .sr(N__52976));
    defparam sRAM_pointer_write_4_LC_13_18_4.C_ON=1'b1;
    defparam sRAM_pointer_write_4_LC_13_18_4.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_4_LC_13_18_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_4_LC_13_18_4 (
            .in0(N__33558),
            .in1(N__32873),
            .in2(_gnd_net_),
            .in3(N__32862),
            .lcout(sRAM_pointer_writeZ0Z_4),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_3),
            .carryout(sRAM_pointer_write_cry_4),
            .clk(N__47818),
            .ce(N__33306),
            .sr(N__52976));
    defparam sRAM_pointer_write_5_LC_13_18_5.C_ON=1'b1;
    defparam sRAM_pointer_write_5_LC_13_18_5.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_5_LC_13_18_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_5_LC_13_18_5 (
            .in0(N__33554),
            .in1(N__32852),
            .in2(_gnd_net_),
            .in3(N__32841),
            .lcout(sRAM_pointer_writeZ0Z_5),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_4),
            .carryout(sRAM_pointer_write_cry_5),
            .clk(N__47818),
            .ce(N__33306),
            .sr(N__52976));
    defparam sRAM_pointer_write_6_LC_13_18_6.C_ON=1'b1;
    defparam sRAM_pointer_write_6_LC_13_18_6.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_6_LC_13_18_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_6_LC_13_18_6 (
            .in0(N__33559),
            .in1(N__32834),
            .in2(_gnd_net_),
            .in3(N__32823),
            .lcout(sRAM_pointer_writeZ0Z_6),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_5),
            .carryout(sRAM_pointer_write_cry_6),
            .clk(N__47818),
            .ce(N__33306),
            .sr(N__52976));
    defparam sRAM_pointer_write_7_LC_13_18_7.C_ON=1'b1;
    defparam sRAM_pointer_write_7_LC_13_18_7.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_7_LC_13_18_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_7_LC_13_18_7 (
            .in0(N__33555),
            .in1(N__32816),
            .in2(_gnd_net_),
            .in3(N__32805),
            .lcout(sRAM_pointer_writeZ0Z_7),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_6),
            .carryout(sRAM_pointer_write_cry_7),
            .clk(N__47818),
            .ce(N__33306),
            .sr(N__52976));
    defparam sRAM_pointer_write_8_LC_13_19_0.C_ON=1'b1;
    defparam sRAM_pointer_write_8_LC_13_19_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_8_LC_13_19_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_8_LC_13_19_0 (
            .in0(N__33567),
            .in1(N__32795),
            .in2(_gnd_net_),
            .in3(N__32784),
            .lcout(sRAM_pointer_writeZ0Z_8),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(sRAM_pointer_write_cry_8),
            .clk(N__47825),
            .ce(N__33305),
            .sr(N__52973));
    defparam sRAM_pointer_write_9_LC_13_19_1.C_ON=1'b1;
    defparam sRAM_pointer_write_9_LC_13_19_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_9_LC_13_19_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_9_LC_13_19_1 (
            .in0(N__33563),
            .in1(N__32771),
            .in2(_gnd_net_),
            .in3(N__32760),
            .lcout(sRAM_pointer_writeZ0Z_9),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_8),
            .carryout(sRAM_pointer_write_cry_9),
            .clk(N__47825),
            .ce(N__33305),
            .sr(N__52973));
    defparam sRAM_pointer_write_10_LC_13_19_2.C_ON=1'b1;
    defparam sRAM_pointer_write_10_LC_13_19_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_10_LC_13_19_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_10_LC_13_19_2 (
            .in0(N__33564),
            .in1(N__33092),
            .in2(_gnd_net_),
            .in3(N__33081),
            .lcout(sRAM_pointer_writeZ0Z_10),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_9),
            .carryout(sRAM_pointer_write_cry_10),
            .clk(N__47825),
            .ce(N__33305),
            .sr(N__52973));
    defparam sRAM_pointer_write_11_LC_13_19_3.C_ON=1'b1;
    defparam sRAM_pointer_write_11_LC_13_19_3.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_11_LC_13_19_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_11_LC_13_19_3 (
            .in0(N__33560),
            .in1(N__33071),
            .in2(_gnd_net_),
            .in3(N__33060),
            .lcout(sRAM_pointer_writeZ0Z_11),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_10),
            .carryout(sRAM_pointer_write_cry_11),
            .clk(N__47825),
            .ce(N__33305),
            .sr(N__52973));
    defparam sRAM_pointer_write_12_LC_13_19_4.C_ON=1'b1;
    defparam sRAM_pointer_write_12_LC_13_19_4.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_12_LC_13_19_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_12_LC_13_19_4 (
            .in0(N__33565),
            .in1(N__33050),
            .in2(_gnd_net_),
            .in3(N__33039),
            .lcout(sRAM_pointer_writeZ0Z_12),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_11),
            .carryout(sRAM_pointer_write_cry_12),
            .clk(N__47825),
            .ce(N__33305),
            .sr(N__52973));
    defparam sRAM_pointer_write_13_LC_13_19_5.C_ON=1'b1;
    defparam sRAM_pointer_write_13_LC_13_19_5.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_13_LC_13_19_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_13_LC_13_19_5 (
            .in0(N__33561),
            .in1(N__33029),
            .in2(_gnd_net_),
            .in3(N__33018),
            .lcout(sRAM_pointer_writeZ0Z_13),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_12),
            .carryout(sRAM_pointer_write_cry_13),
            .clk(N__47825),
            .ce(N__33305),
            .sr(N__52973));
    defparam sRAM_pointer_write_14_LC_13_19_6.C_ON=1'b1;
    defparam sRAM_pointer_write_14_LC_13_19_6.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_14_LC_13_19_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_14_LC_13_19_6 (
            .in0(N__33566),
            .in1(N__33008),
            .in2(_gnd_net_),
            .in3(N__32997),
            .lcout(sRAM_pointer_writeZ0Z_14),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_13),
            .carryout(sRAM_pointer_write_cry_14),
            .clk(N__47825),
            .ce(N__33305),
            .sr(N__52973));
    defparam sRAM_pointer_write_15_LC_13_19_7.C_ON=1'b1;
    defparam sRAM_pointer_write_15_LC_13_19_7.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_15_LC_13_19_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_15_LC_13_19_7 (
            .in0(N__33562),
            .in1(N__32987),
            .in2(_gnd_net_),
            .in3(N__32976),
            .lcout(sRAM_pointer_writeZ0Z_15),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_14),
            .carryout(sRAM_pointer_write_cry_15),
            .clk(N__47825),
            .ce(N__33305),
            .sr(N__52973));
    defparam sRAM_pointer_write_16_LC_13_20_0.C_ON=1'b1;
    defparam sRAM_pointer_write_16_LC_13_20_0.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_16_LC_13_20_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_16_LC_13_20_0 (
            .in0(N__33542),
            .in1(N__32969),
            .in2(_gnd_net_),
            .in3(N__32955),
            .lcout(sRAM_pointer_writeZ0Z_16),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(sRAM_pointer_write_cry_16),
            .clk(N__47835),
            .ce(N__33304),
            .sr(N__52969));
    defparam sRAM_pointer_write_17_LC_13_20_1.C_ON=1'b1;
    defparam sRAM_pointer_write_17_LC_13_20_1.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_17_LC_13_20_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_17_LC_13_20_1 (
            .in0(N__33541),
            .in1(N__32942),
            .in2(_gnd_net_),
            .in3(N__32931),
            .lcout(sRAM_pointer_writeZ0Z_17),
            .ltout(),
            .carryin(sRAM_pointer_write_cry_16),
            .carryout(sRAM_pointer_write_cry_17),
            .clk(N__47835),
            .ce(N__33304),
            .sr(N__52969));
    defparam sRAM_pointer_write_18_LC_13_20_2.C_ON=1'b0;
    defparam sRAM_pointer_write_18_LC_13_20_2.SEQ_MODE=4'b1010;
    defparam sRAM_pointer_write_18_LC_13_20_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 sRAM_pointer_write_18_LC_13_20_2 (
            .in0(N__33543),
            .in1(N__33320),
            .in2(_gnd_net_),
            .in3(N__33330),
            .lcout(sRAM_pointer_writeZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47835),
            .ce(N__33304),
            .sr(N__52969));
    defparam sDAC_mem_pointer_RNIF3GH_6_LC_14_1_3.C_ON=1'b0;
    defparam sDAC_mem_pointer_RNIF3GH_6_LC_14_1_3.SEQ_MODE=4'b0000;
    defparam sDAC_mem_pointer_RNIF3GH_6_LC_14_1_3.LUT_INIT=16'b0000000000110011;
    LogicCell40 sDAC_mem_pointer_RNIF3GH_6_LC_14_1_3 (
            .in0(_gnd_net_),
            .in1(N__37272),
            .in2(_gnd_net_),
            .in3(N__37278),
            .lcout(un17_sdacdyn_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1_1_LC_14_2_0 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1_1_LC_14_2_0 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1_1_LC_14_2_0 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1_1_LC_14_2_0  (
            .in0(N__33277),
            .in1(N__38553),
            .in2(N__37188),
            .in3(N__52415),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_i_RNI0OVC1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIOASC_5_LC_14_2_1 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIOASC_5_LC_14_2_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIOASC_5_LC_14_2_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNIOASC_5_LC_14_2_1  (
            .in0(N__37103),
            .in1(N__37118),
            .in2(N__37244),
            .in3(N__37343),
            .lcout(),
            .ltout(\spi_slave_inst.tx_data_count_neg_sclk_i6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI1DAJ_1_LC_14_2_2 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI1DAJ_1_LC_14_2_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNI1DAJ_1_LC_14_2_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNI1DAJ_1_LC_14_2_2  (
            .in0(N__37138),
            .in1(_gnd_net_),
            .in2(N__33234),
            .in3(N__37207),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_i6 ),
            .ltout(\spi_slave_inst.tx_data_count_neg_sclk_i6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_done_neg_sclk_i_LC_14_2_3 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_done_neg_sclk_i_LC_14_2_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_done_neg_sclk_i_LC_14_2_3 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \spi_slave_inst.tx_done_neg_sclk_i_LC_14_2_3  (
            .in0(_gnd_net_),
            .in1(N__33213),
            .in2(N__33162),
            .in3(N__33149),
            .lcout(\spi_slave_inst.tx_done_neg_sclk_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVspi_slave_inst.tx_done_neg_sclk_iC_net ),
            .ce(),
            .sr(N__53125));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIKKJ63_0_LC_14_2_5 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIKKJ63_0_LC_14_2_5 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIKKJ63_0_LC_14_2_5 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNIKKJ63_0_LC_14_2_5  (
            .in0(N__38554),
            .in1(N__38594),
            .in2(N__33138),
            .in3(N__52314),
            .lcout(spi_miso_rpi_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_13_3_LC_14_4_0.C_ON=1'b0;
    defparam sDAC_data_RNO_13_3_LC_14_4_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_3_LC_14_4_0.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_13_3_LC_14_4_0 (
            .in0(N__52156),
            .in1(N__41661),
            .in2(N__43666),
            .in3(N__33606),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_3_LC_14_4_1.C_ON=1'b0;
    defparam sDAC_data_RNO_5_3_LC_14_4_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_3_LC_14_4_1.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_5_3_LC_14_4_1 (
            .in0(N__52161),
            .in1(N__40068),
            .in2(N__33099),
            .in3(N__37296),
            .lcout(sDAC_data_RNO_5Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_6_0_LC_14_4_2.C_ON=1'b0;
    defparam sDAC_mem_6_0_LC_14_4_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_0_LC_14_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_0_LC_14_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50986),
            .lcout(sDAC_mem_6Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47810),
            .ce(N__43071),
            .sr(N__53098));
    defparam sDAC_data_RNO_13_4_LC_14_4_3.C_ON=1'b0;
    defparam sDAC_data_RNO_13_4_LC_14_4_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_4_LC_14_4_3.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_13_4_LC_14_4_3 (
            .in0(N__52160),
            .in1(N__33600),
            .in2(N__43668),
            .in3(N__33591),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_4_LC_14_4_4.C_ON=1'b0;
    defparam sDAC_data_RNO_5_4_LC_14_4_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_4_LC_14_4_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_5_4_LC_14_4_4 (
            .in0(N__52157),
            .in1(N__40059),
            .in2(N__33594),
            .in3(N__37290),
            .lcout(sDAC_data_RNO_5Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_6_1_LC_14_4_5.C_ON=1'b0;
    defparam sDAC_mem_6_1_LC_14_4_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_1_LC_14_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_1_LC_14_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50600),
            .lcout(sDAC_mem_6Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47810),
            .ce(N__43071),
            .sr(N__53098));
    defparam sDAC_data_RNO_13_5_LC_14_4_6.C_ON=1'b0;
    defparam sDAC_data_RNO_13_5_LC_14_4_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_5_LC_14_4_6.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_13_5_LC_14_4_6 (
            .in0(N__52158),
            .in1(N__41646),
            .in2(N__43667),
            .in3(N__33585),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_5_LC_14_4_7.C_ON=1'b0;
    defparam sDAC_data_RNO_5_5_LC_14_4_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_5_LC_14_4_7.LUT_INIT=16'b1100101100001011;
    LogicCell40 sDAC_data_RNO_5_5_LC_14_4_7 (
            .in0(N__40182),
            .in1(N__52159),
            .in2(N__33579),
            .in3(N__37368),
            .lcout(sDAC_data_RNO_5Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_12_5_LC_14_5_0.C_ON=1'b0;
    defparam sDAC_data_RNO_12_5_LC_14_5_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_5_LC_14_5_0.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_12_5_LC_14_5_0 (
            .in0(N__51910),
            .in1(N__38733),
            .in2(N__43673),
            .in3(N__33573),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_5_LC_14_5_1.C_ON=1'b0;
    defparam sDAC_data_RNO_4_5_LC_14_5_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_5_LC_14_5_1.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_5_LC_14_5_1 (
            .in0(N__52138),
            .in1(N__38769),
            .in2(N__33576),
            .in3(N__37359),
            .lcout(sDAC_data_RNO_4Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_4_2_LC_14_5_2.C_ON=1'b0;
    defparam sDAC_mem_4_2_LC_14_5_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_2_LC_14_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_2_LC_14_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50106),
            .lcout(sDAC_mem_4Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47799),
            .ce(N__39627),
            .sr(N__53085));
    defparam sDAC_data_RNO_12_6_LC_14_5_3.C_ON=1'b0;
    defparam sDAC_data_RNO_12_6_LC_14_5_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_6_LC_14_5_3.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_12_6_LC_14_5_3 (
            .in0(N__52137),
            .in1(N__38721),
            .in2(N__43671),
            .in3(N__33648),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_6_LC_14_5_4.C_ON=1'b0;
    defparam sDAC_data_RNO_4_6_LC_14_5_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_6_LC_14_5_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_6_LC_14_5_4 (
            .in0(N__51907),
            .in1(N__38760),
            .in2(N__33651),
            .in3(N__37353),
            .lcout(sDAC_data_RNO_4Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_4_3_LC_14_5_5.C_ON=1'b0;
    defparam sDAC_mem_4_3_LC_14_5_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_3_LC_14_5_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_4_3_LC_14_5_5 (
            .in0(N__49608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_4Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47799),
            .ce(N__39627),
            .sr(N__53085));
    defparam sDAC_data_RNO_12_7_LC_14_5_6.C_ON=1'b0;
    defparam sDAC_data_RNO_12_7_LC_14_5_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_7_LC_14_5_6.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_12_7_LC_14_5_6 (
            .in0(N__51908),
            .in1(N__38709),
            .in2(N__43672),
            .in3(N__33642),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_7_LC_14_5_7.C_ON=1'b0;
    defparam sDAC_data_RNO_4_7_LC_14_5_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_7_LC_14_5_7.LUT_INIT=16'b1010110000001111;
    LogicCell40 sDAC_data_RNO_4_7_LC_14_5_7 (
            .in0(N__37413),
            .in1(N__38751),
            .in2(N__33630),
            .in3(N__51909),
            .lcout(sDAC_data_RNO_4Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_3_0_LC_14_6_0.C_ON=1'b0;
    defparam sDAC_mem_3_0_LC_14_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_0_LC_14_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_3_0_LC_14_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51040),
            .lcout(sDAC_mem_3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47784),
            .ce(N__42960),
            .sr(N__53073));
    defparam sDAC_data_RNO_28_3_LC_14_6_1.C_ON=1'b0;
    defparam sDAC_data_RNO_28_3_LC_14_6_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_3_LC_14_6_1.LUT_INIT=16'b0100010101100111;
    LogicCell40 sDAC_data_RNO_28_3_LC_14_6_1 (
            .in0(N__43606),
            .in1(N__51902),
            .in2(N__33627),
            .in3(N__37332),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_3_LC_14_6_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_3_LC_14_6_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_3_LC_14_6_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_3_LC_14_6_2 (
            .in0(N__51903),
            .in1(N__40230),
            .in2(N__33618),
            .in3(N__33615),
            .lcout(sDAC_data_RNO_15Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_5_LC_14_6_3.C_ON=1'b0;
    defparam sDAC_data_RNO_17_5_LC_14_6_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_5_LC_14_6_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_5_LC_14_6_3 (
            .in0(N__43607),
            .in1(N__44184),
            .in2(_gnd_net_),
            .in3(N__44319),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_5_LC_14_6_4.C_ON=1'b0;
    defparam sDAC_data_RNO_8_5_LC_14_6_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_5_LC_14_6_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 sDAC_data_RNO_8_5_LC_14_6_4 (
            .in0(N__51904),
            .in1(_gnd_net_),
            .in2(N__33609),
            .in3(N__45207),
            .lcout(sDAC_data_RNO_8Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_5_LC_14_6_5.C_ON=1'b0;
    defparam sDAC_data_RNO_16_5_LC_14_6_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_5_LC_14_6_5.LUT_INIT=16'b0000110100111101;
    LogicCell40 sDAC_data_RNO_16_5_LC_14_6_5 (
            .in0(N__38742),
            .in1(N__51905),
            .in2(N__43665),
            .in3(N__41832),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_5_LC_14_6_6.C_ON=1'b0;
    defparam sDAC_data_RNO_7_5_LC_14_6_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_5_LC_14_6_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_7_5_LC_14_6_6 (
            .in0(N__51906),
            .in1(N__43974),
            .in2(N__33717),
            .in3(N__47193),
            .lcout(),
            .ltout(sDAC_data_RNO_7Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_5_LC_14_6_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_5_LC_14_6_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_5_LC_14_6_7.LUT_INIT=16'b0111001101100010;
    LogicCell40 sDAC_data_RNO_2_5_LC_14_6_7 (
            .in0(N__45874),
            .in1(N__34065),
            .in2(N__33714),
            .in3(N__33711),
            .lcout(sDAC_data_RNO_2Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_5_LC_14_7_0.C_ON=1'b0;
    defparam sDAC_data_RNO_10_5_LC_14_7_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_5_LC_14_7_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_10_5_LC_14_7_0 (
            .in0(N__33705),
            .in1(N__41919),
            .in2(N__45908),
            .in3(N__33693),
            .lcout(),
            .ltout(sDAC_data_RNO_10Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_5_LC_14_7_1.C_ON=1'b0;
    defparam sDAC_data_RNO_3_5_LC_14_7_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_5_LC_14_7_1.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_3_5_LC_14_7_1 (
            .in0(N__42528),
            .in1(N__42638),
            .in2(N__33696),
            .in3(N__38412),
            .lcout(sDAC_data_2_41_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_5_LC_14_7_2.C_ON=1'b0;
    defparam sDAC_data_RNO_22_5_LC_14_7_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_5_LC_14_7_2.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_22_5_LC_14_7_2 (
            .in0(N__45861),
            .in1(N__45518),
            .in2(N__36681),
            .in3(N__34104),
            .lcout(sDAC_data_2_32_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_5_LC_14_7_3.C_ON=1'b0;
    defparam sDAC_data_RNO_6_5_LC_14_7_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_5_LC_14_7_3.LUT_INIT=16'b0100010101100111;
    LogicCell40 sDAC_data_RNO_6_5_LC_14_7_3 (
            .in0(N__45519),
            .in1(N__45865),
            .in2(N__33918),
            .in3(N__33738),
            .lcout(),
            .ltout(sDAC_data_2_14_ns_1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_5_LC_14_7_4.C_ON=1'b0;
    defparam sDAC_data_RNO_1_5_LC_14_7_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_5_LC_14_7_4.LUT_INIT=16'b1100101100001011;
    LogicCell40 sDAC_data_RNO_1_5_LC_14_7_4 (
            .in0(N__33687),
            .in1(N__45866),
            .in2(N__33678),
            .in3(N__33675),
            .lcout(),
            .ltout(sDAC_data_RNO_1Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_5_LC_14_7_5.C_ON=1'b0;
    defparam sDAC_data_RNO_0_5_LC_14_7_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_5_LC_14_7_5.LUT_INIT=16'b0101000011101110;
    LogicCell40 sDAC_data_RNO_0_5_LC_14_7_5 (
            .in0(N__42529),
            .in1(N__33666),
            .in2(N__33660),
            .in3(N__33657),
            .lcout(),
            .ltout(sDAC_data_2_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_5_LC_14_7_6.C_ON=1'b0;
    defparam sDAC_data_5_LC_14_7_6.SEQ_MODE=4'b1010;
    defparam sDAC_data_5_LC_14_7_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 sDAC_data_5_LC_14_7_6 (
            .in0(_gnd_net_),
            .in1(N__45990),
            .in2(N__33771),
            .in3(N__42381),
            .lcout(sDAC_dataZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53248),
            .ce(N__42230),
            .sr(N__53061));
    defparam sDAC_mem_3_2_LC_14_8_0.C_ON=1'b0;
    defparam sDAC_mem_3_2_LC_14_8_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_2_LC_14_8_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_3_2_LC_14_8_0 (
            .in0(N__50187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_3Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47758),
            .ce(N__42977),
            .sr(N__53051));
    defparam sDAC_data_RNO_28_5_LC_14_8_1.C_ON=1'b0;
    defparam sDAC_data_RNO_28_5_LC_14_8_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_5_LC_14_8_1.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_28_5_LC_14_8_1 (
            .in0(N__51815),
            .in1(N__37320),
            .in2(N__43621),
            .in3(N__33756),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_5_LC_14_8_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_5_LC_14_8_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_5_LC_14_8_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_5_LC_14_8_2 (
            .in0(N__51818),
            .in1(N__40221),
            .in2(N__33747),
            .in3(N__33744),
            .lcout(sDAC_data_RNO_15Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_7_LC_14_8_3.C_ON=1'b0;
    defparam sDAC_data_RNO_16_7_LC_14_8_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_7_LC_14_8_3.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_16_7_LC_14_8_3 (
            .in0(N__51814),
            .in1(N__41808),
            .in2(N__43620),
            .in3(N__38829),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_7_LC_14_8_4.C_ON=1'b0;
    defparam sDAC_data_RNO_7_7_LC_14_8_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_7_LC_14_8_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_7_7_LC_14_8_4 (
            .in0(N__51817),
            .in1(N__44259),
            .in2(N__33732),
            .in3(N__47166),
            .lcout(sDAC_data_RNO_7Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_7_LC_14_8_5.C_ON=1'b0;
    defparam sDAC_data_RNO_17_7_LC_14_8_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_7_LC_14_8_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_7_LC_14_8_5 (
            .in0(N__43542),
            .in1(N__44157),
            .in2(_gnd_net_),
            .in3(N__44292),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_7_LC_14_8_6.C_ON=1'b0;
    defparam sDAC_data_RNO_8_7_LC_14_8_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_7_LC_14_8_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_8_7_LC_14_8_6 (
            .in0(_gnd_net_),
            .in1(N__51816),
            .in2(N__33729),
            .in3(N__45180),
            .lcout(),
            .ltout(sDAC_data_RNO_8Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_7_LC_14_8_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_7_LC_14_8_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_7_LC_14_8_7.LUT_INIT=16'b0111011000110010;
    LogicCell40 sDAC_data_RNO_2_7_LC_14_8_7 (
            .in0(N__45783),
            .in1(N__43914),
            .in2(N__33726),
            .in3(N__33723),
            .lcout(sDAC_data_RNO_2Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_27_8_LC_14_9_0.C_ON=1'b0;
    defparam sDAC_data_RNO_27_8_LC_14_9_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_8_LC_14_9_0.LUT_INIT=16'b1111101111001000;
    LogicCell40 sDAC_data_RNO_27_8_LC_14_9_0 (
            .in0(N__43520),
            .in1(N__51555),
            .in2(N__33834),
            .in3(N__33849),
            .lcout(),
            .ltout(sDAC_data_RNO_27Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_8_LC_14_9_1.C_ON=1'b0;
    defparam sDAC_data_RNO_14_8_LC_14_9_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_8_LC_14_9_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 sDAC_data_RNO_14_8_LC_14_9_1 (
            .in0(N__33864),
            .in1(_gnd_net_),
            .in2(N__33852),
            .in3(N__33840),
            .lcout(sDAC_data_RNO_14Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_26_8_LC_14_9_2.C_ON=1'b0;
    defparam sDAC_data_RNO_26_8_LC_14_9_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_8_LC_14_9_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 sDAC_data_RNO_26_8_LC_14_9_2 (
            .in0(N__43518),
            .in1(N__51553),
            .in2(N__33833),
            .in3(N__33848),
            .lcout(sDAC_data_RNO_26Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_1_5_LC_14_9_3.C_ON=1'b0;
    defparam sDAC_mem_1_5_LC_14_9_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_5_LC_14_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_5_LC_14_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47016),
            .lcout(sDAC_mem_1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47744),
            .ce(N__42032),
            .sr(N__53041));
    defparam sDAC_data_RNO_26_9_LC_14_9_4.C_ON=1'b0;
    defparam sDAC_data_RNO_26_9_LC_14_9_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_9_LC_14_9_4.LUT_INIT=16'b0111010000110000;
    LogicCell40 sDAC_data_RNO_26_9_LC_14_9_4 (
            .in0(N__43519),
            .in1(N__51554),
            .in2(N__33804),
            .in3(N__33780),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_9_LC_14_9_5.C_ON=1'b0;
    defparam sDAC_data_RNO_14_9_LC_14_9_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_9_LC_14_9_5.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_14_9_LC_14_9_5 (
            .in0(_gnd_net_),
            .in1(N__33819),
            .in2(N__33807),
            .in3(N__33786),
            .lcout(sDAC_data_RNO_14Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_27_9_LC_14_9_6.C_ON=1'b0;
    defparam sDAC_data_RNO_27_9_LC_14_9_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_9_LC_14_9_6.LUT_INIT=16'b1111110010111000;
    LogicCell40 sDAC_data_RNO_27_9_LC_14_9_6 (
            .in0(N__43517),
            .in1(N__51552),
            .in2(N__33803),
            .in3(N__33779),
            .lcout(sDAC_data_RNO_27Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_1_6_LC_14_9_7.C_ON=1'b0;
    defparam sDAC_mem_1_6_LC_14_9_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_6_LC_14_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_6_LC_14_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48233),
            .lcout(sDAC_mem_1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47744),
            .ce(N__42032),
            .sr(N__53041));
    defparam sDAC_mem_3_6_LC_14_10_0.C_ON=1'b0;
    defparam sDAC_mem_3_6_LC_14_10_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_6_LC_14_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_3_6_LC_14_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48255),
            .lcout(sDAC_mem_3Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47733),
            .ce(N__42978),
            .sr(N__53032));
    defparam sDAC_data_RNO_28_9_LC_14_10_1.C_ON=1'b0;
    defparam sDAC_data_RNO_28_9_LC_14_10_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_9_LC_14_10_1.LUT_INIT=16'b0100010101100111;
    LogicCell40 sDAC_data_RNO_28_9_LC_14_10_1 (
            .in0(N__43514),
            .in1(N__51599),
            .in2(N__34008),
            .in3(N__37308),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_9_LC_14_10_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_9_LC_14_10_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_9_LC_14_10_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_9_LC_14_10_2 (
            .in0(N__51601),
            .in1(N__40722),
            .in2(N__33993),
            .in3(N__33990),
            .lcout(sDAC_data_RNO_15Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_26_4_LC_14_10_3.C_ON=1'b0;
    defparam sDAC_data_RNO_26_4_LC_14_10_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_4_LC_14_10_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 sDAC_data_RNO_26_4_LC_14_10_3 (
            .in0(N__43515),
            .in1(N__51600),
            .in2(N__33969),
            .in3(N__33947),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_4_LC_14_10_4.C_ON=1'b0;
    defparam sDAC_data_RNO_14_4_LC_14_10_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_4_LC_14_10_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_14_4_LC_14_10_4 (
            .in0(_gnd_net_),
            .in1(N__33984),
            .in2(N__33972),
            .in3(N__33939),
            .lcout(sDAC_data_RNO_14Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_27_4_LC_14_10_5.C_ON=1'b0;
    defparam sDAC_data_RNO_27_4_LC_14_10_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_4_LC_14_10_5.LUT_INIT=16'b1111101111001000;
    LogicCell40 sDAC_data_RNO_27_4_LC_14_10_5 (
            .in0(N__43513),
            .in1(N__51598),
            .in2(N__33968),
            .in3(N__33948),
            .lcout(sDAC_data_RNO_27Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_26_5_LC_14_10_6.C_ON=1'b0;
    defparam sDAC_data_RNO_26_5_LC_14_10_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_5_LC_14_10_6.LUT_INIT=16'b0111001001010000;
    LogicCell40 sDAC_data_RNO_26_5_LC_14_10_6 (
            .in0(N__51602),
            .in1(N__43516),
            .in2(N__33906),
            .in3(N__33891),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_5_LC_14_10_7.C_ON=1'b0;
    defparam sDAC_data_RNO_14_5_LC_14_10_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_5_LC_14_10_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 sDAC_data_RNO_14_5_LC_14_10_7 (
            .in0(N__33933),
            .in1(_gnd_net_),
            .in2(N__33921),
            .in3(N__33873),
            .lcout(sDAC_data_RNO_14Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_27_3_LC_14_11_0.C_ON=1'b0;
    defparam sDAC_data_RNO_27_3_LC_14_11_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_3_LC_14_11_0.LUT_INIT=16'b1111101111001000;
    LogicCell40 sDAC_data_RNO_27_3_LC_14_11_0 (
            .in0(N__43501),
            .in1(N__52083),
            .in2(N__39296),
            .in3(N__39263),
            .lcout(sDAC_data_RNO_27Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_27_5_LC_14_11_1.C_ON=1'b0;
    defparam sDAC_data_RNO_27_5_LC_14_11_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_5_LC_14_11_1.LUT_INIT=16'b1110111011100100;
    LogicCell40 sDAC_data_RNO_27_5_LC_14_11_1 (
            .in0(N__52082),
            .in1(N__33902),
            .in2(N__43550),
            .in3(N__33890),
            .lcout(sDAC_data_RNO_27Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_10_LC_14_11_2.C_ON=1'b0;
    defparam sDAC_data_RNO_17_10_LC_14_11_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_10_LC_14_11_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_10_LC_14_11_2 (
            .in0(N__43502),
            .in1(N__44355),
            .in2(_gnd_net_),
            .in3(N__34038),
            .lcout(sDAC_data_RNO_17Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_pointer_RNIAIV21_3_LC_14_11_3.C_ON=1'b0;
    defparam sDAC_mem_pointer_RNIAIV21_3_LC_14_11_3.SEQ_MODE=4'b0000;
    defparam sDAC_mem_pointer_RNIAIV21_3_LC_14_11_3.LUT_INIT=16'b1110000011000000;
    LogicCell40 sDAC_mem_pointer_RNIAIV21_3_LC_14_11_3 (
            .in0(N__52081),
            .in1(N__45639),
            .in2(N__42614),
            .in3(N__45372),
            .lcout(),
            .ltout(op_le_op_le_un15_sdacdynlt4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_pointer_RNI4LV52_4_LC_14_11_4.C_ON=1'b0;
    defparam sDAC_mem_pointer_RNI4LV52_4_LC_14_11_4.SEQ_MODE=4'b0000;
    defparam sDAC_mem_pointer_RNI4LV52_4_LC_14_11_4.LUT_INIT=16'b0101011100000000;
    LogicCell40 sDAC_mem_pointer_RNI4LV52_4_LC_14_11_4 (
            .in0(N__43500),
            .in1(N__42447),
            .in2(N__34050),
            .in3(N__34047),
            .lcout(un17_sdacdyn_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_10_7_LC_14_11_5.C_ON=1'b0;
    defparam sDAC_mem_10_7_LC_14_11_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_7_LC_14_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_7_LC_14_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48777),
            .lcout(sDAC_mem_10Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47724),
            .ce(N__45000),
            .sr(N__53022));
    defparam sDAC_data_RNO_9_10_LC_14_11_7.C_ON=1'b0;
    defparam sDAC_data_RNO_9_10_LC_14_11_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_10_LC_14_11_7.LUT_INIT=16'b0011000001011111;
    LogicCell40 sDAC_data_RNO_9_10_LC_14_11_7 (
            .in0(N__47274),
            .in1(N__51288),
            .in2(N__45807),
            .in3(N__45373),
            .lcout(sDAC_data_2_24_ns_1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_30_10_LC_14_12_0.C_ON=1'b0;
    defparam sDAC_data_RNO_30_10_LC_14_12_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_10_LC_14_12_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_30_10_LC_14_12_0 (
            .in0(N__34026),
            .in1(N__51597),
            .in2(_gnd_net_),
            .in3(N__34032),
            .lcout(sDAC_data_RNO_30Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_18_7_LC_14_12_1.C_ON=1'b0;
    defparam sDAC_mem_18_7_LC_14_12_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_7_LC_14_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_7_LC_14_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48816),
            .lcout(sDAC_mem_18Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47734),
            .ce(N__34088),
            .sr(N__53017));
    defparam sDAC_data_RNO_30_3_LC_14_12_2.C_ON=1'b0;
    defparam sDAC_data_RNO_30_3_LC_14_12_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_3_LC_14_12_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_30_3_LC_14_12_2 (
            .in0(N__34014),
            .in1(N__51596),
            .in2(_gnd_net_),
            .in3(N__34020),
            .lcout(sDAC_data_RNO_30Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_18_0_LC_14_12_3.C_ON=1'b0;
    defparam sDAC_mem_18_0_LC_14_12_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_0_LC_14_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_0_LC_14_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51246),
            .lcout(sDAC_mem_18Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47734),
            .ce(N__34088),
            .sr(N__53017));
    defparam sDAC_data_RNO_30_4_LC_14_12_4.C_ON=1'b0;
    defparam sDAC_data_RNO_30_4_LC_14_12_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_4_LC_14_12_4.LUT_INIT=16'b1111001111000000;
    LogicCell40 sDAC_data_RNO_30_4_LC_14_12_4 (
            .in0(_gnd_net_),
            .in1(N__51594),
            .in2(N__34125),
            .in3(N__34116),
            .lcout(sDAC_data_RNO_30Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_18_1_LC_14_12_5.C_ON=1'b0;
    defparam sDAC_mem_18_1_LC_14_12_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_1_LC_14_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_1_LC_14_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50575),
            .lcout(sDAC_mem_18Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47734),
            .ce(N__34088),
            .sr(N__53017));
    defparam sDAC_data_RNO_30_5_LC_14_12_6.C_ON=1'b0;
    defparam sDAC_data_RNO_30_5_LC_14_12_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_5_LC_14_12_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_30_5_LC_14_12_6 (
            .in0(N__34095),
            .in1(N__51595),
            .in2(_gnd_net_),
            .in3(N__34110),
            .lcout(sDAC_data_RNO_30Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_18_2_LC_14_12_7.C_ON=1'b0;
    defparam sDAC_mem_18_2_LC_14_12_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_18_2_LC_14_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_18_2_LC_14_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50261),
            .lcout(sDAC_mem_18Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47734),
            .ce(N__34088),
            .sr(N__53017));
    defparam sDAC_data_RNO_19_5_LC_14_13_0.C_ON=1'b0;
    defparam sDAC_data_RNO_19_5_LC_14_13_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_5_LC_14_13_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_19_5_LC_14_13_0 (
            .in0(N__43740),
            .in1(N__51865),
            .in2(_gnd_net_),
            .in3(N__45090),
            .lcout(sDAC_data_RNO_19Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_5_LC_14_13_1.C_ON=1'b0;
    defparam sDAC_data_RNO_18_5_LC_14_13_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_5_LC_14_13_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_5_LC_14_13_1 (
            .in0(N__51866),
            .in1(N__49857),
            .in2(_gnd_net_),
            .in3(N__34137),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_5_LC_14_13_2.C_ON=1'b0;
    defparam sDAC_data_RNO_9_5_LC_14_13_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_5_LC_14_13_2.LUT_INIT=16'b0001010110011101;
    LogicCell40 sDAC_data_RNO_9_5_LC_14_13_2 (
            .in0(N__45421),
            .in1(N__45859),
            .in2(N__34074),
            .in3(N__34071),
            .lcout(sDAC_data_2_24_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_6_LC_14_13_3.C_ON=1'b0;
    defparam sDAC_data_RNO_18_6_LC_14_13_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_6_LC_14_13_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_6_LC_14_13_3 (
            .in0(N__51867),
            .in1(N__49383),
            .in2(_gnd_net_),
            .in3(N__34131),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_6_LC_14_13_4.C_ON=1'b0;
    defparam sDAC_data_RNO_9_6_LC_14_13_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_6_LC_14_13_4.LUT_INIT=16'b0001010110011101;
    LogicCell40 sDAC_data_RNO_9_6_LC_14_13_4 (
            .in0(N__45422),
            .in1(N__45860),
            .in2(N__34053),
            .in3(N__34143),
            .lcout(sDAC_data_2_24_ns_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_19_6_LC_14_13_5.C_ON=1'b0;
    defparam sDAC_data_RNO_19_6_LC_14_13_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_6_LC_14_13_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_6_LC_14_13_5 (
            .in0(N__51864),
            .in1(N__45075),
            .in2(_gnd_net_),
            .in3(N__43728),
            .lcout(sDAC_data_RNO_19Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_12_2_LC_14_13_6.C_ON=1'b0;
    defparam sDAC_mem_12_2_LC_14_13_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_2_LC_14_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_2_LC_14_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50105),
            .lcout(sDAC_mem_12Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47745),
            .ce(N__47384),
            .sr(N__53011));
    defparam sDAC_mem_12_3_LC_14_13_7.C_ON=1'b0;
    defparam sDAC_mem_12_3_LC_14_13_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_3_LC_14_13_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_12_3_LC_14_13_7 (
            .in0(N__49795),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_12Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47745),
            .ce(N__47384),
            .sr(N__53011));
    defparam sDAC_mem_31_0_LC_14_14_0.C_ON=1'b0;
    defparam sDAC_mem_31_0_LC_14_14_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_0_LC_14_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_0_LC_14_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51261),
            .lcout(sDAC_mem_31Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47759),
            .ce(N__34380),
            .sr(N__53003));
    defparam sDAC_mem_31_1_LC_14_14_1.C_ON=1'b0;
    defparam sDAC_mem_31_1_LC_14_14_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_1_LC_14_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_1_LC_14_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50733),
            .lcout(sDAC_mem_31Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47759),
            .ce(N__34380),
            .sr(N__53003));
    defparam sDAC_mem_31_2_LC_14_14_2.C_ON=1'b0;
    defparam sDAC_mem_31_2_LC_14_14_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_2_LC_14_14_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_31_2_LC_14_14_2 (
            .in0(N__50262),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_31Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47759),
            .ce(N__34380),
            .sr(N__53003));
    defparam sDAC_mem_31_3_LC_14_14_3.C_ON=1'b0;
    defparam sDAC_mem_31_3_LC_14_14_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_3_LC_14_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_3_LC_14_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49796),
            .lcout(sDAC_mem_31Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47759),
            .ce(N__34380),
            .sr(N__53003));
    defparam sDAC_mem_31_4_LC_14_14_4.C_ON=1'b0;
    defparam sDAC_mem_31_4_LC_14_14_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_4_LC_14_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_4_LC_14_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49222),
            .lcout(sDAC_mem_31Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47759),
            .ce(N__34380),
            .sr(N__53003));
    defparam sDAC_mem_31_5_LC_14_14_5.C_ON=1'b0;
    defparam sDAC_mem_31_5_LC_14_14_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_5_LC_14_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_5_LC_14_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47073),
            .lcout(sDAC_mem_31Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47759),
            .ce(N__34380),
            .sr(N__53003));
    defparam sDAC_mem_31_6_LC_14_14_6.C_ON=1'b0;
    defparam sDAC_mem_31_6_LC_14_14_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_6_LC_14_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_6_LC_14_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48324),
            .lcout(sDAC_mem_31Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47759),
            .ce(N__34380),
            .sr(N__53003));
    defparam sDAC_mem_31_7_LC_14_14_7.C_ON=1'b0;
    defparam sDAC_mem_31_7_LC_14_14_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_31_7_LC_14_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_31_7_LC_14_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48842),
            .lcout(sDAC_mem_31Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47759),
            .ce(N__34380),
            .sr(N__53003));
    defparam sEEADC_freq_RNI4KIA1_2_LC_14_15_0.C_ON=1'b0;
    defparam sEEADC_freq_RNI4KIA1_2_LC_14_15_0.SEQ_MODE=4'b0000;
    defparam sEEADC_freq_RNI4KIA1_2_LC_14_15_0.LUT_INIT=16'b1000001001000001;
    LogicCell40 sEEADC_freq_RNI4KIA1_2_LC_14_15_0 (
            .in0(N__34335),
            .in1(N__34365),
            .in2(N__34329),
            .in3(N__34349),
            .lcout(un11_sacqtime_NE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEADC_freq_2_LC_14_15_1.C_ON=1'b0;
    defparam sEEADC_freq_2_LC_14_15_1.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_2_LC_14_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEADC_freq_2_LC_14_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50264),
            .lcout(sEEADC_freqZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47769),
            .ce(N__44127),
            .sr(_gnd_net_));
    defparam sEEADC_freq_3_LC_14_15_2.C_ON=1'b0;
    defparam sEEADC_freq_3_LC_14_15_2.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_3_LC_14_15_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEADC_freq_3_LC_14_15_2 (
            .in0(N__49798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEADC_freqZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47769),
            .ce(N__44127),
            .sr(_gnd_net_));
    defparam sEEADC_freq_RNICSIA1_4_LC_14_15_3.C_ON=1'b0;
    defparam sEEADC_freq_RNICSIA1_4_LC_14_15_3.SEQ_MODE=4'b0000;
    defparam sEEADC_freq_RNICSIA1_4_LC_14_15_3.LUT_INIT=16'b1000001001000001;
    LogicCell40 sEEADC_freq_RNICSIA1_4_LC_14_15_3 (
            .in0(N__34290),
            .in1(N__34319),
            .in2(N__34284),
            .in3(N__34305),
            .lcout(un11_sacqtime_NE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEADC_freq_4_LC_14_15_4.C_ON=1'b0;
    defparam sEEADC_freq_4_LC_14_15_4.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_4_LC_14_15_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEADC_freq_4_LC_14_15_4 (
            .in0(N__49165),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEADC_freqZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47769),
            .ce(N__44127),
            .sr(_gnd_net_));
    defparam sEEADC_freq_5_LC_14_15_5.C_ON=1'b0;
    defparam sEEADC_freq_5_LC_14_15_5.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_5_LC_14_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEADC_freq_5_LC_14_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47126),
            .lcout(sEEADC_freqZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47769),
            .ce(N__44127),
            .sr(_gnd_net_));
    defparam sEEADC_freq_RNIK4JA1_6_LC_14_15_6.C_ON=1'b0;
    defparam sEEADC_freq_RNIK4JA1_6_LC_14_15_6.SEQ_MODE=4'b0000;
    defparam sEEADC_freq_RNIK4JA1_6_LC_14_15_6.LUT_INIT=16'b1001000000001001;
    LogicCell40 sEEADC_freq_RNIK4JA1_6_LC_14_15_6 (
            .in0(N__34275),
            .in1(N__41451),
            .in2(N__41442),
            .in3(N__34260),
            .lcout(un11_sacqtime_NE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_0_c_inv_LC_14_16_0.C_ON=1'b1;
    defparam un5_sdacdyn_cry_0_c_inv_LC_14_16_0.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_0_c_inv_LC_14_16_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_0_c_inv_LC_14_16_0 (
            .in0(_gnd_net_),
            .in1(N__35088),
            .in2(N__34244),
            .in3(N__34161),
            .lcout(sEEACQ_i_0),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(un5_sdacdyn_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_1_c_inv_LC_14_16_1.C_ON=1'b1;
    defparam un5_sdacdyn_cry_1_c_inv_LC_14_16_1.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_1_c_inv_LC_14_16_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_sdacdyn_cry_1_c_inv_LC_14_16_1 (
            .in0(N__35082),
            .in1(N__35062),
            .in2(N__34977),
            .in3(_gnd_net_),
            .lcout(sEEACQ_i_1),
            .ltout(),
            .carryin(un5_sdacdyn_cry_0),
            .carryout(un5_sdacdyn_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_2_c_inv_LC_14_16_2.C_ON=1'b1;
    defparam un5_sdacdyn_cry_2_c_inv_LC_14_16_2.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_2_c_inv_LC_14_16_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_2_c_inv_LC_14_16_2 (
            .in0(_gnd_net_),
            .in1(N__34956),
            .in2(N__34866),
            .in3(N__34884),
            .lcout(sEEACQ_i_2),
            .ltout(),
            .carryin(un5_sdacdyn_cry_1),
            .carryout(un5_sdacdyn_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_3_c_inv_LC_14_16_3.C_ON=1'b1;
    defparam un5_sdacdyn_cry_3_c_inv_LC_14_16_3.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_3_c_inv_LC_14_16_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_3_c_inv_LC_14_16_3 (
            .in0(_gnd_net_),
            .in1(N__34856),
            .in2(N__34761),
            .in3(N__34779),
            .lcout(sEEACQ_i_3),
            .ltout(),
            .carryin(un5_sdacdyn_cry_2),
            .carryout(un5_sdacdyn_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_4_c_inv_LC_14_16_4.C_ON=1'b1;
    defparam un5_sdacdyn_cry_4_c_inv_LC_14_16_4.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_4_c_inv_LC_14_16_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_sdacdyn_cry_4_c_inv_LC_14_16_4 (
            .in0(N__34752),
            .in1(N__34734),
            .in2(N__36884),
            .in3(_gnd_net_),
            .lcout(sEEACQ_i_4),
            .ltout(),
            .carryin(un5_sdacdyn_cry_3),
            .carryout(un5_sdacdyn_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_5_c_inv_LC_14_16_5.C_ON=1'b1;
    defparam un5_sdacdyn_cry_5_c_inv_LC_14_16_5.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_5_c_inv_LC_14_16_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_5_c_inv_LC_14_16_5 (
            .in0(_gnd_net_),
            .in1(N__34726),
            .in2(N__34629),
            .in3(N__34647),
            .lcout(sEEACQ_i_5),
            .ltout(),
            .carryin(un5_sdacdyn_cry_4),
            .carryout(un5_sdacdyn_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_6_c_inv_LC_14_16_6.C_ON=1'b1;
    defparam un5_sdacdyn_cry_6_c_inv_LC_14_16_6.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_6_c_inv_LC_14_16_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_6_c_inv_LC_14_16_6 (
            .in0(_gnd_net_),
            .in1(N__34612),
            .in2(N__34503),
            .in3(N__34521),
            .lcout(sEEACQ_i_6),
            .ltout(),
            .carryin(un5_sdacdyn_cry_5),
            .carryout(un5_sdacdyn_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_7_c_inv_LC_14_16_7.C_ON=1'b1;
    defparam un5_sdacdyn_cry_7_c_inv_LC_14_16_7.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_7_c_inv_LC_14_16_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_7_c_inv_LC_14_16_7 (
            .in0(_gnd_net_),
            .in1(N__34386),
            .in2(N__34493),
            .in3(N__34404),
            .lcout(sEEACQ_i_7),
            .ltout(),
            .carryin(un5_sdacdyn_cry_6),
            .carryout(un5_sdacdyn_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_8_c_inv_LC_14_17_0.C_ON=1'b1;
    defparam un5_sdacdyn_cry_8_c_inv_LC_14_17_0.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_8_c_inv_LC_14_17_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_8_c_inv_LC_14_17_0 (
            .in0(_gnd_net_),
            .in1(N__35775),
            .in2(N__35888),
            .in3(N__35793),
            .lcout(sEEACQ_i_8),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(un5_sdacdyn_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_9_c_inv_LC_14_17_1.C_ON=1'b1;
    defparam un5_sdacdyn_cry_9_c_inv_LC_14_17_1.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_9_c_inv_LC_14_17_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_9_c_inv_LC_14_17_1 (
            .in0(_gnd_net_),
            .in1(N__35769),
            .in2(N__35664),
            .in3(N__35682),
            .lcout(sEEACQ_i_9),
            .ltout(),
            .carryin(un5_sdacdyn_cry_8),
            .carryout(un5_sdacdyn_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_10_c_inv_LC_14_17_2.C_ON=1'b1;
    defparam un5_sdacdyn_cry_10_c_inv_LC_14_17_2.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_10_c_inv_LC_14_17_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_10_c_inv_LC_14_17_2 (
            .in0(_gnd_net_),
            .in1(N__35646),
            .in2(N__35550),
            .in3(N__35571),
            .lcout(sEEACQ_i_10),
            .ltout(),
            .carryin(un5_sdacdyn_cry_9),
            .carryout(un5_sdacdyn_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_11_c_inv_LC_14_17_3.C_ON=1'b1;
    defparam un5_sdacdyn_cry_11_c_inv_LC_14_17_3.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_11_c_inv_LC_14_17_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_11_c_inv_LC_14_17_3 (
            .in0(_gnd_net_),
            .in1(N__35540),
            .in2(N__35445),
            .in3(N__35463),
            .lcout(sEEACQ_i_11),
            .ltout(),
            .carryin(un5_sdacdyn_cry_10),
            .carryout(un5_sdacdyn_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_12_c_inv_LC_14_17_4.C_ON=1'b1;
    defparam un5_sdacdyn_cry_12_c_inv_LC_14_17_4.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_12_c_inv_LC_14_17_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_sdacdyn_cry_12_c_inv_LC_14_17_4 (
            .in0(N__35436),
            .in1(N__35409),
            .in2(N__35328),
            .in3(_gnd_net_),
            .lcout(sEEACQ_i_12),
            .ltout(),
            .carryin(un5_sdacdyn_cry_11),
            .carryout(un5_sdacdyn_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_13_c_inv_LC_14_17_5.C_ON=1'b1;
    defparam un5_sdacdyn_cry_13_c_inv_LC_14_17_5.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_13_c_inv_LC_14_17_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_13_c_inv_LC_14_17_5 (
            .in0(_gnd_net_),
            .in1(N__35214),
            .in2(N__35319),
            .in3(N__35235),
            .lcout(sEEACQ_i_13),
            .ltout(),
            .carryin(un5_sdacdyn_cry_12),
            .carryout(un5_sdacdyn_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_14_c_inv_LC_14_17_6.C_ON=1'b1;
    defparam un5_sdacdyn_cry_14_c_inv_LC_14_17_6.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_14_c_inv_LC_14_17_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_14_c_inv_LC_14_17_6 (
            .in0(_gnd_net_),
            .in1(N__35203),
            .in2(N__35097),
            .in3(N__35115),
            .lcout(sEEACQ_i_14),
            .ltout(),
            .carryin(un5_sdacdyn_cry_13),
            .carryout(un5_sdacdyn_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_15_c_inv_LC_14_17_7.C_ON=1'b1;
    defparam un5_sdacdyn_cry_15_c_inv_LC_14_17_7.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_15_c_inv_LC_14_17_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_sdacdyn_cry_15_c_inv_LC_14_17_7 (
            .in0(_gnd_net_),
            .in1(N__36660),
            .in2(N__36555),
            .in3(N__36573),
            .lcout(sEEACQ_i_15),
            .ltout(),
            .carryin(un5_sdacdyn_cry_14),
            .carryout(un5_sdacdyn_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_16_c_LC_14_18_0.C_ON=1'b1;
    defparam un5_sdacdyn_cry_16_c_LC_14_18_0.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_16_c_LC_14_18_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_16_c_LC_14_18_0 (
            .in0(_gnd_net_),
            .in1(N__36541),
            .in2(N__38075),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(un5_sdacdyn_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_17_c_LC_14_18_1.C_ON=1'b1;
    defparam un5_sdacdyn_cry_17_c_LC_14_18_1.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_17_c_LC_14_18_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_17_c_LC_14_18_1 (
            .in0(_gnd_net_),
            .in1(N__36442),
            .in2(N__38079),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_16),
            .carryout(un5_sdacdyn_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_18_c_LC_14_18_2.C_ON=1'b1;
    defparam un5_sdacdyn_cry_18_c_LC_14_18_2.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_18_c_LC_14_18_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_18_c_LC_14_18_2 (
            .in0(_gnd_net_),
            .in1(N__36347),
            .in2(N__38076),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_17),
            .carryout(un5_sdacdyn_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_19_c_LC_14_18_3.C_ON=1'b1;
    defparam un5_sdacdyn_cry_19_c_LC_14_18_3.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_19_c_LC_14_18_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_19_c_LC_14_18_3 (
            .in0(_gnd_net_),
            .in1(N__36255),
            .in2(N__38080),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_18),
            .carryout(un5_sdacdyn_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_20_c_LC_14_18_4.C_ON=1'b1;
    defparam un5_sdacdyn_cry_20_c_LC_14_18_4.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_20_c_LC_14_18_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_20_c_LC_14_18_4 (
            .in0(_gnd_net_),
            .in1(N__36170),
            .in2(N__38077),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_19),
            .carryout(un5_sdacdyn_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_21_c_LC_14_18_5.C_ON=1'b1;
    defparam un5_sdacdyn_cry_21_c_LC_14_18_5.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_21_c_LC_14_18_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_21_c_LC_14_18_5 (
            .in0(_gnd_net_),
            .in1(N__36081),
            .in2(N__38081),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_20),
            .carryout(un5_sdacdyn_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_22_c_LC_14_18_6.C_ON=1'b1;
    defparam un5_sdacdyn_cry_22_c_LC_14_18_6.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_22_c_LC_14_18_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_22_c_LC_14_18_6 (
            .in0(_gnd_net_),
            .in1(N__35994),
            .in2(N__38078),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_21),
            .carryout(un5_sdacdyn_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_23_c_LC_14_18_7.C_ON=1'b1;
    defparam un5_sdacdyn_cry_23_c_LC_14_18_7.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_23_c_LC_14_18_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_sdacdyn_cry_23_c_LC_14_18_7 (
            .in0(_gnd_net_),
            .in1(N__37087),
            .in2(N__38082),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un5_sdacdyn_cry_22),
            .carryout(un5_sdacdyn_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_sdacdyn_cry_23_c_RNIELG28_LC_14_19_0.C_ON=1'b0;
    defparam un5_sdacdyn_cry_23_c_RNIELG28_LC_14_19_0.SEQ_MODE=4'b0000;
    defparam un5_sdacdyn_cry_23_c_RNIELG28_LC_14_19_0.LUT_INIT=16'b0000000010101000;
    LogicCell40 un5_sdacdyn_cry_23_c_RNIELG28_LC_14_19_0 (
            .in0(N__36993),
            .in1(N__36978),
            .in2(N__36888),
            .in3(N__36723),
            .lcout(un5_sdacdyn_cry_23_c_RNIELGZ0Z28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_pointer_0_LC_14_19_1.C_ON=1'b0;
    defparam sDAC_mem_pointer_0_LC_14_19_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_0_LC_14_19_1.LUT_INIT=16'b0111011101110111;
    LogicCell40 sDAC_mem_pointer_0_LC_14_19_1 (
            .in0(N__51541),
            .in1(N__42298),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_pointerZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53278),
            .ce(N__42232),
            .sr(N__52977));
    defparam sDAC_data_RNO_31_6_LC_14_19_3.C_ON=1'b0;
    defparam sDAC_data_RNO_31_6_LC_14_19_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_6_LC_14_19_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_31_6_LC_14_19_3 (
            .in0(N__51540),
            .in1(N__36720),
            .in2(_gnd_net_),
            .in3(N__40098),
            .lcout(sDAC_data_RNO_31Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_31_9_LC_14_19_4.C_ON=1'b0;
    defparam sDAC_data_RNO_31_9_LC_14_19_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_9_LC_14_19_4.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_31_9_LC_14_19_4 (
            .in0(N__36708),
            .in1(N__51539),
            .in2(_gnd_net_),
            .in3(N__40107),
            .lcout(sDAC_data_RNO_31Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_32_3_LC_14_19_5.C_ON=1'b0;
    defparam sDAC_data_RNO_32_3_LC_14_19_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_32_3_LC_14_19_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_32_3_LC_14_19_5 (
            .in0(N__51537),
            .in1(N__45261),
            .in2(_gnd_net_),
            .in3(N__38112),
            .lcout(sDAC_data_RNO_32Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_32_9_LC_14_19_7.C_ON=1'b0;
    defparam sDAC_data_RNO_32_9_LC_14_19_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_32_9_LC_14_19_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_32_9_LC_14_19_7 (
            .in0(N__51538),
            .in1(N__41487),
            .in2(_gnd_net_),
            .in3(N__38094),
            .lcout(sDAC_data_RNO_32Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_16_7_LC_14_20_1.C_ON=1'b0;
    defparam sDAC_mem_16_7_LC_14_20_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_7_LC_14_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_7_LC_14_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48808),
            .lcout(sDAC_mem_16Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47826),
            .ce(N__46635),
            .sr(N__52974));
    defparam sDAC_mem_16_0_LC_14_20_3.C_ON=1'b0;
    defparam sDAC_mem_16_0_LC_14_20_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_0_LC_14_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_0_LC_14_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51276),
            .lcout(sDAC_mem_16Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47826),
            .ce(N__46635),
            .sr(N__52974));
    defparam sDAC_data_RNO_29_5_LC_14_20_6.C_ON=1'b0;
    defparam sDAC_data_RNO_29_5_LC_14_20_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_5_LC_14_20_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_29_5_LC_14_20_6 (
            .in0(N__36696),
            .in1(N__51480),
            .in2(_gnd_net_),
            .in3(N__37284),
            .lcout(sDAC_data_RNO_29Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_16_2_LC_14_20_7.C_ON=1'b0;
    defparam sDAC_mem_16_2_LC_14_20_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_2_LC_14_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_2_LC_14_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50310),
            .lcout(sDAC_mem_16Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47826),
            .ce(N__46635),
            .sr(N__52974));
    defparam sDAC_mem_pointer_6_LC_15_1_1.C_ON=1'b0;
    defparam sDAC_mem_pointer_6_LC_15_1_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_6_LC_15_1_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_pointer_6_LC_15_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_mem_pointerZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53242),
            .ce(N__42231),
            .sr(N__53137));
    defparam sDAC_mem_pointer_7_LC_15_1_2.C_ON=1'b0;
    defparam sDAC_mem_pointer_7_LC_15_1_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_7_LC_15_1_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_pointer_7_LC_15_1_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_mem_pointerZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53242),
            .ce(N__42231),
            .sr(N__53137));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_0_LC_15_2_0 .C_ON=1'b1;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_0_LC_15_2_0 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_0_LC_15_2_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_0_LC_15_2_0  (
            .in0(N__37186),
            .in1(N__37240),
            .in2(N__37266),
            .in3(N__37265),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_2_0_),
            .carryout(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0 ),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53132));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_1_LC_15_2_1 .C_ON=1'b1;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_1_LC_15_2_1 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_1_LC_15_2_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_1_LC_15_2_1  (
            .in0(N__37185),
            .in1(N__37208),
            .in2(_gnd_net_),
            .in3(N__37191),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_1 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_0 ),
            .carryout(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1 ),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53132));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_2_LC_15_2_2 .C_ON=1'b1;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_2_LC_15_2_2 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_2_LC_15_2_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_2_LC_15_2_2  (
            .in0(N__37187),
            .in1(N__37139),
            .in2(_gnd_net_),
            .in3(N__37122),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_2 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_1 ),
            .carryout(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2 ),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53132));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_3_LC_15_2_3 .C_ON=1'b1;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_3_LC_15_2_3 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_3_LC_15_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_3_LC_15_2_3  (
            .in0(_gnd_net_),
            .in1(N__37119),
            .in2(_gnd_net_),
            .in3(N__37107),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_3 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_2 ),
            .carryout(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3 ),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53132));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_4_LC_15_2_4 .C_ON=1'b1;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_4_LC_15_2_4 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_4_LC_15_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_4_LC_15_2_4  (
            .in0(_gnd_net_),
            .in1(N__37104),
            .in2(_gnd_net_),
            .in3(N__37092),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_4 ),
            .ltout(),
            .carryin(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_3 ),
            .carryout(\spi_slave_inst.un1_tx_data_count_neg_sclk_i_cry_4 ),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53132));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_5_LC_15_2_5 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_5_LC_15_2_5 .SEQ_MODE=4'b1010;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_5_LC_15_2_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_5_LC_15_2_5  (
            .in0(_gnd_net_),
            .in1(N__37344),
            .in2(_gnd_net_),
            .in3(N__37347),
            .lcout(\spi_slave_inst.tx_data_count_neg_sclk_iZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVspi_slave_inst.tx_data_count_neg_sclk_i_0C_net ),
            .ce(),
            .sr(N__53132));
    defparam sDAC_mem_34_0_LC_15_3_0.C_ON=1'b0;
    defparam sDAC_mem_34_0_LC_15_3_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_0_LC_15_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_0_LC_15_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50882),
            .lcout(sDAC_mem_34Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__40089),
            .sr(N__53126));
    defparam sDAC_mem_34_2_LC_15_3_2.C_ON=1'b0;
    defparam sDAC_mem_34_2_LC_15_3_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_2_LC_15_3_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_2_LC_15_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50004),
            .lcout(sDAC_mem_34Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__40089),
            .sr(N__53126));
    defparam sDAC_mem_34_4_LC_15_3_4.C_ON=1'b0;
    defparam sDAC_mem_34_4_LC_15_3_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_4_LC_15_3_4.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_34_4_LC_15_3_4 (
            .in0(_gnd_net_),
            .in1(N__49188),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_34Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__40089),
            .sr(N__53126));
    defparam sDAC_mem_34_5_LC_15_3_5.C_ON=1'b0;
    defparam sDAC_mem_34_5_LC_15_3_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_5_LC_15_3_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_5_LC_15_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46769),
            .lcout(sDAC_mem_34Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__40089),
            .sr(N__53126));
    defparam sDAC_mem_34_6_LC_15_3_6.C_ON=1'b0;
    defparam sDAC_mem_34_6_LC_15_3_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_6_LC_15_3_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_34_6_LC_15_3_6 (
            .in0(N__47975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_34Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__40089),
            .sr(N__53126));
    defparam sDAC_mem_34_7_LC_15_3_7.C_ON=1'b0;
    defparam sDAC_mem_34_7_LC_15_3_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_7_LC_15_3_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_7_LC_15_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48545),
            .lcout(sDAC_mem_34Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47811),
            .ce(N__40089),
            .sr(N__53126));
    defparam sDAC_mem_7_0_LC_15_4_0.C_ON=1'b0;
    defparam sDAC_mem_7_0_LC_15_4_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_0_LC_15_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_7_0_LC_15_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50987),
            .lcout(sDAC_mem_7Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47800),
            .ce(N__37383),
            .sr(N__53111));
    defparam sDAC_mem_7_1_LC_15_4_1.C_ON=1'b0;
    defparam sDAC_mem_7_1_LC_15_4_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_1_LC_15_4_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_7_1_LC_15_4_1 (
            .in0(N__50601),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_7Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47800),
            .ce(N__37383),
            .sr(N__53111));
    defparam sDAC_mem_7_2_LC_15_4_2.C_ON=1'b0;
    defparam sDAC_mem_7_2_LC_15_4_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_2_LC_15_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_7_2_LC_15_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50107),
            .lcout(sDAC_mem_7Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47800),
            .ce(N__37383),
            .sr(N__53111));
    defparam sDAC_mem_7_3_LC_15_4_3.C_ON=1'b0;
    defparam sDAC_mem_7_3_LC_15_4_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_3_LC_15_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_7_3_LC_15_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49609),
            .lcout(sDAC_mem_7Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47800),
            .ce(N__37383),
            .sr(N__53111));
    defparam sDAC_mem_7_4_LC_15_4_4.C_ON=1'b0;
    defparam sDAC_mem_7_4_LC_15_4_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_4_LC_15_4_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_7_4_LC_15_4_4 (
            .in0(N__49186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_7Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47800),
            .ce(N__37383),
            .sr(N__53111));
    defparam sDAC_mem_7_5_LC_15_4_5.C_ON=1'b0;
    defparam sDAC_mem_7_5_LC_15_4_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_5_LC_15_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_7_5_LC_15_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46876),
            .lcout(sDAC_mem_7Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47800),
            .ce(N__37383),
            .sr(N__53111));
    defparam sDAC_mem_7_6_LC_15_4_6.C_ON=1'b0;
    defparam sDAC_mem_7_6_LC_15_4_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_6_LC_15_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_7_6_LC_15_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48189),
            .lcout(sDAC_mem_7Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47800),
            .ce(N__37383),
            .sr(N__53111));
    defparam sDAC_mem_7_7_LC_15_4_7.C_ON=1'b0;
    defparam sDAC_mem_7_7_LC_15_4_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_7_7_LC_15_4_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_7_7_LC_15_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48746),
            .lcout(sDAC_mem_7Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47800),
            .ce(N__37383),
            .sr(N__53111));
    defparam sDAC_mem_5_0_LC_15_5_0.C_ON=1'b0;
    defparam sDAC_mem_5_0_LC_15_5_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_0_LC_15_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_0_LC_15_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51099),
            .lcout(sDAC_mem_5Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47785),
            .ce(N__37395),
            .sr(N__53099));
    defparam sDAC_mem_5_1_LC_15_5_1.C_ON=1'b0;
    defparam sDAC_mem_5_1_LC_15_5_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_1_LC_15_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_1_LC_15_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50685),
            .lcout(sDAC_mem_5Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47785),
            .ce(N__37395),
            .sr(N__53099));
    defparam sDAC_mem_5_2_LC_15_5_2.C_ON=1'b0;
    defparam sDAC_mem_5_2_LC_15_5_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_2_LC_15_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_2_LC_15_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50108),
            .lcout(sDAC_mem_5Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47785),
            .ce(N__37395),
            .sr(N__53099));
    defparam sDAC_mem_5_3_LC_15_5_3.C_ON=1'b0;
    defparam sDAC_mem_5_3_LC_15_5_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_3_LC_15_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_3_LC_15_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49610),
            .lcout(sDAC_mem_5Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47785),
            .ce(N__37395),
            .sr(N__53099));
    defparam sDAC_mem_5_4_LC_15_5_4.C_ON=1'b0;
    defparam sDAC_mem_5_4_LC_15_5_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_4_LC_15_5_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_5_4_LC_15_5_4 (
            .in0(N__49187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_5Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47785),
            .ce(N__37395),
            .sr(N__53099));
    defparam sDAC_mem_5_5_LC_15_5_5.C_ON=1'b0;
    defparam sDAC_mem_5_5_LC_15_5_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_5_LC_15_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_5_LC_15_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46878),
            .lcout(sDAC_mem_5Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47785),
            .ce(N__37395),
            .sr(N__53099));
    defparam sDAC_mem_5_6_LC_15_5_6.C_ON=1'b0;
    defparam sDAC_mem_5_6_LC_15_5_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_6_LC_15_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_6_LC_15_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48191),
            .lcout(sDAC_mem_5Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47785),
            .ce(N__37395),
            .sr(N__53099));
    defparam sDAC_mem_5_7_LC_15_5_7.C_ON=1'b0;
    defparam sDAC_mem_5_7_LC_15_5_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_5_7_LC_15_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_5_7_LC_15_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48747),
            .lcout(sDAC_mem_5Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47785),
            .ce(N__37395),
            .sr(N__53099));
    defparam sAddress_RNI9IH12_10_3_LC_15_6_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_10_3_LC_15_6_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_10_3_LC_15_6_0.LUT_INIT=16'b0000010000000000;
    LogicCell40 sAddress_RNI9IH12_10_3_LC_15_6_0 (
            .in0(N__40584),
            .in1(N__40398),
            .in2(N__46449),
            .in3(N__37494),
            .lcout(sDAC_mem_2_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_17_3_LC_15_6_1.C_ON=1'b0;
    defparam sAddress_RNI9IH12_17_3_LC_15_6_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_17_3_LC_15_6_1.LUT_INIT=16'b0000000000100000;
    LogicCell40 sAddress_RNI9IH12_17_3_LC_15_6_1 (
            .in0(N__37490),
            .in1(N__40585),
            .in2(N__46246),
            .in3(N__40401),
            .lcout(sDAC_mem_5_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_15_3_LC_15_6_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_15_3_LC_15_6_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_15_3_LC_15_6_2.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNI9IH12_15_3_LC_15_6_2 (
            .in0(N__40583),
            .in1(N__40397),
            .in2(N__44586),
            .in3(N__37489),
            .lcout(sDAC_mem_7_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_2_3_LC_15_6_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_2_3_LC_15_6_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_2_3_LC_15_6_3.LUT_INIT=16'b0010000000000000;
    LogicCell40 sAddress_RNI9IH12_2_3_LC_15_6_3 (
            .in0(N__37492),
            .in1(N__40586),
            .in2(N__44587),
            .in3(N__40402),
            .lcout(sDAC_mem_8_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_19_3_LC_15_6_4.C_ON=1'b0;
    defparam sAddress_RNI9IH12_19_3_LC_15_6_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_19_3_LC_15_6_4.LUT_INIT=16'b0000001000000000;
    LogicCell40 sAddress_RNI9IH12_19_3_LC_15_6_4 (
            .in0(N__43282),
            .in1(N__40396),
            .in2(N__40604),
            .in3(N__37491),
            .lcout(sDAC_mem_3_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_4_3_LC_15_6_5.C_ON=1'b0;
    defparam sAddress_RNI9IH12_4_3_LC_15_6_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_4_3_LC_15_6_5.LUT_INIT=16'b0010000000000000;
    LogicCell40 sAddress_RNI9IH12_4_3_LC_15_6_5 (
            .in0(N__37493),
            .in1(N__40582),
            .in2(N__46245),
            .in3(N__40399),
            .lcout(sDAC_mem_6_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIVREN1_1_4_LC_15_6_6.C_ON=1'b0;
    defparam sAddress_RNIVREN1_1_4_LC_15_6_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNIVREN1_1_4_LC_15_6_6.LUT_INIT=16'b0100000000000000;
    LogicCell40 sAddress_RNIVREN1_1_4_LC_15_6_6 (
            .in0(N__46528),
            .in1(N__44645),
            .in2(N__44808),
            .in3(N__44741),
            .lcout(N_279),
            .ltout(N_279_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_6_3_LC_15_6_7.C_ON=1'b0;
    defparam sAddress_RNI9IH12_6_3_LC_15_6_7.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_6_3_LC_15_6_7.LUT_INIT=16'b0100000000000000;
    LogicCell40 sAddress_RNI9IH12_6_3_LC_15_6_7 (
            .in0(N__40575),
            .in1(N__40400),
            .in2(N__37473),
            .in3(N__43283),
            .lcout(sDAC_mem_4_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_7_LC_15_7_0.C_ON=1'b0;
    defparam sDAC_data_RNO_10_7_LC_15_7_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_7_LC_15_7_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_10_7_LC_15_7_0 (
            .in0(N__37470),
            .in1(N__38790),
            .in2(N__45875),
            .in3(N__38862),
            .lcout(sDAC_data_RNO_10Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_7_LC_15_7_2.C_ON=1'b0;
    defparam sDAC_data_RNO_6_7_LC_15_7_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_7_LC_15_7_2.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_6_7_LC_15_7_2 (
            .in0(N__45803),
            .in1(N__45520),
            .in2(N__42093),
            .in3(N__39072),
            .lcout(),
            .ltout(sDAC_data_2_14_ns_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_7_LC_15_7_3.C_ON=1'b0;
    defparam sDAC_data_RNO_1_7_LC_15_7_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_7_LC_15_7_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_1_7_LC_15_7_3 (
            .in0(N__45867),
            .in1(N__38892),
            .in2(N__37461),
            .in3(N__37458),
            .lcout(sDAC_data_RNO_1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_7_LC_15_7_4.C_ON=1'b0;
    defparam sDAC_data_RNO_3_7_LC_15_7_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_7_LC_15_7_4.LUT_INIT=16'b0010010101110101;
    LogicCell40 sDAC_data_RNO_3_7_LC_15_7_4 (
            .in0(N__42631),
            .in1(N__38469),
            .in2(N__42534),
            .in3(N__37449),
            .lcout(),
            .ltout(sDAC_data_2_41_ns_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_7_LC_15_7_5.C_ON=1'b0;
    defparam sDAC_data_RNO_0_7_LC_15_7_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_7_LC_15_7_5.LUT_INIT=16'b0101111000001110;
    LogicCell40 sDAC_data_RNO_0_7_LC_15_7_5 (
            .in0(N__42518),
            .in1(N__37443),
            .in2(N__37437),
            .in3(N__37434),
            .lcout(),
            .ltout(sDAC_data_2_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_7_LC_15_7_6.C_ON=1'b0;
    defparam sDAC_data_7_LC_15_7_6.SEQ_MODE=4'b1010;
    defparam sDAC_data_7_LC_15_7_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 sDAC_data_7_LC_15_7_6 (
            .in0(N__45960),
            .in1(_gnd_net_),
            .in2(N__37428),
            .in3(N__42382),
            .lcout(sDAC_dataZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53252),
            .ce(N__42229),
            .sr(N__53074));
    defparam sDAC_data_RNO_17_9_LC_15_8_1.C_ON=1'b0;
    defparam sDAC_data_RNO_17_9_LC_15_8_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_9_LC_15_8_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_9_LC_15_8_1 (
            .in0(N__43581),
            .in1(N__44367),
            .in2(_gnd_net_),
            .in3(N__44271),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_9_LC_15_8_2.C_ON=1'b0;
    defparam sDAC_data_RNO_8_9_LC_15_8_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_9_LC_15_8_2.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_8_9_LC_15_8_2 (
            .in0(_gnd_net_),
            .in1(N__51808),
            .in2(N__37539),
            .in3(N__45156),
            .lcout(),
            .ltout(sDAC_data_RNO_8Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_9_LC_15_8_3.C_ON=1'b0;
    defparam sDAC_data_RNO_2_9_LC_15_8_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_9_LC_15_8_3.LUT_INIT=16'b0111011000110010;
    LogicCell40 sDAC_data_RNO_2_9_LC_15_8_3 (
            .in0(N__45751),
            .in1(N__38295),
            .in2(N__37536),
            .in3(N__37530),
            .lcout(sDAC_data_RNO_2Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_3_4_LC_15_8_4.C_ON=1'b0;
    defparam sDAC_mem_3_4_LC_15_8_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_4_LC_15_8_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_3_4_LC_15_8_4 (
            .in0(N__49260),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_3Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47746),
            .ce(N__42961),
            .sr(N__53062));
    defparam sDAC_data_RNO_16_9_LC_15_8_5.C_ON=1'b0;
    defparam sDAC_data_RNO_16_9_LC_15_8_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_9_LC_15_8_5.LUT_INIT=16'b0011000100111101;
    LogicCell40 sDAC_data_RNO_16_9_LC_15_8_5 (
            .in0(N__38817),
            .in1(N__43580),
            .in2(N__52012),
            .in3(N__41796),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_9_LC_15_8_6.C_ON=1'b0;
    defparam sDAC_data_RNO_7_9_LC_15_8_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_9_LC_15_8_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_7_9_LC_15_8_6 (
            .in0(N__52119),
            .in1(N__44232),
            .in2(N__37533),
            .in3(N__46650),
            .lcout(sDAC_data_RNO_7Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_29_7_LC_15_9_2.C_ON=1'b0;
    defparam sDAC_data_RNO_29_7_LC_15_9_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_7_LC_15_9_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_29_7_LC_15_9_2 (
            .in0(N__37524),
            .in1(N__52014),
            .in2(_gnd_net_),
            .in3(N__37515),
            .lcout(sDAC_data_RNO_29Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_16_4_LC_15_9_3.C_ON=1'b0;
    defparam sDAC_mem_16_4_LC_15_9_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_4_LC_15_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_4_LC_15_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49360),
            .lcout(sDAC_mem_16Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47735),
            .ce(N__46629),
            .sr(N__53052));
    defparam sDAC_data_RNO_29_8_LC_15_9_4.C_ON=1'b0;
    defparam sDAC_data_RNO_29_8_LC_15_9_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_8_LC_15_9_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_29_8_LC_15_9_4 (
            .in0(N__37509),
            .in1(N__52013),
            .in2(_gnd_net_),
            .in3(N__37500),
            .lcout(sDAC_data_RNO_29Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_16_5_LC_15_9_5.C_ON=1'b0;
    defparam sDAC_mem_16_5_LC_15_9_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_5_LC_15_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_5_LC_15_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47017),
            .lcout(sDAC_mem_16Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47735),
            .ce(N__46629),
            .sr(N__53052));
    defparam sDAC_data_RNO_29_9_LC_15_9_6.C_ON=1'b0;
    defparam sDAC_data_RNO_29_9_LC_15_9_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_9_LC_15_9_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_29_9_LC_15_9_6 (
            .in0(N__37569),
            .in1(N__52015),
            .in2(_gnd_net_),
            .in3(N__37560),
            .lcout(sDAC_data_RNO_29Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_16_6_LC_15_9_7.C_ON=1'b0;
    defparam sDAC_mem_16_6_LC_15_9_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_6_LC_15_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_6_LC_15_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48234),
            .lcout(sDAC_mem_16Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47735),
            .ce(N__46629),
            .sr(N__53052));
    defparam sDAC_mem_pointer_RNI3NFH_1_LC_15_10_0.C_ON=1'b1;
    defparam sDAC_mem_pointer_RNI3NFH_1_LC_15_10_0.SEQ_MODE=4'b0000;
    defparam sDAC_mem_pointer_RNI3NFH_1_LC_15_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 sDAC_mem_pointer_RNI3NFH_1_LC_15_10_0 (
            .in0(_gnd_net_),
            .in1(N__52041),
            .in2(N__45491),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(sDAC_mem_pointer_0_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_pointer_2_LC_15_10_1.C_ON=1'b1;
    defparam sDAC_mem_pointer_2_LC_15_10_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_2_LC_15_10_1.LUT_INIT=16'b0010001010001000;
    LogicCell40 sDAC_mem_pointer_2_LC_15_10_1 (
            .in0(N__42373),
            .in1(N__45717),
            .in2(_gnd_net_),
            .in3(N__37554),
            .lcout(sDAC_mem_pointerZ0Z_2),
            .ltout(),
            .carryin(sDAC_mem_pointer_0_cry_1),
            .carryout(sDAC_mem_pointer_0_cry_2),
            .clk(N__53254),
            .ce(N__42225),
            .sr(N__53042));
    defparam sDAC_mem_pointer_3_LC_15_10_2.C_ON=1'b1;
    defparam sDAC_mem_pointer_3_LC_15_10_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_3_LC_15_10_2.LUT_INIT=16'b0010001010001000;
    LogicCell40 sDAC_mem_pointer_3_LC_15_10_2 (
            .in0(N__42376),
            .in1(N__42623),
            .in2(_gnd_net_),
            .in3(N__37551),
            .lcout(sDAC_mem_pointerZ0Z_3),
            .ltout(),
            .carryin(sDAC_mem_pointer_0_cry_2),
            .carryout(sDAC_mem_pointer_0_cry_3),
            .clk(N__53254),
            .ce(N__42225),
            .sr(N__53042));
    defparam sDAC_mem_pointer_4_LC_15_10_3.C_ON=1'b1;
    defparam sDAC_mem_pointer_4_LC_15_10_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_4_LC_15_10_3.LUT_INIT=16'b0010001010001000;
    LogicCell40 sDAC_mem_pointer_4_LC_15_10_3 (
            .in0(N__42374),
            .in1(N__42483),
            .in2(_gnd_net_),
            .in3(N__37548),
            .lcout(sDAC_mem_pointerZ0Z_4),
            .ltout(),
            .carryin(sDAC_mem_pointer_0_cry_3),
            .carryout(sDAC_mem_pointer_0_cry_4),
            .clk(N__53254),
            .ce(N__42225),
            .sr(N__53042));
    defparam sDAC_mem_pointer_5_LC_15_10_4.C_ON=1'b0;
    defparam sDAC_mem_pointer_5_LC_15_10_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_5_LC_15_10_4.LUT_INIT=16'b0100010010001000;
    LogicCell40 sDAC_mem_pointer_5_LC_15_10_4 (
            .in0(N__43479),
            .in1(N__42375),
            .in2(_gnd_net_),
            .in3(N__37545),
            .lcout(sDAC_mem_pointerZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53254),
            .ce(N__42225),
            .sr(N__53042));
    defparam sDAC_data_RNO_23_9_LC_15_11_1.C_ON=1'b0;
    defparam sDAC_data_RNO_23_9_LC_15_11_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_9_LC_15_11_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_9_LC_15_11_1 (
            .in0(N__52017),
            .in1(N__38355),
            .in2(_gnd_net_),
            .in3(N__37629),
            .lcout(),
            .ltout(sDAC_data_RNO_23Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_9_LC_15_11_2.C_ON=1'b0;
    defparam sDAC_data_RNO_11_9_LC_15_11_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_9_LC_15_11_2.LUT_INIT=16'b1010000011011101;
    LogicCell40 sDAC_data_RNO_11_9_LC_15_11_2 (
            .in0(N__45709),
            .in1(N__38169),
            .in2(N__37542),
            .in3(N__38121),
            .lcout(sDAC_data_RNO_11Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_10_LC_15_11_3.C_ON=1'b0;
    defparam sDAC_data_RNO_8_10_LC_15_11_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_10_LC_15_11_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_8_10_LC_15_11_3 (
            .in0(N__37653),
            .in1(N__52019),
            .in2(_gnd_net_),
            .in3(N__45141),
            .lcout(),
            .ltout(sDAC_data_RNO_8Z0Z_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_10_LC_15_11_4.C_ON=1'b0;
    defparam sDAC_data_RNO_2_10_LC_15_11_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_10_LC_15_11_4.LUT_INIT=16'b0111011000110010;
    LogicCell40 sDAC_data_RNO_2_10_LC_15_11_4 (
            .in0(N__45710),
            .in1(N__37647),
            .in2(N__37641),
            .in3(N__37635),
            .lcout(sDAC_data_RNO_2Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_10_LC_15_11_5.C_ON=1'b0;
    defparam sDAC_data_RNO_16_10_LC_15_11_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_10_LC_15_11_5.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_16_10_LC_15_11_5 (
            .in0(N__52016),
            .in1(N__41997),
            .in2(N__43575),
            .in3(N__38808),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_10_LC_15_11_6.C_ON=1'b0;
    defparam sDAC_data_RNO_7_10_LC_15_11_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_10_LC_15_11_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_7_10_LC_15_11_6 (
            .in0(N__52018),
            .in1(N__44220),
            .in2(N__37638),
            .in3(N__47340),
            .lcout(sDAC_data_RNO_7Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_28_6_LC_15_11_7.C_ON=1'b0;
    defparam sDAC_mem_28_6_LC_15_11_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_6_LC_15_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_6_LC_15_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48310),
            .lcout(sDAC_mem_28Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47718),
            .ce(N__41772),
            .sr(N__53033));
    defparam sDAC_mem_pointer_1_LC_15_12_0.C_ON=1'b0;
    defparam sDAC_mem_pointer_1_LC_15_12_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_pointer_1_LC_15_12_0.LUT_INIT=16'b0110011000000000;
    LogicCell40 sDAC_mem_pointer_1_LC_15_12_0 (
            .in0(N__45424),
            .in1(N__52064),
            .in2(_gnd_net_),
            .in3(N__42379),
            .lcout(sDAC_mem_pointerZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53263),
            .ce(N__42228),
            .sr(N__53023));
    defparam sDAC_data_1_LC_15_12_2.C_ON=1'b0;
    defparam sDAC_data_1_LC_15_12_2.SEQ_MODE=4'b1010;
    defparam sDAC_data_1_LC_15_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_1_LC_15_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53263),
            .ce(N__42228),
            .sr(N__53023));
    defparam sDAC_data_11_LC_15_12_3.C_ON=1'b0;
    defparam sDAC_data_11_LC_15_12_3.SEQ_MODE=4'b1010;
    defparam sDAC_data_11_LC_15_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_11_LC_15_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53263),
            .ce(N__42228),
            .sr(N__53023));
    defparam sDAC_data_12_LC_15_12_4.C_ON=1'b0;
    defparam sDAC_data_12_LC_15_12_4.SEQ_MODE=4'b1010;
    defparam sDAC_data_12_LC_15_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_12_LC_15_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38018),
            .lcout(sDAC_dataZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53263),
            .ce(N__42228),
            .sr(N__53023));
    defparam sDAC_data_13_LC_15_12_5.C_ON=1'b0;
    defparam sDAC_data_13_LC_15_12_5.SEQ_MODE=4'b1010;
    defparam sDAC_data_13_LC_15_12_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_data_13_LC_15_12_5 (
            .in0(N__38019),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_dataZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53263),
            .ce(N__42228),
            .sr(N__53023));
    defparam sDAC_data_14_LC_15_12_6.C_ON=1'b0;
    defparam sDAC_data_14_LC_15_12_6.SEQ_MODE=4'b1010;
    defparam sDAC_data_14_LC_15_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_14_LC_15_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53263),
            .ce(N__42228),
            .sr(N__53023));
    defparam sDAC_data_15_LC_15_12_7.C_ON=1'b0;
    defparam sDAC_data_15_LC_15_12_7.SEQ_MODE=4'b1010;
    defparam sDAC_data_15_LC_15_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_data_15_LC_15_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(sDAC_dataZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53263),
            .ce(N__42228),
            .sr(N__53023));
    defparam sDAC_data_RNO_31_8_LC_15_13_0.C_ON=1'b0;
    defparam sDAC_data_RNO_31_8_LC_15_13_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_8_LC_15_13_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_31_8_LC_15_13_0 (
            .in0(N__40128),
            .in1(N__51880),
            .in2(_gnd_net_),
            .in3(N__38157),
            .lcout(),
            .ltout(sDAC_data_RNO_31Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_25_8_LC_15_13_1.C_ON=1'b0;
    defparam sDAC_data_RNO_25_8_LC_15_13_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_8_LC_15_13_1.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_25_8_LC_15_13_1 (
            .in0(N__45848),
            .in1(N__45415),
            .in2(N__37683),
            .in3(N__37677),
            .lcout(),
            .ltout(sDAC_data_2_39_ns_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_8_LC_15_13_2.C_ON=1'b0;
    defparam sDAC_data_RNO_11_8_LC_15_13_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_8_LC_15_13_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_11_8_LC_15_13_2 (
            .in0(N__45828),
            .in1(N__37659),
            .in2(N__37680),
            .in3(N__37671),
            .lcout(sDAC_data_RNO_11Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_32_8_LC_15_13_3.C_ON=1'b0;
    defparam sDAC_data_RNO_32_8_LC_15_13_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_32_8_LC_15_13_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_32_8_LC_15_13_3 (
            .in0(N__51878),
            .in1(N__41499),
            .in2(_gnd_net_),
            .in3(N__38100),
            .lcout(sDAC_data_RNO_32Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_8_LC_15_13_4.C_ON=1'b0;
    defparam sDAC_data_RNO_23_8_LC_15_13_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_8_LC_15_13_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_8_LC_15_13_4 (
            .in0(N__51881),
            .in1(N__38364),
            .in2(_gnd_net_),
            .in3(N__41511),
            .lcout(sDAC_data_RNO_23Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_8_LC_15_13_5.C_ON=1'b0;
    defparam sDAC_data_RNO_24_8_LC_15_13_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_8_LC_15_13_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_8_LC_15_13_5 (
            .in0(N__51879),
            .in1(N__37665),
            .in2(_gnd_net_),
            .in3(N__39708),
            .lcout(sDAC_data_RNO_24Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_24_5_LC_15_13_6.C_ON=1'b0;
    defparam sDAC_mem_24_5_LC_15_13_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_5_LC_15_13_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_5_LC_15_13_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47117),
            .lcout(sDAC_mem_24Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47736),
            .ce(N__39971),
            .sr(N__53018));
    defparam sDAC_data_RNO_25_9_LC_15_13_7.C_ON=1'b0;
    defparam sDAC_data_RNO_25_9_LC_15_13_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_9_LC_15_13_7.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_25_9_LC_15_13_7 (
            .in0(N__45847),
            .in1(N__45414),
            .in2(N__38151),
            .in3(N__38133),
            .lcout(sDAC_data_2_39_ns_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_26_0_LC_15_14_0.C_ON=1'b0;
    defparam sDAC_mem_26_0_LC_15_14_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_0_LC_15_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_26_0_LC_15_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51247),
            .lcout(sDAC_mem_26Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47747),
            .ce(N__39528),
            .sr(N__53012));
    defparam sDAC_mem_26_1_LC_15_14_1.C_ON=1'b0;
    defparam sDAC_mem_26_1_LC_15_14_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_1_LC_15_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_26_1_LC_15_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50723),
            .lcout(sDAC_mem_26Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47747),
            .ce(N__39528),
            .sr(N__53012));
    defparam sDAC_mem_26_2_LC_15_14_2.C_ON=1'b0;
    defparam sDAC_mem_26_2_LC_15_14_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_2_LC_15_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_26_2_LC_15_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50263),
            .lcout(sDAC_mem_26Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47747),
            .ce(N__39528),
            .sr(N__53012));
    defparam sDAC_mem_26_3_LC_15_14_3.C_ON=1'b0;
    defparam sDAC_mem_26_3_LC_15_14_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_3_LC_15_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_26_3_LC_15_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49797),
            .lcout(sDAC_mem_26Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47747),
            .ce(N__39528),
            .sr(N__53012));
    defparam sDAC_mem_26_4_LC_15_14_4.C_ON=1'b0;
    defparam sDAC_mem_26_4_LC_15_14_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_4_LC_15_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_26_4_LC_15_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49177),
            .lcout(sDAC_mem_26Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47747),
            .ce(N__39528),
            .sr(N__53012));
    defparam sDAC_mem_26_5_LC_15_14_5.C_ON=1'b0;
    defparam sDAC_mem_26_5_LC_15_14_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_5_LC_15_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_26_5_LC_15_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47074),
            .lcout(sDAC_mem_26Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47747),
            .ce(N__39528),
            .sr(N__53012));
    defparam sDAC_mem_26_6_LC_15_14_6.C_ON=1'b0;
    defparam sDAC_mem_26_6_LC_15_14_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_6_LC_15_14_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_26_6_LC_15_14_6 (
            .in0(N__48311),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_26Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47747),
            .ce(N__39528),
            .sr(N__53012));
    defparam sDAC_mem_26_7_LC_15_14_7.C_ON=1'b0;
    defparam sDAC_mem_26_7_LC_15_14_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_26_7_LC_15_14_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_26_7_LC_15_14_7 (
            .in0(N__48843),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_26Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47747),
            .ce(N__39528),
            .sr(N__53012));
    defparam sDAC_data_RNO_19_9_LC_15_15_0.C_ON=1'b0;
    defparam sDAC_data_RNO_19_9_LC_15_15_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_9_LC_15_15_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_9_LC_15_15_0 (
            .in0(N__52112),
            .in1(N__45036),
            .in2(_gnd_net_),
            .in3(N__43947),
            .lcout(sDAC_data_RNO_19Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_9_LC_15_15_1.C_ON=1'b0;
    defparam sDAC_data_RNO_18_9_LC_15_15_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_9_LC_15_15_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_9_LC_15_15_1 (
            .in0(N__52114),
            .in1(N__45234),
            .in2(_gnd_net_),
            .in3(N__47868),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_9_LC_15_15_2.C_ON=1'b0;
    defparam sDAC_data_RNO_9_9_LC_15_15_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_9_LC_15_15_2.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_9_9_LC_15_15_2 (
            .in0(N__45736),
            .in1(N__45439),
            .in2(N__38304),
            .in3(N__38301),
            .lcout(sDAC_data_2_24_ns_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEADC_freq_RNISBIA1_0_LC_15_15_4.C_ON=1'b0;
    defparam sEEADC_freq_RNISBIA1_0_LC_15_15_4.SEQ_MODE=4'b0000;
    defparam sEEADC_freq_RNISBIA1_0_LC_15_15_4.LUT_INIT=16'b1000001001000001;
    LogicCell40 sEEADC_freq_RNISBIA1_0_LC_15_15_4 (
            .in0(N__41460),
            .in1(N__38283),
            .in2(N__44142),
            .in3(N__38268),
            .lcout(),
            .ltout(un11_sacqtime_NE_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEADC_freq_RNI01BA5_0_LC_15_15_5.C_ON=1'b0;
    defparam sEEADC_freq_RNI01BA5_0_LC_15_15_5.SEQ_MODE=4'b0000;
    defparam sEEADC_freq_RNI01BA5_0_LC_15_15_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 sEEADC_freq_RNI01BA5_0_LC_15_15_5 (
            .in0(N__38253),
            .in1(N__38247),
            .in2(N__38241),
            .in3(N__38238),
            .lcout(un11_sacqtime_NE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_9_LC_15_15_7.C_ON=1'b0;
    defparam sDAC_data_RNO_24_9_LC_15_15_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_9_LC_15_15_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_24_9_LC_15_15_7 (
            .in0(N__38175),
            .in1(N__52113),
            .in2(_gnd_net_),
            .in3(N__39699),
            .lcout(sDAC_data_RNO_24Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_29_0_LC_15_16_0.C_ON=1'b0;
    defparam sDAC_mem_29_0_LC_15_16_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_0_LC_15_16_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_29_0_LC_15_16_0 (
            .in0(N__51253),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_29Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47770),
            .ce(N__38346),
            .sr(N__52994));
    defparam sDAC_mem_29_1_LC_15_16_1.C_ON=1'b0;
    defparam sDAC_mem_29_1_LC_15_16_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_1_LC_15_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_29_1_LC_15_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50754),
            .lcout(sDAC_mem_29Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47770),
            .ce(N__38346),
            .sr(N__52994));
    defparam sDAC_mem_29_2_LC_15_16_2.C_ON=1'b0;
    defparam sDAC_mem_29_2_LC_15_16_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_2_LC_15_16_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_29_2_LC_15_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50300),
            .lcout(sDAC_mem_29Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47770),
            .ce(N__38346),
            .sr(N__52994));
    defparam sDAC_mem_29_3_LC_15_16_3.C_ON=1'b0;
    defparam sDAC_mem_29_3_LC_15_16_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_3_LC_15_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_29_3_LC_15_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49835),
            .lcout(sDAC_mem_29Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47770),
            .ce(N__38346),
            .sr(N__52994));
    defparam sDAC_mem_29_4_LC_15_16_4.C_ON=1'b0;
    defparam sDAC_mem_29_4_LC_15_16_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_4_LC_15_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_29_4_LC_15_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49326),
            .lcout(sDAC_mem_29Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47770),
            .ce(N__38346),
            .sr(N__52994));
    defparam sDAC_mem_29_5_LC_15_16_5.C_ON=1'b0;
    defparam sDAC_mem_29_5_LC_15_16_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_5_LC_15_16_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_29_5_LC_15_16_5 (
            .in0(N__47134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_29Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47770),
            .ce(N__38346),
            .sr(N__52994));
    defparam sDAC_mem_29_6_LC_15_16_6.C_ON=1'b0;
    defparam sDAC_mem_29_6_LC_15_16_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_6_LC_15_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_29_6_LC_15_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48337),
            .lcout(sDAC_mem_29Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47770),
            .ce(N__38346),
            .sr(N__52994));
    defparam sDAC_mem_29_7_LC_15_16_7.C_ON=1'b0;
    defparam sDAC_mem_29_7_LC_15_16_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_29_7_LC_15_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_29_7_LC_15_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48830),
            .lcout(sDAC_mem_29Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47770),
            .ce(N__38346),
            .sr(N__52994));
    defparam sDAC_data_RNO_11_6_LC_15_17_0.C_ON=1'b0;
    defparam sDAC_data_RNO_11_6_LC_15_17_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_6_LC_15_17_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_11_6_LC_15_17_0 (
            .in0(N__38424),
            .in1(N__38325),
            .in2(N__45841),
            .in3(N__38664),
            .lcout(sDAC_data_RNO_11Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_6_LC_15_17_1.C_ON=1'b0;
    defparam sDAC_data_RNO_23_6_LC_15_17_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_6_LC_15_17_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_6_LC_15_17_1 (
            .in0(N__52075),
            .in1(N__38331),
            .in2(_gnd_net_),
            .in3(N__38457),
            .lcout(sDAC_data_RNO_23Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_31_7_LC_15_17_2.C_ON=1'b0;
    defparam sDAC_data_RNO_31_7_LC_15_17_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_7_LC_15_17_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_31_7_LC_15_17_2 (
            .in0(N__51892),
            .in1(N__38319),
            .in2(_gnd_net_),
            .in3(N__39897),
            .lcout(),
            .ltout(sDAC_data_RNO_31Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_25_7_LC_15_17_3.C_ON=1'b0;
    defparam sDAC_data_RNO_25_7_LC_15_17_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_7_LC_15_17_3.LUT_INIT=16'b0100010101100111;
    LogicCell40 sDAC_data_RNO_25_7_LC_15_17_3 (
            .in0(N__45440),
            .in1(N__45746),
            .in2(N__38307),
            .in3(N__38442),
            .lcout(),
            .ltout(sDAC_data_2_39_ns_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_7_LC_15_17_4.C_ON=1'b0;
    defparam sDAC_data_RNO_11_7_LC_15_17_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_7_LC_15_17_4.LUT_INIT=16'b1100101100001011;
    LogicCell40 sDAC_data_RNO_11_7_LC_15_17_4 (
            .in0(N__39744),
            .in1(N__45750),
            .in2(N__38472),
            .in3(N__38649),
            .lcout(sDAC_data_RNO_11Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_28_3_LC_15_17_5.C_ON=1'b0;
    defparam sDAC_mem_28_3_LC_15_17_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_3_LC_15_17_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_28_3_LC_15_17_5 (
            .in0(N__49837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_28Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47786),
            .ce(N__41778),
            .sr(N__52989));
    defparam sDAC_data_RNO_32_7_LC_15_17_6.C_ON=1'b0;
    defparam sDAC_data_RNO_32_7_LC_15_17_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_32_7_LC_15_17_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_32_7_LC_15_17_6 (
            .in0(N__51891),
            .in1(N__41226),
            .in2(_gnd_net_),
            .in3(N__38451),
            .lcout(sDAC_data_RNO_32Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_6_LC_15_17_7.C_ON=1'b0;
    defparam sDAC_data_RNO_24_6_LC_15_17_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_6_LC_15_17_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_6_LC_15_17_7 (
            .in0(N__52074),
            .in1(N__38436),
            .in2(_gnd_net_),
            .in3(N__39720),
            .lcout(sDAC_data_RNO_24Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_31_5_LC_15_18_0.C_ON=1'b0;
    defparam sDAC_data_RNO_31_5_LC_15_18_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_5_LC_15_18_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_31_5_LC_15_18_0 (
            .in0(N__51495),
            .in1(N__38679),
            .in2(_gnd_net_),
            .in3(N__40134),
            .lcout(),
            .ltout(sDAC_data_RNO_31Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_25_5_LC_15_18_1.C_ON=1'b0;
    defparam sDAC_data_RNO_25_5_LC_15_18_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_5_LC_15_18_1.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_25_5_LC_15_18_1 (
            .in0(N__45734),
            .in1(N__45521),
            .in2(N__38418),
            .in3(N__38388),
            .lcout(),
            .ltout(sDAC_data_2_39_ns_1_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_5_LC_15_18_2.C_ON=1'b0;
    defparam sDAC_data_RNO_11_5_LC_15_18_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_5_LC_15_18_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_11_5_LC_15_18_2 (
            .in0(N__45737),
            .in1(N__38685),
            .in2(N__38415),
            .in3(N__38370),
            .lcout(sDAC_data_RNO_11Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_32_5_LC_15_18_3.C_ON=1'b0;
    defparam sDAC_data_RNO_32_5_LC_15_18_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_32_5_LC_15_18_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_32_5_LC_15_18_3 (
            .in0(N__41256),
            .in1(N__51493),
            .in2(_gnd_net_),
            .in3(N__38397),
            .lcout(sDAC_data_RNO_32Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_5_LC_15_18_4.C_ON=1'b0;
    defparam sDAC_data_RNO_23_5_LC_15_18_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_5_LC_15_18_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_5_LC_15_18_4 (
            .in0(N__51494),
            .in1(N__38379),
            .in2(_gnd_net_),
            .in3(N__41535),
            .lcout(sDAC_data_RNO_23Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_5_LC_15_18_5.C_ON=1'b0;
    defparam sDAC_data_RNO_24_5_LC_15_18_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_5_LC_15_18_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_5_LC_15_18_5 (
            .in0(N__51501),
            .in1(N__38697),
            .in2(_gnd_net_),
            .in3(N__39729),
            .lcout(sDAC_data_RNO_24Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_24_2_LC_15_18_6.C_ON=1'b0;
    defparam sDAC_mem_24_2_LC_15_18_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_2_LC_15_18_6.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_24_2_LC_15_18_6 (
            .in0(_gnd_net_),
            .in1(N__50301),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_24Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47801),
            .ce(N__39972),
            .sr(N__52984));
    defparam sDAC_data_RNO_25_6_LC_15_18_7.C_ON=1'b0;
    defparam sDAC_data_RNO_25_6_LC_15_18_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_6_LC_15_18_7.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_25_6_LC_15_18_7 (
            .in0(N__45735),
            .in1(N__45522),
            .in2(N__38673),
            .in3(N__38631),
            .lcout(sDAC_data_2_39_ns_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_7_LC_15_19_1.C_ON=1'b0;
    defparam sDAC_data_RNO_23_7_LC_15_19_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_7_LC_15_19_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_7_LC_15_19_1 (
            .in0(N__51502),
            .in1(N__38658),
            .in2(_gnd_net_),
            .in3(N__41523),
            .lcout(sDAC_data_RNO_23Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_32_6_LC_15_19_4.C_ON=1'b0;
    defparam sDAC_data_RNO_32_6_LC_15_19_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_32_6_LC_15_19_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_32_6_LC_15_19_4 (
            .in0(N__51478),
            .in1(N__41241),
            .in2(_gnd_net_),
            .in3(N__38640),
            .lcout(sDAC_data_RNO_32Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_31_3_LC_15_19_5.C_ON=1'b0;
    defparam sDAC_data_RNO_31_3_LC_15_19_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_3_LC_15_19_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_31_3_LC_15_19_5 (
            .in0(N__38625),
            .in1(N__51477),
            .in2(_gnd_net_),
            .in3(N__40113),
            .lcout(sDAC_data_RNO_31Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_29_6_LC_15_19_6.C_ON=1'b0;
    defparam sDAC_data_RNO_29_6_LC_15_19_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_6_LC_15_19_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_29_6_LC_15_19_6 (
            .in0(N__51479),
            .in1(N__38610),
            .in2(_gnd_net_),
            .in3(N__44055),
            .lcout(sDAC_data_RNO_29Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ00Q2_0_LC_16_2_3 .C_ON=1'b0;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ00Q2_0_LC_16_2_3 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ00Q2_0_LC_16_2_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \spi_slave_inst.tx_data_count_neg_sclk_i_RNIQ00Q2_0_LC_16_2_3  (
            .in0(N__38595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38563),
            .lcout(spi_miso_ft_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_8_3_LC_16_3_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_8_3_LC_16_3_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_8_3_LC_16_3_0.LUT_INIT=16'b0000010000000000;
    LogicCell40 sAddress_RNI9IH12_8_3_LC_16_3_0 (
            .in0(N__40613),
            .in1(N__40641),
            .in2(N__46452),
            .in3(N__40417),
            .lcout(sDAC_mem_34_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_36_0_LC_16_4_0.C_ON=1'b0;
    defparam sDAC_mem_36_0_LC_16_4_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_0_LC_16_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_0_LC_16_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51082),
            .lcout(sDAC_mem_36Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47787),
            .ce(N__40656),
            .sr(N__53127));
    defparam sDAC_mem_36_1_LC_16_4_1.C_ON=1'b0;
    defparam sDAC_mem_36_1_LC_16_4_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_1_LC_16_4_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_1_LC_16_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50677),
            .lcout(sDAC_mem_36Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47787),
            .ce(N__40656),
            .sr(N__53127));
    defparam sDAC_mem_36_2_LC_16_4_2.C_ON=1'b0;
    defparam sDAC_mem_36_2_LC_16_4_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_2_LC_16_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_2_LC_16_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50151),
            .lcout(sDAC_mem_36Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47787),
            .ce(N__40656),
            .sr(N__53127));
    defparam sDAC_mem_36_3_LC_16_4_3.C_ON=1'b0;
    defparam sDAC_mem_36_3_LC_16_4_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_3_LC_16_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_3_LC_16_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49661),
            .lcout(sDAC_mem_36Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47787),
            .ce(N__40656),
            .sr(N__53127));
    defparam sDAC_mem_36_4_LC_16_4_4.C_ON=1'b0;
    defparam sDAC_mem_36_4_LC_16_4_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_4_LC_16_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_4_LC_16_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49109),
            .lcout(sDAC_mem_36Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47787),
            .ce(N__40656),
            .sr(N__53127));
    defparam sDAC_mem_36_5_LC_16_4_5.C_ON=1'b0;
    defparam sDAC_mem_36_5_LC_16_4_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_5_LC_16_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_5_LC_16_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46877),
            .lcout(sDAC_mem_36Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47787),
            .ce(N__40656),
            .sr(N__53127));
    defparam sDAC_mem_36_6_LC_16_4_6.C_ON=1'b0;
    defparam sDAC_mem_36_6_LC_16_4_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_6_LC_16_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_6_LC_16_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48190),
            .lcout(sDAC_mem_36Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47787),
            .ce(N__40656),
            .sr(N__53127));
    defparam sDAC_mem_36_7_LC_16_4_7.C_ON=1'b0;
    defparam sDAC_mem_36_7_LC_16_4_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_36_7_LC_16_4_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_36_7_LC_16_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48737),
            .lcout(sDAC_mem_36Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47787),
            .ce(N__40656),
            .sr(N__53127));
    defparam sDAC_mem_37_0_LC_16_5_0.C_ON=1'b0;
    defparam sDAC_mem_37_0_LC_16_5_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_0_LC_16_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_0_LC_16_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51100),
            .lcout(sDAC_mem_37Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47771),
            .ce(N__40149),
            .sr(N__53112));
    defparam sDAC_mem_37_1_LC_16_5_1.C_ON=1'b0;
    defparam sDAC_mem_37_1_LC_16_5_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_1_LC_16_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_1_LC_16_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50686),
            .lcout(sDAC_mem_37Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47771),
            .ce(N__40149),
            .sr(N__53112));
    defparam sDAC_mem_37_2_LC_16_5_2.C_ON=1'b0;
    defparam sDAC_mem_37_2_LC_16_5_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_2_LC_16_5_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_37_2_LC_16_5_2 (
            .in0(N__50240),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_37Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47771),
            .ce(N__40149),
            .sr(N__53112));
    defparam sDAC_mem_37_3_LC_16_5_3.C_ON=1'b0;
    defparam sDAC_mem_37_3_LC_16_5_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_3_LC_16_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_3_LC_16_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49765),
            .lcout(sDAC_mem_37Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47771),
            .ce(N__40149),
            .sr(N__53112));
    defparam sDAC_mem_37_4_LC_16_5_4.C_ON=1'b0;
    defparam sDAC_mem_37_4_LC_16_5_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_4_LC_16_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_4_LC_16_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49110),
            .lcout(sDAC_mem_37Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47771),
            .ce(N__40149),
            .sr(N__53112));
    defparam sDAC_mem_37_5_LC_16_5_5.C_ON=1'b0;
    defparam sDAC_mem_37_5_LC_16_5_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_5_LC_16_5_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_37_5_LC_16_5_5 (
            .in0(N__46879),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_37Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47771),
            .ce(N__40149),
            .sr(N__53112));
    defparam sDAC_mem_37_6_LC_16_5_6.C_ON=1'b0;
    defparam sDAC_mem_37_6_LC_16_5_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_6_LC_16_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_6_LC_16_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48192),
            .lcout(sDAC_mem_37Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47771),
            .ce(N__40149),
            .sr(N__53112));
    defparam sDAC_mem_37_7_LC_16_5_7.C_ON=1'b0;
    defparam sDAC_mem_37_7_LC_16_5_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_37_7_LC_16_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_37_7_LC_16_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48738),
            .lcout(sDAC_mem_37Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47771),
            .ce(N__40149),
            .sr(N__53112));
    defparam sDAC_mem_8_0_LC_16_6_0.C_ON=1'b0;
    defparam sDAC_mem_8_0_LC_16_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_0_LC_16_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_0_LC_16_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51101),
            .lcout(sDAC_mem_8Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47760),
            .ce(N__38796),
            .sr(N__53100));
    defparam sDAC_mem_8_1_LC_16_6_1.C_ON=1'b0;
    defparam sDAC_mem_8_1_LC_16_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_1_LC_16_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_1_LC_16_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50687),
            .lcout(sDAC_mem_8Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47760),
            .ce(N__38796),
            .sr(N__53100));
    defparam sDAC_mem_8_2_LC_16_6_2.C_ON=1'b0;
    defparam sDAC_mem_8_2_LC_16_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_2_LC_16_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_2_LC_16_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50241),
            .lcout(sDAC_mem_8Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47760),
            .ce(N__38796),
            .sr(N__53100));
    defparam sDAC_mem_8_3_LC_16_6_3.C_ON=1'b0;
    defparam sDAC_mem_8_3_LC_16_6_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_3_LC_16_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_3_LC_16_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49766),
            .lcout(sDAC_mem_8Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47760),
            .ce(N__38796),
            .sr(N__53100));
    defparam sDAC_mem_8_4_LC_16_6_4.C_ON=1'b0;
    defparam sDAC_mem_8_4_LC_16_6_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_4_LC_16_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_4_LC_16_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49358),
            .lcout(sDAC_mem_8Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47760),
            .ce(N__38796),
            .sr(N__53100));
    defparam sDAC_mem_8_5_LC_16_6_5.C_ON=1'b0;
    defparam sDAC_mem_8_5_LC_16_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_5_LC_16_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_5_LC_16_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46880),
            .lcout(sDAC_mem_8Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47760),
            .ce(N__38796),
            .sr(N__53100));
    defparam sDAC_mem_8_6_LC_16_6_6.C_ON=1'b0;
    defparam sDAC_mem_8_6_LC_16_6_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_6_LC_16_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_6_LC_16_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48211),
            .lcout(sDAC_mem_8Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47760),
            .ce(N__38796),
            .sr(N__53100));
    defparam sDAC_mem_8_7_LC_16_6_7.C_ON=1'b0;
    defparam sDAC_mem_8_7_LC_16_6_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_8_7_LC_16_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_8_7_LC_16_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48740),
            .lcout(sDAC_mem_8Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47760),
            .ce(N__38796),
            .sr(N__53100));
    defparam sDAC_data_RNO_20_7_LC_16_7_0.C_ON=1'b0;
    defparam sDAC_data_RNO_20_7_LC_16_7_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_7_LC_16_7_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_20_7_LC_16_7_0 (
            .in0(N__52002),
            .in1(N__40704),
            .in2(_gnd_net_),
            .in3(N__38781),
            .lcout(sDAC_data_RNO_20Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_20_4_LC_16_7_1.C_ON=1'b0;
    defparam sDAC_mem_20_4_LC_16_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_4_LC_16_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_4_LC_16_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49111),
            .lcout(sDAC_mem_20Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47748),
            .ce(N__44029),
            .sr(N__53086));
    defparam sDAC_data_RNO_20_8_LC_16_7_2.C_ON=1'b0;
    defparam sDAC_data_RNO_20_8_LC_16_7_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_8_LC_16_7_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_20_8_LC_16_7_2 (
            .in0(N__40698),
            .in1(N__51999),
            .in2(_gnd_net_),
            .in3(N__38775),
            .lcout(sDAC_data_RNO_20Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_20_5_LC_16_7_3.C_ON=1'b0;
    defparam sDAC_mem_20_5_LC_16_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_5_LC_16_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_5_LC_16_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46881),
            .lcout(sDAC_mem_20Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47748),
            .ce(N__44029),
            .sr(N__53086));
    defparam sDAC_data_RNO_20_9_LC_16_7_4.C_ON=1'b0;
    defparam sDAC_data_RNO_20_9_LC_16_7_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_9_LC_16_7_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_20_9_LC_16_7_4 (
            .in0(N__52001),
            .in1(N__40692),
            .in2(_gnd_net_),
            .in3(N__38961),
            .lcout(sDAC_data_RNO_20Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_20_6_LC_16_7_5.C_ON=1'b0;
    defparam sDAC_mem_20_6_LC_16_7_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_6_LC_16_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_6_LC_16_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48212),
            .lcout(sDAC_mem_20Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47748),
            .ce(N__44029),
            .sr(N__53086));
    defparam sDAC_data_RNO_21_10_LC_16_7_6.C_ON=1'b0;
    defparam sDAC_data_RNO_21_10_LC_16_7_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_10_LC_16_7_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_10_LC_16_7_6 (
            .in0(N__52000),
            .in1(N__38955),
            .in2(_gnd_net_),
            .in3(N__38946),
            .lcout(sDAC_data_RNO_21Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_21_3_LC_16_7_7.C_ON=1'b0;
    defparam sDAC_data_RNO_21_3_LC_16_7_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_3_LC_16_7_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_3_LC_16_7_7 (
            .in0(N__51998),
            .in1(N__38931),
            .in2(_gnd_net_),
            .in3(N__38922),
            .lcout(sDAC_data_RNO_21Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_13_7_LC_16_8_1.C_ON=1'b0;
    defparam sDAC_data_RNO_13_7_LC_16_8_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_7_LC_16_8_1.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_13_7_LC_16_8_1 (
            .in0(N__52122),
            .in1(N__41625),
            .in2(N__43669),
            .in3(N__40824),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_7_LC_16_8_2.C_ON=1'b0;
    defparam sDAC_data_RNO_5_7_LC_16_8_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_7_LC_16_8_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_5_7_LC_16_8_2 (
            .in0(N__51811),
            .in1(N__40173),
            .in2(N__38907),
            .in3(N__38904),
            .lcout(sDAC_data_RNO_5Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_7_LC_16_8_3.C_ON=1'b0;
    defparam sDAC_data_RNO_22_7_LC_16_8_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_7_LC_16_8_3.LUT_INIT=16'b0100011001010111;
    LogicCell40 sDAC_data_RNO_22_7_LC_16_8_3 (
            .in0(N__45490),
            .in1(N__45799),
            .in2(N__38886),
            .in3(N__38868),
            .lcout(sDAC_data_2_32_ns_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_7_3_LC_16_8_5.C_ON=1'b0;
    defparam sAddress_RNI9IH12_7_3_LC_16_8_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_7_3_LC_16_8_5.LUT_INIT=16'b0000100000000000;
    LogicCell40 sAddress_RNI9IH12_7_3_LC_16_8_5 (
            .in0(N__40416),
            .in1(N__43281),
            .in2(N__40603),
            .in3(N__43190),
            .lcout(sDAC_mem_20_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_28_7_LC_16_8_6.C_ON=1'b0;
    defparam sDAC_data_RNO_28_7_LC_16_8_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_7_LC_16_8_6.LUT_INIT=16'b0010011000110111;
    LogicCell40 sDAC_data_RNO_28_7_LC_16_8_6 (
            .in0(N__51809),
            .in1(N__43624),
            .in2(N__38856),
            .in3(N__38841),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_7_LC_16_8_7.C_ON=1'b0;
    defparam sDAC_data_RNO_15_7_LC_16_8_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_7_LC_16_8_7.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_15_7_LC_16_8_7 (
            .in0(N__39081),
            .in1(N__51810),
            .in2(N__39075),
            .in3(N__40209),
            .lcout(sDAC_data_RNO_15Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_12_8_LC_16_9_0.C_ON=1'b0;
    defparam sDAC_data_RNO_12_8_LC_16_9_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_8_LC_16_9_0.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_12_8_LC_16_9_0 (
            .in0(N__52116),
            .in1(N__39066),
            .in2(N__43565),
            .in3(N__39033),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_8_LC_16_9_1.C_ON=1'b0;
    defparam sDAC_data_RNO_4_8_LC_16_9_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_8_LC_16_9_1.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_8_LC_16_9_1 (
            .in0(N__52105),
            .in1(N__39057),
            .in2(N__39048),
            .in3(N__39045),
            .lcout(sDAC_data_RNO_4Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_4_5_LC_16_9_2.C_ON=1'b0;
    defparam sDAC_mem_4_5_LC_16_9_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_5_LC_16_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_5_LC_16_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47088),
            .lcout(sDAC_mem_4Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47725),
            .ce(N__39631),
            .sr(N__53063));
    defparam sDAC_data_RNO_12_9_LC_16_9_3.C_ON=1'b0;
    defparam sDAC_data_RNO_12_9_LC_16_9_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_9_LC_16_9_3.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_12_9_LC_16_9_3 (
            .in0(N__52106),
            .in1(N__39027),
            .in2(N__43686),
            .in3(N__38994),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_9_LC_16_9_4.C_ON=1'b0;
    defparam sDAC_data_RNO_4_9_LC_16_9_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_9_LC_16_9_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_9_LC_16_9_4 (
            .in0(N__52117),
            .in1(N__39018),
            .in2(N__39009),
            .in3(N__39006),
            .lcout(sDAC_data_RNO_4Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_4_6_LC_16_9_5.C_ON=1'b0;
    defparam sDAC_mem_4_6_LC_16_9_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_6_LC_16_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_6_LC_16_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48235),
            .lcout(sDAC_mem_4Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47725),
            .ce(N__39631),
            .sr(N__53063));
    defparam sDAC_data_RNO_13_10_LC_16_9_6.C_ON=1'b0;
    defparam sDAC_data_RNO_13_10_LC_16_9_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_10_LC_16_9_6.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_13_10_LC_16_9_6 (
            .in0(N__52115),
            .in1(N__41880),
            .in2(N__43564),
            .in3(N__38988),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_10_LC_16_9_7.C_ON=1'b0;
    defparam sDAC_data_RNO_5_10_LC_16_9_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_10_LC_16_9_7.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_5_10_LC_16_9_7 (
            .in0(N__52104),
            .in1(N__40161),
            .in2(N__38976),
            .in3(N__38973),
            .lcout(sDAC_data_RNO_5Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_9_LC_16_10_0.C_ON=1'b0;
    defparam sDAC_data_RNO_1_9_LC_16_10_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_9_LC_16_10_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_1_9_LC_16_10_0 (
            .in0(N__42726),
            .in1(N__39195),
            .in2(N__45808),
            .in3(N__39132),
            .lcout(),
            .ltout(sDAC_data_RNO_1Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_9_LC_16_10_1.C_ON=1'b0;
    defparam sDAC_data_RNO_0_9_LC_16_10_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_9_LC_16_10_1.LUT_INIT=16'b0101000011101110;
    LogicCell40 sDAC_data_RNO_0_9_LC_16_10_1 (
            .in0(N__42517),
            .in1(N__39189),
            .in2(N__39177),
            .in3(N__39087),
            .lcout(),
            .ltout(sDAC_data_2_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_9_LC_16_10_2.C_ON=1'b0;
    defparam sDAC_data_9_LC_16_10_2.SEQ_MODE=4'b1010;
    defparam sDAC_data_9_LC_16_10_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 sDAC_data_9_LC_16_10_2 (
            .in0(_gnd_net_),
            .in1(N__47250),
            .in2(N__39174),
            .in3(N__42380),
            .lcout(sDAC_dataZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53257),
            .ce(N__42222),
            .sr(N__53053));
    defparam sDAC_data_RNO_6_9_LC_16_10_3.C_ON=1'b0;
    defparam sDAC_data_RNO_6_9_LC_16_10_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_9_LC_16_10_3.LUT_INIT=16'b0100011001010111;
    LogicCell40 sDAC_data_RNO_6_9_LC_16_10_3 (
            .in0(N__45533),
            .in1(N__45712),
            .in2(N__39156),
            .in3(N__39144),
            .lcout(sDAC_data_2_14_ns_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_9_LC_16_10_4.C_ON=1'b0;
    defparam sDAC_data_RNO_22_9_LC_16_10_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_9_LC_16_10_4.LUT_INIT=16'b0000101101011011;
    LogicCell40 sDAC_data_RNO_22_9_LC_16_10_4 (
            .in0(N__45711),
            .in1(N__39126),
            .in2(N__45534),
            .in3(N__39120),
            .lcout(),
            .ltout(sDAC_data_2_32_ns_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_9_LC_16_10_5.C_ON=1'b0;
    defparam sDAC_data_RNO_10_9_LC_16_10_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_9_LC_16_10_5.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_10_9_LC_16_10_5 (
            .in0(N__45716),
            .in1(N__39843),
            .in2(N__39108),
            .in3(N__39105),
            .lcout(),
            .ltout(sDAC_data_RNO_10Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_9_LC_16_10_6.C_ON=1'b0;
    defparam sDAC_data_RNO_3_9_LC_16_10_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_9_LC_16_10_6.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_3_9_LC_16_10_6 (
            .in0(N__42479),
            .in1(N__42610),
            .in2(N__39096),
            .in3(N__39093),
            .lcout(sDAC_data_2_41_ns_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_3_5_LC_16_11_0.C_ON=1'b0;
    defparam sDAC_mem_3_5_LC_16_11_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_5_LC_16_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_3_5_LC_16_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47089),
            .lcout(sDAC_mem_3Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47713),
            .ce(N__42984),
            .sr(N__53043));
    defparam sDAC_data_RNO_28_8_LC_16_11_1.C_ON=1'b0;
    defparam sDAC_data_RNO_28_8_LC_16_11_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_8_LC_16_11_1.LUT_INIT=16'b0100010101100111;
    LogicCell40 sDAC_data_RNO_28_8_LC_16_11_1 (
            .in0(N__43450),
            .in1(N__52092),
            .in2(N__39399),
            .in3(N__39384),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_8_LC_16_11_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_8_LC_16_11_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_8_LC_16_11_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_8_LC_16_11_2 (
            .in0(N__52093),
            .in1(N__40194),
            .in2(N__39369),
            .in3(N__39366),
            .lcout(sDAC_data_RNO_15Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_26_10_LC_16_11_3.C_ON=1'b0;
    defparam sDAC_data_RNO_26_10_LC_16_11_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_10_LC_16_11_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 sDAC_data_RNO_26_10_LC_16_11_3 (
            .in0(N__43449),
            .in1(N__52094),
            .in2(N__39342),
            .in3(N__39320),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_10_LC_16_11_4.C_ON=1'b0;
    defparam sDAC_data_RNO_14_10_LC_16_11_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_10_LC_16_11_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_14_10_LC_16_11_4 (
            .in0(_gnd_net_),
            .in1(N__39360),
            .in2(N__39345),
            .in3(N__39306),
            .lcout(sDAC_data_RNO_14Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_27_10_LC_16_11_5.C_ON=1'b0;
    defparam sDAC_data_RNO_27_10_LC_16_11_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_10_LC_16_11_5.LUT_INIT=16'b1111101111001000;
    LogicCell40 sDAC_data_RNO_27_10_LC_16_11_5 (
            .in0(N__43448),
            .in1(N__52091),
            .in2(N__39341),
            .in3(N__39321),
            .lcout(sDAC_data_RNO_27Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_26_3_LC_16_11_6.C_ON=1'b0;
    defparam sDAC_data_RNO_26_3_LC_16_11_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_3_LC_16_11_6.LUT_INIT=16'b0111010100100000;
    LogicCell40 sDAC_data_RNO_26_3_LC_16_11_6 (
            .in0(N__52095),
            .in1(N__43451),
            .in2(N__39300),
            .in3(N__39270),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_3_LC_16_11_7.C_ON=1'b0;
    defparam sDAC_data_RNO_14_3_LC_16_11_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_3_LC_16_11_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_14_3_LC_16_11_7 (
            .in0(_gnd_net_),
            .in1(N__39252),
            .in2(N__39237),
            .in3(N__39234),
            .lcout(sDAC_data_RNO_14Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_10_LC_16_12_0.C_ON=1'b0;
    defparam sDAC_data_RNO_10_10_LC_16_12_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_10_LC_16_12_0.LUT_INIT=16'b1010000011001111;
    LogicCell40 sDAC_data_RNO_10_10_LC_16_12_0 (
            .in0(N__39537),
            .in1(N__39225),
            .in2(N__45882),
            .in3(N__39201),
            .lcout(sDAC_data_RNO_10Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_10_LC_16_12_1.C_ON=1'b0;
    defparam sDAC_data_RNO_22_10_LC_16_12_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_10_LC_16_12_1.LUT_INIT=16'b0010011000110111;
    LogicCell40 sDAC_data_RNO_22_10_LC_16_12_1 (
            .in0(N__45728),
            .in1(N__45423),
            .in2(N__39213),
            .in3(N__41322),
            .lcout(sDAC_data_2_32_ns_1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_10_LC_16_12_2.C_ON=1'b0;
    defparam sDAC_data_RNO_6_10_LC_16_12_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_10_LC_16_12_2.LUT_INIT=16'b0000001111011101;
    LogicCell40 sDAC_data_RNO_6_10_LC_16_12_2 (
            .in0(N__39513),
            .in1(N__45729),
            .in2(N__42849),
            .in3(N__45523),
            .lcout(),
            .ltout(sDAC_data_2_14_ns_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_10_LC_16_12_3.C_ON=1'b0;
    defparam sDAC_data_RNO_1_10_LC_16_12_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_10_LC_16_12_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_1_10_LC_16_12_3 (
            .in0(N__45730),
            .in1(N__39504),
            .in2(N__39495),
            .in3(N__39411),
            .lcout(sDAC_data_RNO_1Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_10_LC_16_12_4.C_ON=1'b0;
    defparam sDAC_data_RNO_3_10_LC_16_12_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_10_LC_16_12_4.LUT_INIT=16'b0000101001110111;
    LogicCell40 sDAC_data_RNO_3_10_LC_16_12_4 (
            .in0(N__42532),
            .in1(N__39492),
            .in2(N__40044),
            .in3(N__42630),
            .lcout(),
            .ltout(sDAC_data_2_41_ns_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_10_LC_16_12_5.C_ON=1'b0;
    defparam sDAC_data_RNO_0_10_LC_16_12_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_10_LC_16_12_5.LUT_INIT=16'b0101111000001110;
    LogicCell40 sDAC_data_RNO_0_10_LC_16_12_5 (
            .in0(N__42533),
            .in1(N__39486),
            .in2(N__39480),
            .in3(N__39477),
            .lcout(),
            .ltout(sDAC_data_2_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_10_LC_16_12_6.C_ON=1'b0;
    defparam sDAC_data_10_LC_16_12_6.SEQ_MODE=4'b1010;
    defparam sDAC_data_10_LC_16_12_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 sDAC_data_10_LC_16_12_6 (
            .in0(_gnd_net_),
            .in1(N__46587),
            .in2(N__39471),
            .in3(N__42378),
            .lcout(sDAC_dataZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53268),
            .ce(N__42227),
            .sr(N__53034));
    defparam sDAC_data_RNO_12_10_LC_16_13_0.C_ON=1'b0;
    defparam sDAC_data_RNO_12_10_LC_16_13_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_10_LC_16_13_0.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_12_10_LC_16_13_0 (
            .in0(N__51971),
            .in1(N__39450),
            .in2(N__43634),
            .in3(N__39405),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_10_LC_16_13_1.C_ON=1'b0;
    defparam sDAC_data_RNO_4_10_LC_16_13_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_10_LC_16_13_1.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_10_LC_16_13_1 (
            .in0(N__51996),
            .in1(N__39438),
            .in2(N__39426),
            .in3(N__39423),
            .lcout(sDAC_data_RNO_4Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_4_7_LC_16_13_2.C_ON=1'b0;
    defparam sDAC_mem_4_7_LC_16_13_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_7_LC_16_13_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_4_7_LC_16_13_2 (
            .in0(N__48834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_4Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47726),
            .ce(N__39639),
            .sr(N__53024));
    defparam sDAC_data_RNO_12_3_LC_16_13_3.C_ON=1'b0;
    defparam sDAC_data_RNO_12_3_LC_16_13_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_3_LC_16_13_3.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_12_3_LC_16_13_3 (
            .in0(N__51997),
            .in1(N__39687),
            .in2(N__43635),
            .in3(N__39645),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_3_LC_16_13_4.C_ON=1'b0;
    defparam sDAC_data_RNO_4_3_LC_16_13_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_3_LC_16_13_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_3_LC_16_13_4 (
            .in0(N__51972),
            .in1(N__39675),
            .in2(N__39660),
            .in3(N__39657),
            .lcout(sDAC_data_RNO_4Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_4_0_LC_16_13_5.C_ON=1'b0;
    defparam sDAC_mem_4_0_LC_16_13_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_4_0_LC_16_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_4_0_LC_16_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51252),
            .lcout(sDAC_mem_4Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47726),
            .ce(N__39639),
            .sr(N__53024));
    defparam sDAC_data_RNO_12_4_LC_16_13_6.C_ON=1'b0;
    defparam sDAC_data_RNO_12_4_LC_16_13_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_12_4_LC_16_13_6.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_12_4_LC_16_13_6 (
            .in0(N__51970),
            .in1(N__39597),
            .in2(N__43633),
            .in3(N__39588),
            .lcout(),
            .ltout(sDAC_data_2_13_am_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_4_4_LC_16_13_7.C_ON=1'b0;
    defparam sDAC_data_RNO_4_4_LC_16_13_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_4_4_LC_16_13_7.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_4_4_LC_16_13_7 (
            .in0(N__51995),
            .in1(N__39570),
            .in2(N__39555),
            .in3(N__39552),
            .lcout(sDAC_data_RNO_4Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_20_10_LC_16_14_0.C_ON=1'b0;
    defparam sDAC_data_RNO_20_10_LC_16_14_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_10_LC_16_14_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_20_10_LC_16_14_0 (
            .in0(N__51985),
            .in1(N__40686),
            .in2(_gnd_net_),
            .in3(N__44046),
            .lcout(sDAC_data_RNO_20Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_4_1_LC_16_14_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_4_1_LC_16_14_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_4_1_LC_16_14_2.LUT_INIT=16'b0100010000000000;
    LogicCell40 sAddress_RNI9IH12_4_1_LC_16_14_2 (
            .in0(N__44410),
            .in1(N__46244),
            .in2(_gnd_net_),
            .in3(N__43179),
            .lcout(sDAC_mem_30_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_2_1_LC_16_14_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_2_1_LC_16_14_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_2_1_LC_16_14_3.LUT_INIT=16'b0010001000000000;
    LogicCell40 sAddress_RNI9IH12_2_1_LC_16_14_3 (
            .in0(N__43178),
            .in1(N__44409),
            .in2(_gnd_net_),
            .in3(N__43254),
            .lcout(sDAC_mem_28_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_0_1_LC_16_14_4.C_ON=1'b0;
    defparam sAddress_RNI9IH12_0_1_LC_16_14_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_0_1_LC_16_14_4.LUT_INIT=16'b0001000100000000;
    LogicCell40 sAddress_RNI9IH12_0_1_LC_16_14_4 (
            .in0(N__44411),
            .in1(N__46418),
            .in2(_gnd_net_),
            .in3(N__43177),
            .lcout(sDAC_mem_26_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI5B15_0_3_LC_16_14_5.C_ON=1'b0;
    defparam sAddress_RNI5B15_0_3_LC_16_14_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNI5B15_0_3_LC_16_14_5.LUT_INIT=16'b0011001111111111;
    LogicCell40 sAddress_RNI5B15_0_3_LC_16_14_5 (
            .in0(_gnd_net_),
            .in1(N__40541),
            .in2(_gnd_net_),
            .in3(N__40359),
            .lcout(N_142),
            .ltout(N_142_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_rpi_ibuf_RNIRGF52_LC_16_14_6.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNIRGF52_LC_16_14_6.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNIRGF52_LC_16_14_6.LUT_INIT=16'b0000110000000000;
    LogicCell40 reset_rpi_ibuf_RNIRGF52_LC_16_14_6 (
            .in0(_gnd_net_),
            .in1(N__46243),
            .in2(N__39732),
            .in3(N__46044),
            .lcout(sEEADC_freq_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_30_0_LC_16_15_0.C_ON=1'b0;
    defparam sDAC_mem_30_0_LC_16_15_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_0_LC_16_15_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_0_LC_16_15_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51248),
            .lcout(sDAC_mem_30Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47749),
            .ce(N__39693),
            .sr(N__53013));
    defparam sDAC_mem_30_1_LC_16_15_1.C_ON=1'b0;
    defparam sDAC_mem_30_1_LC_16_15_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_1_LC_16_15_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_1_LC_16_15_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50724),
            .lcout(sDAC_mem_30Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47749),
            .ce(N__39693),
            .sr(N__53013));
    defparam sDAC_mem_30_2_LC_16_15_2.C_ON=1'b0;
    defparam sDAC_mem_30_2_LC_16_15_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_2_LC_16_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_2_LC_16_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50178),
            .lcout(sDAC_mem_30Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47749),
            .ce(N__39693),
            .sr(N__53013));
    defparam sDAC_mem_30_3_LC_16_15_3.C_ON=1'b0;
    defparam sDAC_mem_30_3_LC_16_15_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_3_LC_16_15_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_3_LC_16_15_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49836),
            .lcout(sDAC_mem_30Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47749),
            .ce(N__39693),
            .sr(N__53013));
    defparam sDAC_mem_30_4_LC_16_15_4.C_ON=1'b0;
    defparam sDAC_mem_30_4_LC_16_15_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_4_LC_16_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_4_LC_16_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49091),
            .lcout(sDAC_mem_30Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47749),
            .ce(N__39693),
            .sr(N__53013));
    defparam sDAC_mem_30_5_LC_16_15_5.C_ON=1'b0;
    defparam sDAC_mem_30_5_LC_16_15_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_5_LC_16_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_5_LC_16_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47135),
            .lcout(sDAC_mem_30Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47749),
            .ce(N__39693),
            .sr(N__53013));
    defparam sDAC_mem_30_6_LC_16_15_6.C_ON=1'b0;
    defparam sDAC_mem_30_6_LC_16_15_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_6_LC_16_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_6_LC_16_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48338),
            .lcout(sDAC_mem_30Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47749),
            .ce(N__39693),
            .sr(N__53013));
    defparam sDAC_mem_30_7_LC_16_15_7.C_ON=1'b0;
    defparam sDAC_mem_30_7_LC_16_15_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_30_7_LC_16_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_30_7_LC_16_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48831),
            .lcout(sDAC_mem_30Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47749),
            .ce(N__39693),
            .sr(N__53013));
    defparam sDAC_data_RNO_21_8_LC_16_16_0.C_ON=1'b0;
    defparam sDAC_data_RNO_21_8_LC_16_16_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_8_LC_16_16_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_8_LC_16_16_0 (
            .in0(N__51888),
            .in1(N__39885),
            .in2(_gnd_net_),
            .in3(N__39867),
            .lcout(sDAC_data_RNO_21Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_22_5_LC_16_16_1.C_ON=1'b0;
    defparam sDAC_mem_22_5_LC_16_16_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_5_LC_16_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_5_LC_16_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47136),
            .lcout(sDAC_mem_22Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47761),
            .ce(N__39825),
            .sr(N__53004));
    defparam sDAC_data_RNO_21_9_LC_16_16_2.C_ON=1'b0;
    defparam sDAC_data_RNO_21_9_LC_16_16_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_9_LC_16_16_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_9_LC_16_16_2 (
            .in0(N__51889),
            .in1(N__39861),
            .in2(_gnd_net_),
            .in3(N__39831),
            .lcout(sDAC_data_RNO_21Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_22_6_LC_16_16_3.C_ON=1'b0;
    defparam sDAC_mem_22_6_LC_16_16_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_22_6_LC_16_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_22_6_LC_16_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48339),
            .lcout(sDAC_mem_22Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47761),
            .ce(N__39825),
            .sr(N__53004));
    defparam sDAC_data_RNO_23_4_LC_16_16_4.C_ON=1'b0;
    defparam sDAC_data_RNO_23_4_LC_16_16_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_4_LC_16_16_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_23_4_LC_16_16_4 (
            .in0(N__39786),
            .in1(N__51886),
            .in2(_gnd_net_),
            .in3(N__41541),
            .lcout(sDAC_data_RNO_23Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_4_LC_16_16_6.C_ON=1'b0;
    defparam sDAC_data_RNO_24_4_LC_16_16_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_4_LC_16_16_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_24_4_LC_16_16_6 (
            .in0(N__51887),
            .in1(N__39780),
            .in2(_gnd_net_),
            .in3(N__39774),
            .lcout(sDAC_data_RNO_24Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_7_LC_16_16_7.C_ON=1'b0;
    defparam sDAC_data_RNO_24_7_LC_16_16_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_7_LC_16_16_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_7_LC_16_16_7 (
            .in0(N__51885),
            .in1(N__39762),
            .in2(_gnd_net_),
            .in3(N__39750),
            .lcout(sDAC_data_RNO_24Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_31_10_LC_16_17_0.C_ON=1'b0;
    defparam sDAC_data_RNO_31_10_LC_16_17_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_10_LC_16_17_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_31_10_LC_16_17_0 (
            .in0(N__51895),
            .in1(N__39978),
            .in2(_gnd_net_),
            .in3(N__39891),
            .lcout(),
            .ltout(sDAC_data_RNO_31Z0Z_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_25_10_LC_16_17_1.C_ON=1'b0;
    defparam sDAC_data_RNO_25_10_LC_16_17_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_10_LC_16_17_1.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_25_10_LC_16_17_1 (
            .in0(N__45877),
            .in1(N__45481),
            .in2(N__39735),
            .in3(N__40023),
            .lcout(),
            .ltout(sDAC_data_2_39_ns_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_10_LC_16_17_2.C_ON=1'b0;
    defparam sDAC_data_RNO_11_10_LC_16_17_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_10_LC_16_17_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_11_10_LC_16_17_2 (
            .in0(N__45878),
            .in1(N__39984),
            .in2(N__40047),
            .in3(N__40011),
            .lcout(sDAC_data_RNO_11Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_32_10_LC_16_17_3.C_ON=1'b0;
    defparam sDAC_data_RNO_32_10_LC_16_17_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_32_10_LC_16_17_3.LUT_INIT=16'b1111001111000000;
    LogicCell40 sDAC_data_RNO_32_10_LC_16_17_3 (
            .in0(_gnd_net_),
            .in1(N__51893),
            .in2(N__41472),
            .in3(N__40032),
            .lcout(sDAC_data_RNO_32Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_10_LC_16_17_4.C_ON=1'b0;
    defparam sDAC_data_RNO_23_10_LC_16_17_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_10_LC_16_17_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_10_LC_16_17_4 (
            .in0(N__51894),
            .in1(N__40017),
            .in2(_gnd_net_),
            .in3(N__41784),
            .lcout(sDAC_data_RNO_23Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_10_LC_16_17_5.C_ON=1'b0;
    defparam sDAC_data_RNO_24_10_LC_16_17_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_10_LC_16_17_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_10_LC_16_17_5 (
            .in0(N__51896),
            .in1(N__40005),
            .in2(_gnd_net_),
            .in3(N__39993),
            .lcout(sDAC_data_RNO_24Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_24_7_LC_16_17_6.C_ON=1'b0;
    defparam sDAC_mem_24_7_LC_16_17_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_24_7_LC_16_17_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_24_7_LC_16_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48799),
            .lcout(sDAC_mem_24Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47772),
            .ce(N__39967),
            .sr(N__52995));
    defparam sDAC_data_RNO_25_3_LC_16_17_7.C_ON=1'b0;
    defparam sDAC_data_RNO_25_3_LC_16_17_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_3_LC_16_17_7.LUT_INIT=16'b0010011000110111;
    LogicCell40 sDAC_data_RNO_25_3_LC_16_17_7 (
            .in0(N__45876),
            .in1(N__45480),
            .in2(N__39921),
            .in3(N__39906),
            .lcout(sDAC_data_2_39_ns_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_25_4_LC_16_18_2.C_ON=1'b0;
    defparam sDAC_mem_25_4_LC_16_18_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_4_LC_16_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_4_LC_16_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49327),
            .lcout(sDAC_mem_25Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47788),
            .ce(N__41723),
            .sr(N__52990));
    defparam sDAC_mem_25_7_LC_16_18_3.C_ON=1'b0;
    defparam sDAC_mem_25_7_LC_16_18_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_7_LC_16_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_7_LC_16_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48801),
            .lcout(sDAC_mem_25Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47788),
            .ce(N__41723),
            .sr(N__52990));
    defparam sDAC_mem_25_2_LC_16_18_4.C_ON=1'b0;
    defparam sDAC_mem_25_2_LC_16_18_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_2_LC_16_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_2_LC_16_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50299),
            .lcout(sDAC_mem_25Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47788),
            .ce(N__41723),
            .sr(N__52990));
    defparam sDAC_mem_25_5_LC_16_18_6.C_ON=1'b0;
    defparam sDAC_mem_25_5_LC_16_18_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_5_LC_16_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_5_LC_16_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47131),
            .lcout(sDAC_mem_25Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47788),
            .ce(N__41723),
            .sr(N__52990));
    defparam sDAC_mem_25_0_LC_16_19_0.C_ON=1'b0;
    defparam sDAC_mem_25_0_LC_16_19_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_0_LC_16_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_0_LC_16_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51271),
            .lcout(sDAC_mem_25Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47802),
            .ce(N__41727),
            .sr(N__52985));
    defparam sDAC_mem_25_6_LC_16_19_2.C_ON=1'b0;
    defparam sDAC_mem_25_6_LC_16_19_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_6_LC_16_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_6_LC_16_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48342),
            .lcout(sDAC_mem_25Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47802),
            .ce(N__41727),
            .sr(N__52985));
    defparam sDAC_mem_25_3_LC_16_19_5.C_ON=1'b0;
    defparam sDAC_mem_25_3_LC_16_19_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_3_LC_16_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_3_LC_16_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49833),
            .lcout(sDAC_mem_25Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47802),
            .ce(N__41727),
            .sr(N__52985));
    defparam sDAC_mem_34_1_LC_17_3_0.C_ON=1'b0;
    defparam sDAC_mem_34_1_LC_17_3_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_1_LC_17_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_1_LC_17_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50500),
            .lcout(sDAC_mem_34Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47789),
            .ce(N__40088),
            .sr(N__53138));
    defparam sDAC_mem_34_3_LC_17_3_2.C_ON=1'b0;
    defparam sDAC_mem_34_3_LC_17_3_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_34_3_LC_17_3_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_34_3_LC_17_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49626),
            .lcout(sDAC_mem_34Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47789),
            .ce(N__40088),
            .sr(N__53138));
    defparam sDAC_mem_39_0_LC_17_4_0.C_ON=1'b0;
    defparam sDAC_mem_39_0_LC_17_4_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_0_LC_17_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_39_0_LC_17_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51083),
            .lcout(sDAC_mem_39Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47773),
            .ce(N__40140),
            .sr(N__53133));
    defparam sDAC_mem_39_1_LC_17_4_1.C_ON=1'b0;
    defparam sDAC_mem_39_1_LC_17_4_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_1_LC_17_4_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_39_1_LC_17_4_1 (
            .in0(N__50678),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_39Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47773),
            .ce(N__40140),
            .sr(N__53133));
    defparam sDAC_mem_39_2_LC_17_4_2.C_ON=1'b0;
    defparam sDAC_mem_39_2_LC_17_4_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_2_LC_17_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_39_2_LC_17_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50255),
            .lcout(sDAC_mem_39Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47773),
            .ce(N__40140),
            .sr(N__53133));
    defparam sDAC_mem_39_3_LC_17_4_3.C_ON=1'b0;
    defparam sDAC_mem_39_3_LC_17_4_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_3_LC_17_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_39_3_LC_17_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49784),
            .lcout(sDAC_mem_39Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47773),
            .ce(N__40140),
            .sr(N__53133));
    defparam sDAC_mem_39_4_LC_17_4_4.C_ON=1'b0;
    defparam sDAC_mem_39_4_LC_17_4_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_4_LC_17_4_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_39_4_LC_17_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49357),
            .lcout(sDAC_mem_39Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47773),
            .ce(N__40140),
            .sr(N__53133));
    defparam sDAC_mem_39_5_LC_17_4_5.C_ON=1'b0;
    defparam sDAC_mem_39_5_LC_17_4_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_5_LC_17_4_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_39_5_LC_17_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46985),
            .lcout(sDAC_mem_39Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47773),
            .ce(N__40140),
            .sr(N__53133));
    defparam sDAC_mem_39_6_LC_17_4_6.C_ON=1'b0;
    defparam sDAC_mem_39_6_LC_17_4_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_6_LC_17_4_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_39_6_LC_17_4_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48210),
            .lcout(sDAC_mem_39Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47773),
            .ce(N__40140),
            .sr(N__53133));
    defparam sDAC_mem_39_7_LC_17_4_7.C_ON=1'b0;
    defparam sDAC_mem_39_7_LC_17_4_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_39_7_LC_17_4_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_39_7_LC_17_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48739),
            .lcout(sDAC_mem_39Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47773),
            .ce(N__40140),
            .sr(N__53133));
    defparam sAddress_RNI9IH12_0_3_LC_17_5_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_0_3_LC_17_5_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_0_3_LC_17_5_0.LUT_INIT=16'b0100000000000000;
    LogicCell40 sAddress_RNI9IH12_0_3_LC_17_5_0 (
            .in0(N__40609),
            .in1(N__40407),
            .in2(N__44593),
            .in3(N__40633),
            .lcout(sDAC_mem_40_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_13_3_LC_17_5_1.C_ON=1'b0;
    defparam sAddress_RNI9IH12_13_3_LC_17_5_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_13_3_LC_17_5_1.LUT_INIT=16'b0000000000001000;
    LogicCell40 sAddress_RNI9IH12_13_3_LC_17_5_1 (
            .in0(N__40636),
            .in1(N__46250),
            .in2(N__40418),
            .in3(N__40610),
            .lcout(sDAC_mem_37_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_12_3_LC_17_5_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_12_3_LC_17_5_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_12_3_LC_17_5_2.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNI9IH12_12_3_LC_17_5_2 (
            .in0(N__40611),
            .in1(N__40412),
            .in2(N__44594),
            .in3(N__40635),
            .lcout(sDAC_mem_39_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_11_3_LC_17_5_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_11_3_LC_17_5_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_11_3_LC_17_5_3.LUT_INIT=16'b0000001000000000;
    LogicCell40 sAddress_RNI9IH12_11_3_LC_17_5_3 (
            .in0(N__40634),
            .in1(N__40612),
            .in2(N__40419),
            .in3(N__43255),
            .lcout(sDAC_mem_35_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_3_LC_17_5_4.C_ON=1'b0;
    defparam sAddress_RNI9IH12_3_LC_17_5_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_3_LC_17_5_4.LUT_INIT=16'b0000100000000000;
    LogicCell40 sAddress_RNI9IH12_3_LC_17_5_4 (
            .in0(N__43256),
            .in1(N__40406),
            .in2(N__40614),
            .in3(N__40637),
            .lcout(sDAC_mem_36_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIVREN1_4_LC_17_5_5.C_ON=1'b0;
    defparam sAddress_RNIVREN1_4_LC_17_5_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNIVREN1_4_LC_17_5_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 sAddress_RNIVREN1_4_LC_17_5_5 (
            .in0(N__46573),
            .in1(N__44649),
            .in2(N__44807),
            .in3(N__44750),
            .lcout(N_288),
            .ltout(N_288_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_1_3_LC_17_5_6.C_ON=1'b0;
    defparam sAddress_RNI9IH12_1_3_LC_17_5_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_1_3_LC_17_5_6.LUT_INIT=16'b0100000000000000;
    LogicCell40 sAddress_RNI9IH12_1_3_LC_17_5_6 (
            .in0(N__40608),
            .in1(N__46249),
            .in2(N__40422),
            .in3(N__40408),
            .lcout(sDAC_mem_38_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_35_0_LC_17_6_0.C_ON=1'b0;
    defparam sDAC_mem_35_0_LC_17_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_0_LC_17_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_0_LC_17_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51155),
            .lcout(sDAC_mem_35Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47750),
            .ce(N__40710),
            .sr(N__53113));
    defparam sDAC_mem_35_1_LC_17_6_1.C_ON=1'b0;
    defparam sDAC_mem_35_1_LC_17_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_1_LC_17_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_1_LC_17_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50707),
            .lcout(sDAC_mem_35Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47750),
            .ce(N__40710),
            .sr(N__53113));
    defparam sDAC_mem_35_2_LC_17_6_2.C_ON=1'b0;
    defparam sDAC_mem_35_2_LC_17_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_2_LC_17_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_2_LC_17_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50242),
            .lcout(sDAC_mem_35Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47750),
            .ce(N__40710),
            .sr(N__53113));
    defparam sDAC_mem_35_3_LC_17_6_3.C_ON=1'b0;
    defparam sDAC_mem_35_3_LC_17_6_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_3_LC_17_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_3_LC_17_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49767),
            .lcout(sDAC_mem_35Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47750),
            .ce(N__40710),
            .sr(N__53113));
    defparam sDAC_mem_35_4_LC_17_6_4.C_ON=1'b0;
    defparam sDAC_mem_35_4_LC_17_6_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_4_LC_17_6_4.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_35_4_LC_17_6_4 (
            .in0(_gnd_net_),
            .in1(N__49356),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_35Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47750),
            .ce(N__40710),
            .sr(N__53113));
    defparam sDAC_mem_35_5_LC_17_6_5.C_ON=1'b0;
    defparam sDAC_mem_35_5_LC_17_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_5_LC_17_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_5_LC_17_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46986),
            .lcout(sDAC_mem_35Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47750),
            .ce(N__40710),
            .sr(N__53113));
    defparam sDAC_mem_35_6_LC_17_6_6.C_ON=1'b0;
    defparam sDAC_mem_35_6_LC_17_6_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_6_LC_17_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_6_LC_17_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48213),
            .lcout(sDAC_mem_35Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47750),
            .ce(N__40710),
            .sr(N__53113));
    defparam sDAC_mem_35_7_LC_17_6_7.C_ON=1'b0;
    defparam sDAC_mem_35_7_LC_17_6_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_35_7_LC_17_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_35_7_LC_17_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48797),
            .lcout(sDAC_mem_35Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47750),
            .ce(N__40710),
            .sr(N__53113));
    defparam sDAC_mem_21_0_LC_17_7_0.C_ON=1'b0;
    defparam sDAC_mem_21_0_LC_17_7_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_0_LC_17_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_0_LC_17_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51157),
            .lcout(sDAC_mem_21Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47737),
            .ce(N__40674),
            .sr(N__53101));
    defparam sDAC_mem_21_1_LC_17_7_1.C_ON=1'b0;
    defparam sDAC_mem_21_1_LC_17_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_1_LC_17_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_1_LC_17_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50708),
            .lcout(sDAC_mem_21Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47737),
            .ce(N__40674),
            .sr(N__53101));
    defparam sDAC_mem_21_2_LC_17_7_2.C_ON=1'b0;
    defparam sDAC_mem_21_2_LC_17_7_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_2_LC_17_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_2_LC_17_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50243),
            .lcout(sDAC_mem_21Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47737),
            .ce(N__40674),
            .sr(N__53101));
    defparam sDAC_mem_21_3_LC_17_7_3.C_ON=1'b0;
    defparam sDAC_mem_21_3_LC_17_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_3_LC_17_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_3_LC_17_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49768),
            .lcout(sDAC_mem_21Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47737),
            .ce(N__40674),
            .sr(N__53101));
    defparam sDAC_mem_21_4_LC_17_7_4.C_ON=1'b0;
    defparam sDAC_mem_21_4_LC_17_7_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_4_LC_17_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_4_LC_17_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49207),
            .lcout(sDAC_mem_21Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47737),
            .ce(N__40674),
            .sr(N__53101));
    defparam sDAC_mem_21_5_LC_17_7_5.C_ON=1'b0;
    defparam sDAC_mem_21_5_LC_17_7_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_5_LC_17_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_5_LC_17_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46983),
            .lcout(sDAC_mem_21Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47737),
            .ce(N__40674),
            .sr(N__53101));
    defparam sDAC_mem_21_6_LC_17_7_6.C_ON=1'b0;
    defparam sDAC_mem_21_6_LC_17_7_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_6_LC_17_7_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_21_6_LC_17_7_6 (
            .in0(N__48214),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_21Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47737),
            .ce(N__40674),
            .sr(N__53101));
    defparam sDAC_mem_21_7_LC_17_7_7.C_ON=1'b0;
    defparam sDAC_mem_21_7_LC_17_7_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_21_7_LC_17_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_21_7_LC_17_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48741),
            .lcout(sDAC_mem_21Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47737),
            .ce(N__40674),
            .sr(N__53101));
    defparam sDAC_data_RNO_13_6_LC_17_8_0.C_ON=1'b0;
    defparam sDAC_data_RNO_13_6_LC_17_8_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_6_LC_17_8_0.LUT_INIT=16'b0001110000011111;
    LogicCell40 sDAC_data_RNO_13_6_LC_17_8_0 (
            .in0(N__41634),
            .in1(N__51812),
            .in2(N__43636),
            .in3(N__40830),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_6_LC_17_8_1.C_ON=1'b0;
    defparam sDAC_data_RNO_5_6_LC_17_8_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_6_LC_17_8_1.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_5_6_LC_17_8_1 (
            .in0(N__40857),
            .in1(N__52120),
            .in2(N__40845),
            .in3(N__40842),
            .lcout(sDAC_data_RNO_5Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_6_3_LC_17_8_2.C_ON=1'b0;
    defparam sDAC_mem_6_3_LC_17_8_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_3_LC_17_8_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_6_3_LC_17_8_2 (
            .in0(N__49769),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_6Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47727),
            .ce(N__43085),
            .sr(N__53087));
    defparam sDAC_mem_6_4_LC_17_8_5.C_ON=1'b0;
    defparam sDAC_mem_6_4_LC_17_8_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_4_LC_17_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_4_LC_17_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49312),
            .lcout(sDAC_mem_6Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47727),
            .ce(N__43085),
            .sr(N__53087));
    defparam sDAC_data_RNO_13_8_LC_17_8_6.C_ON=1'b0;
    defparam sDAC_data_RNO_13_8_LC_17_8_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_8_LC_17_8_6.LUT_INIT=16'b0001110000011111;
    LogicCell40 sDAC_data_RNO_13_8_LC_17_8_6 (
            .in0(N__41889),
            .in1(N__51813),
            .in2(N__43637),
            .in3(N__40818),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_8_LC_17_8_7.C_ON=1'b0;
    defparam sDAC_data_RNO_5_8_LC_17_8_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_8_LC_17_8_7.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_5_8_LC_17_8_7 (
            .in0(N__40806),
            .in1(N__52121),
            .in2(N__40794),
            .in3(N__40791),
            .lcout(sDAC_data_RNO_5Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_8_LC_17_9_0.C_ON=1'b0;
    defparam sDAC_data_RNO_10_8_LC_17_9_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_8_LC_17_9_0.LUT_INIT=16'b1100101100001011;
    LogicCell40 sDAC_data_RNO_10_8_LC_17_9_0 (
            .in0(N__40779),
            .in1(N__45870),
            .in2(N__40734),
            .in3(N__40767),
            .lcout(sDAC_data_RNO_10Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_8_LC_17_9_1.C_ON=1'b0;
    defparam sDAC_data_RNO_22_8_LC_17_9_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_8_LC_17_9_1.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_22_8_LC_17_9_1 (
            .in0(N__45868),
            .in1(N__45526),
            .in2(N__40758),
            .in3(N__40746),
            .lcout(sDAC_data_2_32_ns_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_8_LC_17_9_2.C_ON=1'b0;
    defparam sDAC_data_RNO_6_8_LC_17_9_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_8_LC_17_9_2.LUT_INIT=16'b0100011001010111;
    LogicCell40 sDAC_data_RNO_6_8_LC_17_9_2 (
            .in0(N__45527),
            .in1(N__45869),
            .in2(N__40989),
            .in3(N__40977),
            .lcout(),
            .ltout(sDAC_data_2_14_ns_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_8_LC_17_9_3.C_ON=1'b0;
    defparam sDAC_data_RNO_1_8_LC_17_9_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_8_LC_17_9_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_1_8_LC_17_9_3 (
            .in0(N__45871),
            .in1(N__40968),
            .in2(N__40962),
            .in3(N__40959),
            .lcout(sDAC_data_RNO_1Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_8_LC_17_9_4.C_ON=1'b0;
    defparam sDAC_data_RNO_3_8_LC_17_9_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_8_LC_17_9_4.LUT_INIT=16'b0001101101010101;
    LogicCell40 sDAC_data_RNO_3_8_LC_17_9_4 (
            .in0(N__42639),
            .in1(N__40953),
            .in2(N__40947),
            .in3(N__42525),
            .lcout(),
            .ltout(sDAC_data_2_41_ns_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_8_LC_17_9_5.C_ON=1'b0;
    defparam sDAC_data_RNO_0_8_LC_17_9_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_8_LC_17_9_5.LUT_INIT=16'b0101111000001110;
    LogicCell40 sDAC_data_RNO_0_8_LC_17_9_5 (
            .in0(N__42526),
            .in1(N__42771),
            .in2(N__40929),
            .in3(N__40926),
            .lcout(),
            .ltout(sDAC_data_2_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_8_LC_17_9_6.C_ON=1'b0;
    defparam sDAC_data_8_LC_17_9_6.SEQ_MODE=4'b1010;
    defparam sDAC_data_8_LC_17_9_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 sDAC_data_8_LC_17_9_6 (
            .in0(_gnd_net_),
            .in1(N__47262),
            .in2(N__40920),
            .in3(N__42383),
            .lcout(sDAC_dataZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53258),
            .ce(N__42223),
            .sr(N__53075));
    defparam sDAC_mem_3_1_LC_17_10_0.C_ON=1'b0;
    defparam sDAC_mem_3_1_LC_17_10_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_1_LC_17_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_3_1_LC_17_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50740),
            .lcout(sDAC_mem_3Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47714),
            .ce(N__42985),
            .sr(N__53064));
    defparam sDAC_data_RNO_28_4_LC_17_10_1.C_ON=1'b0;
    defparam sDAC_data_RNO_28_4_LC_17_10_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_4_LC_17_10_1.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_28_4_LC_17_10_1 (
            .in0(N__52109),
            .in1(N__43628),
            .in2(N__40899),
            .in3(N__40884),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_4_LC_17_10_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_4_LC_17_10_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_4_LC_17_10_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_4_LC_17_10_2 (
            .in0(N__52107),
            .in1(N__40875),
            .in2(N__40866),
            .in3(N__40863),
            .lcout(sDAC_data_RNO_15Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_6_LC_17_10_3.C_ON=1'b0;
    defparam sDAC_data_RNO_17_6_LC_17_10_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_6_LC_17_10_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_6_LC_17_10_3 (
            .in0(N__43629),
            .in1(N__44172),
            .in2(_gnd_net_),
            .in3(N__44304),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_6_LC_17_10_4.C_ON=1'b0;
    defparam sDAC_data_RNO_8_6_LC_17_10_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_6_LC_17_10_4.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_8_6_LC_17_10_4 (
            .in0(_gnd_net_),
            .in1(N__52110),
            .in2(N__41103),
            .in3(N__45192),
            .lcout(sDAC_data_RNO_8Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_6_LC_17_10_5.C_ON=1'b0;
    defparam sDAC_data_RNO_16_6_LC_17_10_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_6_LC_17_10_5.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_16_6_LC_17_10_5 (
            .in0(N__52111),
            .in1(N__41820),
            .in2(N__43670),
            .in3(N__41100),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_6_LC_17_10_6.C_ON=1'b0;
    defparam sDAC_data_RNO_7_6_LC_17_10_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_6_LC_17_10_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_7_6_LC_17_10_6 (
            .in0(N__52108),
            .in1(N__43959),
            .in2(N__41088),
            .in3(N__47178),
            .lcout(),
            .ltout(sDAC_data_RNO_7Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_6_LC_17_10_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_6_LC_17_10_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_6_LC_17_10_7.LUT_INIT=16'b0111001101100010;
    LogicCell40 sDAC_data_RNO_2_6_LC_17_10_7 (
            .in0(N__45873),
            .in1(N__41085),
            .in2(N__41073),
            .in3(N__41070),
            .lcout(sDAC_data_RNO_2Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_4_LC_17_11_0.C_ON=1'b0;
    defparam sDAC_data_RNO_10_4_LC_17_11_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_4_LC_17_11_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_10_4_LC_17_11_0 (
            .in0(N__41265),
            .in1(N__41943),
            .in2(N__45945),
            .in3(N__41049),
            .lcout(),
            .ltout(sDAC_data_RNO_10Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_4_LC_17_11_1.C_ON=1'b0;
    defparam sDAC_data_RNO_3_4_LC_17_11_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_4_LC_17_11_1.LUT_INIT=16'b0001010110011101;
    LogicCell40 sDAC_data_RNO_3_4_LC_17_11_1 (
            .in0(N__42641),
            .in1(N__42531),
            .in2(N__41064),
            .in3(N__41577),
            .lcout(sDAC_data_2_41_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_4_LC_17_11_2.C_ON=1'b0;
    defparam sDAC_data_RNO_22_4_LC_17_11_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_4_LC_17_11_2.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_22_4_LC_17_11_2 (
            .in0(N__45938),
            .in1(N__45528),
            .in2(N__41676),
            .in3(N__41061),
            .lcout(sDAC_data_2_32_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_4_LC_17_11_3.C_ON=1'b0;
    defparam sDAC_data_RNO_6_4_LC_17_11_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_4_LC_17_11_3.LUT_INIT=16'b0100011001010111;
    LogicCell40 sDAC_data_RNO_6_4_LC_17_11_3 (
            .in0(N__45529),
            .in1(N__45942),
            .in2(N__41043),
            .in3(N__41031),
            .lcout(),
            .ltout(sDAC_data_2_14_ns_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_4_LC_17_11_4.C_ON=1'b0;
    defparam sDAC_data_RNO_1_4_LC_17_11_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_4_LC_17_11_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_1_4_LC_17_11_4 (
            .in0(N__45943),
            .in1(N__41019),
            .in2(N__41004),
            .in3(N__41001),
            .lcout(),
            .ltout(sDAC_data_RNO_1Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_4_LC_17_11_5.C_ON=1'b0;
    defparam sDAC_data_RNO_0_4_LC_17_11_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_4_LC_17_11_5.LUT_INIT=16'b0101000011101110;
    LogicCell40 sDAC_data_RNO_0_4_LC_17_11_5 (
            .in0(N__42530),
            .in1(N__43299),
            .in2(N__41214),
            .in3(N__41211),
            .lcout(),
            .ltout(sDAC_data_2_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_4_LC_17_11_6.C_ON=1'b0;
    defparam sDAC_data_4_LC_17_11_6.SEQ_MODE=4'b1010;
    defparam sDAC_data_4_LC_17_11_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 sDAC_data_4_LC_17_11_6 (
            .in0(_gnd_net_),
            .in1(N__46002),
            .in2(N__41205),
            .in3(N__42366),
            .lcout(sDAC_dataZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53269),
            .ce(N__42224),
            .sr(N__53054));
    defparam sDAC_data_RNO_10_3_LC_17_12_0.C_ON=1'b0;
    defparam sDAC_data_RNO_10_3_LC_17_12_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_3_LC_17_12_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_10_3_LC_17_12_0 (
            .in0(N__41190),
            .in1(N__41967),
            .in2(N__45909),
            .in3(N__41166),
            .lcout(),
            .ltout(sDAC_data_RNO_10Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_3_LC_17_12_1.C_ON=1'b0;
    defparam sDAC_data_RNO_3_3_LC_17_12_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_3_LC_17_12_1.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_3_3_LC_17_12_1 (
            .in0(N__42522),
            .in1(N__42642),
            .in2(N__41178),
            .in3(N__41385),
            .lcout(sDAC_data_2_41_ns_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_3_LC_17_12_2.C_ON=1'b0;
    defparam sDAC_data_RNO_22_3_LC_17_12_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_3_LC_17_12_2.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_22_3_LC_17_12_2 (
            .in0(N__45883),
            .in1(N__45457),
            .in2(N__44070),
            .in3(N__41175),
            .lcout(sDAC_data_2_32_ns_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_3_LC_17_12_3.C_ON=1'b0;
    defparam sDAC_data_RNO_6_3_LC_17_12_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_3_LC_17_12_3.LUT_INIT=16'b0100011001010111;
    LogicCell40 sDAC_data_RNO_6_3_LC_17_12_3 (
            .in0(N__45458),
            .in1(N__45887),
            .in2(N__41160),
            .in3(N__41142),
            .lcout(),
            .ltout(sDAC_data_2_14_ns_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_1_3_LC_17_12_4.C_ON=1'b0;
    defparam sDAC_data_RNO_1_3_LC_17_12_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_3_LC_17_12_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_1_3_LC_17_12_4 (
            .in0(N__45888),
            .in1(N__41136),
            .in2(N__41121),
            .in3(N__41118),
            .lcout(),
            .ltout(sDAC_data_RNO_1Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_3_LC_17_12_5.C_ON=1'b0;
    defparam sDAC_data_RNO_0_3_LC_17_12_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_3_LC_17_12_5.LUT_INIT=16'b0101000011101110;
    LogicCell40 sDAC_data_RNO_0_3_LC_17_12_5 (
            .in0(N__42523),
            .in1(N__43002),
            .in2(N__41112),
            .in3(N__41109),
            .lcout(),
            .ltout(sDAC_data_2_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_3_LC_17_12_6.C_ON=1'b0;
    defparam sDAC_data_3_LC_17_12_6.SEQ_MODE=4'b1010;
    defparam sDAC_data_3_LC_17_12_6.LUT_INIT=16'b1110010011100100;
    LogicCell40 sDAC_data_3_LC_17_12_6 (
            .in0(N__42377),
            .in1(N__46017),
            .in2(N__41373),
            .in3(_gnd_net_),
            .lcout(sDAC_dataZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53271),
            .ce(N__42226),
            .sr(N__53044));
    defparam sDAC_data_RNO_29_10_LC_17_13_0.C_ON=1'b0;
    defparam sDAC_data_RNO_29_10_LC_17_13_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_10_LC_17_13_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_29_10_LC_17_13_0 (
            .in0(N__41352),
            .in1(N__51993),
            .in2(_gnd_net_),
            .in3(N__41337),
            .lcout(sDAC_data_RNO_29Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_30_6_LC_17_13_2.C_ON=1'b0;
    defparam sDAC_data_RNO_30_6_LC_17_13_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_30_6_LC_17_13_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_30_6_LC_17_13_2 (
            .in0(N__41316),
            .in1(N__51994),
            .in2(_gnd_net_),
            .in3(N__41304),
            .lcout(sDAC_data_RNO_30Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_3_5_LC_17_13_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_3_5_LC_17_13_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_3_5_LC_17_13_3.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNI9IH12_3_5_LC_17_13_3 (
            .in0(N__44430),
            .in1(N__46574),
            .in2(N__46251),
            .in3(N__46322),
            .lcout(sDAC_mem_14_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_21_4_LC_17_13_6.C_ON=1'b0;
    defparam sDAC_data_RNO_21_4_LC_17_13_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_21_4_LC_17_13_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_21_4_LC_17_13_6 (
            .in0(N__52153),
            .in1(N__41295),
            .in2(_gnd_net_),
            .in3(N__41280),
            .lcout(sDAC_data_RNO_21Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_27_1_LC_17_14_1.C_ON=1'b0;
    defparam sDAC_mem_27_1_LC_17_14_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_1_LC_17_14_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_27_1_LC_17_14_1 (
            .in0(N__50761),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_27Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47728),
            .ce(N__45245),
            .sr(N__53025));
    defparam sDAC_mem_27_2_LC_17_14_2.C_ON=1'b0;
    defparam sDAC_mem_27_2_LC_17_14_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_2_LC_17_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_2_LC_17_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50174),
            .lcout(sDAC_mem_27Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47728),
            .ce(N__45245),
            .sr(N__53025));
    defparam sDAC_mem_27_3_LC_17_14_3.C_ON=1'b0;
    defparam sDAC_mem_27_3_LC_17_14_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_3_LC_17_14_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_27_3_LC_17_14_3 (
            .in0(N__49794),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_27Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47728),
            .ce(N__45245),
            .sr(N__53025));
    defparam sDAC_mem_27_4_LC_17_14_4.C_ON=1'b0;
    defparam sDAC_mem_27_4_LC_17_14_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_4_LC_17_14_4.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_27_4_LC_17_14_4 (
            .in0(_gnd_net_),
            .in1(N__49231),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_27Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47728),
            .ce(N__45245),
            .sr(N__53025));
    defparam sDAC_mem_27_5_LC_17_14_5.C_ON=1'b0;
    defparam sDAC_mem_27_5_LC_17_14_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_5_LC_17_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_5_LC_17_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47081),
            .lcout(sDAC_mem_27Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47728),
            .ce(N__45245),
            .sr(N__53025));
    defparam sDAC_mem_27_6_LC_17_14_6.C_ON=1'b0;
    defparam sDAC_mem_27_6_LC_17_14_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_6_LC_17_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_6_LC_17_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48331),
            .lcout(sDAC_mem_27Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47728),
            .ce(N__45245),
            .sr(N__53025));
    defparam sDAC_mem_27_7_LC_17_14_7.C_ON=1'b0;
    defparam sDAC_mem_27_7_LC_17_14_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_7_LC_17_14_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_27_7_LC_17_14_7 (
            .in0(_gnd_net_),
            .in1(N__48841),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_27Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47728),
            .ce(N__45245),
            .sr(N__53025));
    defparam sEEADC_freq_0_LC_17_15_0.C_ON=1'b0;
    defparam sEEADC_freq_0_LC_17_15_0.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_0_LC_17_15_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEADC_freq_0_LC_17_15_0 (
            .in0(N__51269),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEADC_freqZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47738),
            .ce(N__44122),
            .sr(_gnd_net_));
    defparam sEEADC_freq_6_LC_17_15_1.C_ON=1'b0;
    defparam sEEADC_freq_6_LC_17_15_1.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_6_LC_17_15_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 sEEADC_freq_6_LC_17_15_1 (
            .in0(_gnd_net_),
            .in1(N__48332),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEADC_freqZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47738),
            .ce(N__44122),
            .sr(_gnd_net_));
    defparam sEEADC_freq_7_LC_17_15_2.C_ON=1'b0;
    defparam sEEADC_freq_7_LC_17_15_2.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_7_LC_17_15_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEADC_freq_7_LC_17_15_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48818),
            .lcout(sEEADC_freqZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47738),
            .ce(N__44122),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_24_3_LC_17_16_0.C_ON=1'b0;
    defparam sDAC_data_RNO_24_3_LC_17_16_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_24_3_LC_17_16_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_24_3_LC_17_16_0 (
            .in0(N__51771),
            .in1(N__41427),
            .in2(_gnd_net_),
            .in3(N__41415),
            .lcout(sDAC_data_RNO_24Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_23_3_LC_17_16_1.C_ON=1'b0;
    defparam sDAC_data_RNO_23_3_LC_17_16_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_23_3_LC_17_16_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_23_3_LC_17_16_1 (
            .in0(N__52073),
            .in1(N__41409),
            .in2(_gnd_net_),
            .in3(N__41613),
            .lcout(),
            .ltout(sDAC_data_RNO_23Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_3_LC_17_16_2.C_ON=1'b0;
    defparam sDAC_data_RNO_11_3_LC_17_16_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_3_LC_17_16_2.LUT_INIT=16'b1010000011011101;
    LogicCell40 sDAC_data_RNO_11_3_LC_17_16_2 (
            .in0(N__45879),
            .in1(N__41400),
            .in2(N__41394),
            .in3(N__41391),
            .lcout(sDAC_data_RNO_11Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_28_0_LC_17_16_3.C_ON=1'b0;
    defparam sDAC_mem_28_0_LC_17_16_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_0_LC_17_16_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_0_LC_17_16_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51272),
            .lcout(sDAC_mem_28Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47751),
            .ce(N__41777),
            .sr(N__53014));
    defparam sDAC_data_RNO_31_4_LC_17_16_4.C_ON=1'b0;
    defparam sDAC_data_RNO_31_4_LC_17_16_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_31_4_LC_17_16_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 sDAC_data_RNO_31_4_LC_17_16_4 (
            .in0(N__51772),
            .in1(N__41607),
            .in2(_gnd_net_),
            .in3(N__41736),
            .lcout(),
            .ltout(sDAC_data_RNO_31Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_25_4_LC_17_16_5.C_ON=1'b0;
    defparam sDAC_data_RNO_25_4_LC_17_16_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_25_4_LC_17_16_5.LUT_INIT=16'b0010001101100111;
    LogicCell40 sDAC_data_RNO_25_4_LC_17_16_5 (
            .in0(N__45881),
            .in1(N__45501),
            .in2(N__41595),
            .in3(N__41547),
            .lcout(),
            .ltout(sDAC_data_2_39_ns_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_11_4_LC_17_16_6.C_ON=1'b0;
    defparam sDAC_data_RNO_11_4_LC_17_16_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_11_4_LC_17_16_6.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_11_4_LC_17_16_6 (
            .in0(N__45880),
            .in1(N__41592),
            .in2(N__41586),
            .in3(N__41583),
            .lcout(sDAC_data_RNO_11Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_32_4_LC_17_16_7.C_ON=1'b0;
    defparam sDAC_data_RNO_32_4_LC_17_16_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_32_4_LC_17_16_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 sDAC_data_RNO_32_4_LC_17_16_7 (
            .in0(N__41568),
            .in1(N__51770),
            .in2(_gnd_net_),
            .in3(N__41556),
            .lcout(sDAC_data_RNO_32Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_28_1_LC_17_17_0.C_ON=1'b0;
    defparam sDAC_mem_28_1_LC_17_17_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_1_LC_17_17_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_1_LC_17_17_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50771),
            .lcout(sDAC_mem_28Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47762),
            .ce(N__41776),
            .sr(N__53005));
    defparam sDAC_mem_28_2_LC_17_17_1.C_ON=1'b0;
    defparam sDAC_mem_28_2_LC_17_17_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_2_LC_17_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_2_LC_17_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50256),
            .lcout(sDAC_mem_28Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47762),
            .ce(N__41776),
            .sr(N__53005));
    defparam sDAC_mem_28_4_LC_17_17_2.C_ON=1'b0;
    defparam sDAC_mem_28_4_LC_17_17_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_4_LC_17_17_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_4_LC_17_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49305),
            .lcout(sDAC_mem_28Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47762),
            .ce(N__41776),
            .sr(N__53005));
    defparam sDAC_mem_28_5_LC_17_17_3.C_ON=1'b0;
    defparam sDAC_mem_28_5_LC_17_17_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_5_LC_17_17_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_5_LC_17_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47133),
            .lcout(sDAC_mem_28Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47762),
            .ce(N__41776),
            .sr(N__53005));
    defparam sDAC_mem_28_7_LC_17_17_4.C_ON=1'b0;
    defparam sDAC_mem_28_7_LC_17_17_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_28_7_LC_17_17_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_28_7_LC_17_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48800),
            .lcout(sDAC_mem_28Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47762),
            .ce(N__41776),
            .sr(N__53005));
    defparam sAddress_RNI9IH12_1_LC_17_18_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_1_LC_17_18_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_1_LC_17_18_0.LUT_INIT=16'b0001000100000000;
    LogicCell40 sAddress_RNI9IH12_1_LC_17_18_0 (
            .in0(N__46428),
            .in1(N__46132),
            .in2(_gnd_net_),
            .in3(N__43189),
            .lcout(sDAC_mem_25_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_25_1_LC_17_18_2.C_ON=1'b0;
    defparam sDAC_mem_25_1_LC_17_18_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_25_1_LC_17_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_25_1_LC_17_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50772),
            .lcout(sDAC_mem_25Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47774),
            .ce(N__41716),
            .sr(N__52996));
    defparam sDAC_data_RNO_29_4_LC_17_19_4.C_ON=1'b0;
    defparam sDAC_data_RNO_29_4_LC_17_19_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_4_LC_17_19_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_29_4_LC_17_19_4 (
            .in0(N__41694),
            .in1(N__51551),
            .in2(_gnd_net_),
            .in3(N__45219),
            .lcout(sDAC_data_RNO_29Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_38_6_LC_18_4_0.C_ON=1'b0;
    defparam sDAC_mem_38_6_LC_18_4_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_6_LC_18_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_6_LC_18_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48227),
            .lcout(sDAC_mem_38Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47763),
            .ce(N__41867),
            .sr(N__53139));
    defparam sDAC_mem_38_0_LC_18_5_0.C_ON=1'b0;
    defparam sDAC_mem_38_0_LC_18_5_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_0_LC_18_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_0_LC_18_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51156),
            .lcout(sDAC_mem_38Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47752),
            .ce(N__41866),
            .sr(N__53134));
    defparam sDAC_mem_38_2_LC_18_5_2.C_ON=1'b0;
    defparam sDAC_mem_38_2_LC_18_5_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_2_LC_18_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_2_LC_18_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50078),
            .lcout(sDAC_mem_38Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47752),
            .ce(N__41866),
            .sr(N__53134));
    defparam sDAC_mem_38_3_LC_18_5_3.C_ON=1'b0;
    defparam sDAC_mem_38_3_LC_18_5_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_3_LC_18_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_3_LC_18_5_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49734),
            .lcout(sDAC_mem_38Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47752),
            .ce(N__41866),
            .sr(N__53134));
    defparam sDAC_mem_38_4_LC_18_5_4.C_ON=1'b0;
    defparam sDAC_mem_38_4_LC_18_5_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_4_LC_18_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_4_LC_18_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49362),
            .lcout(sDAC_mem_38Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47752),
            .ce(N__41866),
            .sr(N__53134));
    defparam sDAC_mem_38_5_LC_18_5_5.C_ON=1'b0;
    defparam sDAC_mem_38_5_LC_18_5_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_5_LC_18_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_5_LC_18_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47099),
            .lcout(sDAC_mem_38Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47752),
            .ce(N__41866),
            .sr(N__53134));
    defparam sDAC_mem_38_7_LC_18_5_7.C_ON=1'b0;
    defparam sDAC_mem_38_7_LC_18_5_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_38_7_LC_18_5_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_38_7_LC_18_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48742),
            .lcout(sDAC_mem_38Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47752),
            .ce(N__41866),
            .sr(N__53134));
    defparam sDAC_mem_40_0_LC_18_6_0.C_ON=1'b0;
    defparam sDAC_mem_40_0_LC_18_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_0_LC_18_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_0_LC_18_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51158),
            .lcout(sDAC_mem_40Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47739),
            .ce(N__41985),
            .sr(N__53128));
    defparam sDAC_mem_40_1_LC_18_6_1.C_ON=1'b0;
    defparam sDAC_mem_40_1_LC_18_6_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_1_LC_18_6_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_1_LC_18_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50709),
            .lcout(sDAC_mem_40Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47739),
            .ce(N__41985),
            .sr(N__53128));
    defparam sDAC_mem_40_2_LC_18_6_2.C_ON=1'b0;
    defparam sDAC_mem_40_2_LC_18_6_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_2_LC_18_6_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_2_LC_18_6_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50079),
            .lcout(sDAC_mem_40Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47739),
            .ce(N__41985),
            .sr(N__53128));
    defparam sDAC_mem_40_3_LC_18_6_3.C_ON=1'b0;
    defparam sDAC_mem_40_3_LC_18_6_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_3_LC_18_6_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_40_3_LC_18_6_3 (
            .in0(N__49735),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_40Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47739),
            .ce(N__41985),
            .sr(N__53128));
    defparam sDAC_mem_40_4_LC_18_6_4.C_ON=1'b0;
    defparam sDAC_mem_40_4_LC_18_6_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_4_LC_18_6_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_4_LC_18_6_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49363),
            .lcout(sDAC_mem_40Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47739),
            .ce(N__41985),
            .sr(N__53128));
    defparam sDAC_mem_40_5_LC_18_6_5.C_ON=1'b0;
    defparam sDAC_mem_40_5_LC_18_6_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_5_LC_18_6_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_5_LC_18_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47071),
            .lcout(sDAC_mem_40Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47739),
            .ce(N__41985),
            .sr(N__53128));
    defparam sDAC_mem_40_6_LC_18_6_6.C_ON=1'b0;
    defparam sDAC_mem_40_6_LC_18_6_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_6_LC_18_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_6_LC_18_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48228),
            .lcout(sDAC_mem_40Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47739),
            .ce(N__41985),
            .sr(N__53128));
    defparam sDAC_mem_40_7_LC_18_6_7.C_ON=1'b0;
    defparam sDAC_mem_40_7_LC_18_6_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_40_7_LC_18_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_40_7_LC_18_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48743),
            .lcout(sDAC_mem_40Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47739),
            .ce(N__41985),
            .sr(N__53128));
    defparam sDAC_data_RNO_20_3_LC_18_7_0.C_ON=1'b0;
    defparam sDAC_data_RNO_20_3_LC_18_7_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_3_LC_18_7_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_20_3_LC_18_7_0 (
            .in0(N__52003),
            .in1(N__41973),
            .in2(_gnd_net_),
            .in3(N__41955),
            .lcout(sDAC_data_RNO_20Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_20_0_LC_18_7_1.C_ON=1'b0;
    defparam sDAC_mem_20_0_LC_18_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_0_LC_18_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_0_LC_18_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51164),
            .lcout(sDAC_mem_20Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47729),
            .ce(N__44030),
            .sr(N__53114));
    defparam sDAC_data_RNO_20_4_LC_18_7_2.C_ON=1'b0;
    defparam sDAC_data_RNO_20_4_LC_18_7_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_4_LC_18_7_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_20_4_LC_18_7_2 (
            .in0(N__52004),
            .in1(N__41949),
            .in2(_gnd_net_),
            .in3(N__41931),
            .lcout(sDAC_data_RNO_20Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_20_1_LC_18_7_3.C_ON=1'b0;
    defparam sDAC_mem_20_1_LC_18_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_1_LC_18_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_1_LC_18_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50710),
            .lcout(sDAC_mem_20Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47729),
            .ce(N__44030),
            .sr(N__53114));
    defparam sDAC_data_RNO_20_5_LC_18_7_4.C_ON=1'b0;
    defparam sDAC_data_RNO_20_5_LC_18_7_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_5_LC_18_7_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_20_5_LC_18_7_4 (
            .in0(N__52005),
            .in1(N__41925),
            .in2(_gnd_net_),
            .in3(N__41910),
            .lcout(sDAC_data_RNO_20Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_20_2_LC_18_7_5.C_ON=1'b0;
    defparam sDAC_mem_20_2_LC_18_7_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_2_LC_18_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_2_LC_18_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50080),
            .lcout(sDAC_mem_20Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47729),
            .ce(N__44030),
            .sr(N__53114));
    defparam sDAC_data_RNO_20_6_LC_18_7_6.C_ON=1'b0;
    defparam sDAC_data_RNO_20_6_LC_18_7_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_20_6_LC_18_7_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_20_6_LC_18_7_6 (
            .in0(N__52006),
            .in1(N__41904),
            .in2(_gnd_net_),
            .in3(N__41895),
            .lcout(sDAC_data_RNO_20Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_20_3_LC_18_7_7.C_ON=1'b0;
    defparam sDAC_mem_20_3_LC_18_7_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_3_LC_18_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_3_LC_18_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49736),
            .lcout(sDAC_mem_20Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47729),
            .ce(N__44030),
            .sr(N__53114));
    defparam sDAC_data_RNO_26_6_LC_18_8_0.C_ON=1'b0;
    defparam sDAC_data_RNO_26_6_LC_18_8_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_6_LC_18_8_0.LUT_INIT=16'b0111010000110000;
    LogicCell40 sDAC_data_RNO_26_6_LC_18_8_0 (
            .in0(N__43579),
            .in1(N__51804),
            .in2(N__42144),
            .in3(N__42114),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_6_LC_18_8_1.C_ON=1'b0;
    defparam sDAC_data_RNO_14_6_LC_18_8_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_6_LC_18_8_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_14_6_LC_18_8_1 (
            .in0(_gnd_net_),
            .in1(N__42159),
            .in2(N__42147),
            .in3(N__42120),
            .lcout(sDAC_data_RNO_14Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_27_6_LC_18_8_2.C_ON=1'b0;
    defparam sDAC_data_RNO_27_6_LC_18_8_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_6_LC_18_8_2.LUT_INIT=16'b1111110010111000;
    LogicCell40 sDAC_data_RNO_27_6_LC_18_8_2 (
            .in0(N__43577),
            .in1(N__51802),
            .in2(N__42143),
            .in3(N__42113),
            .lcout(sDAC_data_RNO_27Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_1_3_LC_18_8_3.C_ON=1'b0;
    defparam sDAC_mem_1_3_LC_18_8_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_3_LC_18_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_1_3_LC_18_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49824),
            .lcout(sDAC_mem_1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47719),
            .ce(N__42039),
            .sr(N__53102));
    defparam sDAC_data_RNO_26_7_LC_18_8_4.C_ON=1'b0;
    defparam sDAC_data_RNO_26_7_LC_18_8_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_26_7_LC_18_8_4.LUT_INIT=16'b0111010000110000;
    LogicCell40 sDAC_data_RNO_26_7_LC_18_8_4 (
            .in0(N__43578),
            .in1(N__51803),
            .in2(N__42078),
            .in3(N__42048),
            .lcout(),
            .ltout(sDAC_data_RNO_26Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_14_7_LC_18_8_5.C_ON=1'b0;
    defparam sDAC_data_RNO_14_7_LC_18_8_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_14_7_LC_18_8_5.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_14_7_LC_18_8_5 (
            .in0(_gnd_net_),
            .in1(N__42105),
            .in2(N__42096),
            .in3(N__42054),
            .lcout(sDAC_data_RNO_14Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_27_7_LC_18_8_6.C_ON=1'b0;
    defparam sDAC_data_RNO_27_7_LC_18_8_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_27_7_LC_18_8_6.LUT_INIT=16'b1111110010111000;
    LogicCell40 sDAC_data_RNO_27_7_LC_18_8_6 (
            .in0(N__43576),
            .in1(N__51801),
            .in2(N__42077),
            .in3(N__42047),
            .lcout(sDAC_data_RNO_27Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_1_4_LC_18_8_7.C_ON=1'b0;
    defparam sDAC_mem_1_4_LC_18_8_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_1_4_LC_18_8_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_1_4_LC_18_8_7 (
            .in0(N__49334),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47719),
            .ce(N__42039),
            .sr(N__53102));
    defparam sDAC_data_RNO_1_6_LC_18_9_0.C_ON=1'b0;
    defparam sDAC_data_RNO_1_6_LC_18_9_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_1_6_LC_18_9_0.LUT_INIT=16'b1100000010101111;
    LogicCell40 sDAC_data_RNO_1_6_LC_18_9_0 (
            .in0(N__42015),
            .in1(N__42009),
            .in2(N__45944),
            .in3(N__42708),
            .lcout(sDAC_data_RNO_1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_6_6_LC_18_9_1.C_ON=1'b0;
    defparam sDAC_data_RNO_6_6_LC_18_9_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_6_6_LC_18_9_1.LUT_INIT=16'b0010011000110111;
    LogicCell40 sDAC_data_RNO_6_6_LC_18_9_1 (
            .in0(N__45932),
            .in1(N__45524),
            .in2(N__42816),
            .in3(N__42714),
            .lcout(sDAC_data_2_14_ns_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_22_6_LC_18_9_2.C_ON=1'b0;
    defparam sDAC_data_RNO_22_6_LC_18_9_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_22_6_LC_18_9_2.LUT_INIT=16'b0100010101100111;
    LogicCell40 sDAC_data_RNO_22_6_LC_18_9_2 (
            .in0(N__45525),
            .in1(N__45933),
            .in2(N__42702),
            .in3(N__42681),
            .lcout(),
            .ltout(sDAC_data_2_32_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_10_6_LC_18_9_3.C_ON=1'b0;
    defparam sDAC_data_RNO_10_6_LC_18_9_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_10_6_LC_18_9_3.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_10_6_LC_18_9_3 (
            .in0(N__45934),
            .in1(N__42669),
            .in2(N__42654),
            .in3(N__42651),
            .lcout(),
            .ltout(sDAC_data_RNO_10Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_3_6_LC_18_9_4.C_ON=1'b0;
    defparam sDAC_data_RNO_3_6_LC_18_9_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_3_6_LC_18_9_4.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_3_6_LC_18_9_4 (
            .in0(N__42524),
            .in1(N__42640),
            .in2(N__42555),
            .in3(N__42552),
            .lcout(),
            .ltout(sDAC_data_2_41_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_0_6_LC_18_9_5.C_ON=1'b0;
    defparam sDAC_data_RNO_0_6_LC_18_9_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_0_6_LC_18_9_5.LUT_INIT=16'b0101111000001110;
    LogicCell40 sDAC_data_RNO_0_6_LC_18_9_5 (
            .in0(N__42527),
            .in1(N__42399),
            .in2(N__42393),
            .in3(N__42390),
            .lcout(),
            .ltout(sDAC_data_2_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_6_LC_18_9_6.C_ON=1'b0;
    defparam sDAC_data_6_LC_18_9_6.SEQ_MODE=4'b1010;
    defparam sDAC_data_6_LC_18_9_6.LUT_INIT=16'b1110010011100100;
    LogicCell40 sDAC_data_6_LC_18_9_6 (
            .in0(N__42384),
            .in1(N__45975),
            .in2(N__42255),
            .in3(_gnd_net_),
            .lcout(sDAC_dataZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53264),
            .ce(N__42221),
            .sr(N__53088));
    defparam sDAC_mem_3_3_LC_18_10_0.C_ON=1'b0;
    defparam sDAC_mem_3_3_LC_18_10_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_3_LC_18_10_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_3_3_LC_18_10_0 (
            .in0(N__49818),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_3Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47708),
            .ce(N__42992),
            .sr(N__53076));
    defparam sDAC_data_RNO_28_6_LC_18_10_1.C_ON=1'b0;
    defparam sDAC_data_RNO_28_6_LC_18_10_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_6_LC_18_10_1.LUT_INIT=16'b0100010101100111;
    LogicCell40 sDAC_data_RNO_28_6_LC_18_10_1 (
            .in0(N__43543),
            .in1(N__52141),
            .in2(N__42186),
            .in3(N__42171),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_6_LC_18_10_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_6_LC_18_10_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_6_LC_18_10_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_6_LC_18_10_2 (
            .in0(N__52142),
            .in1(N__42837),
            .in2(N__42825),
            .in3(N__42822),
            .lcout(sDAC_data_RNO_15Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_8_LC_18_10_3.C_ON=1'b0;
    defparam sDAC_data_RNO_17_8_LC_18_10_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_8_LC_18_10_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 sDAC_data_RNO_17_8_LC_18_10_3 (
            .in0(N__44376),
            .in1(_gnd_net_),
            .in2(N__43622),
            .in3(N__44277),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_8_LC_18_10_4.C_ON=1'b0;
    defparam sDAC_data_RNO_8_8_LC_18_10_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_8_LC_18_10_4.LUT_INIT=16'b1101100011011000;
    LogicCell40 sDAC_data_RNO_8_8_LC_18_10_4 (
            .in0(N__52143),
            .in1(N__45165),
            .in2(N__42807),
            .in3(_gnd_net_),
            .lcout(sDAC_data_RNO_8Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_8_LC_18_10_5.C_ON=1'b0;
    defparam sDAC_data_RNO_16_8_LC_18_10_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_8_LC_18_10_5.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_16_8_LC_18_10_5 (
            .in0(N__52144),
            .in1(N__42804),
            .in2(N__43623),
            .in3(N__42795),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_8_LC_18_10_6.C_ON=1'b0;
    defparam sDAC_data_RNO_7_8_LC_18_10_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_8_LC_18_10_6.LUT_INIT=16'b1000111110000011;
    LogicCell40 sDAC_data_RNO_7_8_LC_18_10_6 (
            .in0(N__46662),
            .in1(N__52145),
            .in2(N__42783),
            .in3(N__44244),
            .lcout(),
            .ltout(sDAC_data_RNO_7Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_8_LC_18_10_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_8_LC_18_10_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_8_LC_18_10_7.LUT_INIT=16'b0111001101100010;
    LogicCell40 sDAC_data_RNO_2_8_LC_18_10_7 (
            .in0(N__45872),
            .in1(N__43896),
            .in2(N__42780),
            .in3(N__42777),
            .lcout(sDAC_data_RNO_2Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_13_9_LC_18_11_0.C_ON=1'b0;
    defparam sDAC_data_RNO_13_9_LC_18_11_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_13_9_LC_18_11_0.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_13_9_LC_18_11_0 (
            .in0(N__52154),
            .in1(N__42765),
            .in2(N__43689),
            .in3(N__43095),
            .lcout(),
            .ltout(sDAC_data_2_13_bm_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_5_9_LC_18_11_1.C_ON=1'b0;
    defparam sDAC_data_RNO_5_9_LC_18_11_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_5_9_LC_18_11_1.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_5_9_LC_18_11_1 (
            .in0(N__52079),
            .in1(N__42756),
            .in2(N__42744),
            .in3(N__42741),
            .lcout(sDAC_data_RNO_5Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_6_6_LC_18_11_2.C_ON=1'b0;
    defparam sDAC_mem_6_6_LC_18_11_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_6_6_LC_18_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_6_6_LC_18_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48329),
            .lcout(sDAC_mem_6Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47704),
            .ce(N__43089),
            .sr(N__53065));
    defparam sDAC_data_RNO_16_3_LC_18_11_3.C_ON=1'b0;
    defparam sDAC_data_RNO_16_3_LC_18_11_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_3_LC_18_11_3.LUT_INIT=16'b0001101000011111;
    LogicCell40 sDAC_data_RNO_16_3_LC_18_11_3 (
            .in0(N__52078),
            .in1(N__43041),
            .in2(N__43688),
            .in3(N__43032),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_3_LC_18_11_4.C_ON=1'b0;
    defparam sDAC_data_RNO_7_3_LC_18_11_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_3_LC_18_11_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_7_3_LC_18_11_4 (
            .in0(N__52155),
            .in1(N__43998),
            .in2(N__43017),
            .in3(N__47217),
            .lcout(sDAC_data_RNO_7Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_3_LC_18_11_5.C_ON=1'b0;
    defparam sDAC_data_RNO_17_3_LC_18_11_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_3_LC_18_11_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_3_LC_18_11_5 (
            .in0(N__43682),
            .in1(N__44208),
            .in2(_gnd_net_),
            .in3(N__44340),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_3_LC_18_11_6.C_ON=1'b0;
    defparam sDAC_data_RNO_8_3_LC_18_11_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_3_LC_18_11_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_8_3_LC_18_11_6 (
            .in0(_gnd_net_),
            .in1(N__52080),
            .in2(N__43014),
            .in3(N__45012),
            .lcout(),
            .ltout(sDAC_data_RNO_8Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_3_LC_18_11_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_3_LC_18_11_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_3_LC_18_11_7.LUT_INIT=16'b0111011001010100;
    LogicCell40 sDAC_data_RNO_2_3_LC_18_11_7 (
            .in0(N__45099),
            .in1(N__45931),
            .in2(N__43011),
            .in3(N__43008),
            .lcout(sDAC_data_RNO_2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_3_7_LC_18_12_0.C_ON=1'b0;
    defparam sDAC_mem_3_7_LC_18_12_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_3_7_LC_18_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_3_7_LC_18_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48778),
            .lcout(sDAC_mem_3Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47709),
            .ce(N__42996),
            .sr(N__53055));
    defparam sDAC_data_RNO_28_10_LC_18_12_1.C_ON=1'b0;
    defparam sDAC_data_RNO_28_10_LC_18_12_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_28_10_LC_18_12_1.LUT_INIT=16'b0100011001010111;
    LogicCell40 sDAC_data_RNO_28_10_LC_18_12_1 (
            .in0(N__43674),
            .in1(N__52065),
            .in2(N__42906),
            .in3(N__42885),
            .lcout(),
            .ltout(sDAC_data_2_6_bm_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_15_10_LC_18_12_2.C_ON=1'b0;
    defparam sDAC_data_RNO_15_10_LC_18_12_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_15_10_LC_18_12_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 sDAC_data_RNO_15_10_LC_18_12_2 (
            .in0(N__52067),
            .in1(N__42870),
            .in2(N__42858),
            .in3(N__42855),
            .lcout(sDAC_data_RNO_15Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_16_4_LC_18_12_3.C_ON=1'b0;
    defparam sDAC_data_RNO_16_4_LC_18_12_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_16_4_LC_18_12_3.LUT_INIT=16'b0001110000011111;
    LogicCell40 sDAC_data_RNO_16_4_LC_18_12_3 (
            .in0(N__43716),
            .in1(N__52066),
            .in2(N__43687),
            .in3(N__43707),
            .lcout(),
            .ltout(sDAC_data_2_20_am_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_7_4_LC_18_12_4.C_ON=1'b0;
    defparam sDAC_data_RNO_7_4_LC_18_12_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_7_4_LC_18_12_4.LUT_INIT=16'b1100101000001111;
    LogicCell40 sDAC_data_RNO_7_4_LC_18_12_4 (
            .in0(N__43986),
            .in1(N__47205),
            .in2(N__43692),
            .in3(N__52139),
            .lcout(sDAC_data_RNO_7Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_17_4_LC_18_12_5.C_ON=1'b0;
    defparam sDAC_data_RNO_17_4_LC_18_12_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_17_4_LC_18_12_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_17_4_LC_18_12_5 (
            .in0(N__43678),
            .in1(N__44196),
            .in2(_gnd_net_),
            .in3(N__44331),
            .lcout(),
            .ltout(sDAC_data_RNO_17Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_8_4_LC_18_12_6.C_ON=1'b0;
    defparam sDAC_data_RNO_8_4_LC_18_12_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_8_4_LC_18_12_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 sDAC_data_RNO_8_4_LC_18_12_6 (
            .in0(_gnd_net_),
            .in1(N__52140),
            .in2(N__43311),
            .in3(N__45006),
            .lcout(),
            .ltout(sDAC_data_RNO_8Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_2_4_LC_18_12_7.C_ON=1'b0;
    defparam sDAC_data_RNO_2_4_LC_18_12_7.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_2_4_LC_18_12_7.LUT_INIT=16'b0111011001010100;
    LogicCell40 sDAC_data_RNO_2_4_LC_18_12_7 (
            .in0(N__45300),
            .in1(N__45889),
            .in2(N__43308),
            .in3(N__43305),
            .lcout(sDAC_data_RNO_2Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI5B15_2_1_LC_18_13_0.C_ON=1'b0;
    defparam sAddress_RNI5B15_2_1_LC_18_13_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI5B15_2_1_LC_18_13_0.LUT_INIT=16'b0011001100000000;
    LogicCell40 sAddress_RNI5B15_2_1_LC_18_13_0 (
            .in0(_gnd_net_),
            .in1(N__44896),
            .in2(_gnd_net_),
            .in3(N__44831),
            .lcout(N_284),
            .ltout(N_284_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_4_5_LC_18_13_1.C_ON=1'b0;
    defparam sAddress_RNI9IH12_4_5_LC_18_13_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_4_5_LC_18_13_1.LUT_INIT=16'b0000000000100000;
    LogicCell40 sAddress_RNI9IH12_4_5_LC_18_13_1 (
            .in0(N__46321),
            .in1(N__44445),
            .in2(N__43290),
            .in3(N__46569),
            .lcout(sDAC_mem_12_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_8_5_LC_18_13_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_8_5_LC_18_13_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_8_5_LC_18_13_2.LUT_INIT=16'b0000001000000000;
    LogicCell40 sAddress_RNI9IH12_8_5_LC_18_13_2 (
            .in0(N__43226),
            .in1(N__46119),
            .in2(N__46575),
            .in3(N__46320),
            .lcout(sDAC_mem_11_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_3_1_LC_18_13_3.C_ON=1'b0;
    defparam sAddress_RNI9IH12_3_1_LC_18_13_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_3_1_LC_18_13_3.LUT_INIT=16'b0100010000000000;
    LogicCell40 sAddress_RNI9IH12_3_1_LC_18_13_3 (
            .in0(N__46118),
            .in1(N__43225),
            .in2(_gnd_net_),
            .in3(N__43191),
            .lcout(sDAC_mem_27_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_1_LC_18_13_5.C_ON=1'b0;
    defparam sAddress_1_LC_18_13_5.SEQ_MODE=4'b1010;
    defparam sAddress_1_LC_18_13_5.LUT_INIT=16'b0000000011001100;
    LogicCell40 sAddress_1_LC_18_13_5 (
            .in0(_gnd_net_),
            .in1(N__50672),
            .in2(_gnd_net_),
            .in3(N__43868),
            .lcout(sAddressZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47715),
            .ce(N__43779),
            .sr(N__53045));
    defparam sAddress_RNI5B15_1_LC_18_13_6.C_ON=1'b0;
    defparam sAddress_RNI5B15_1_LC_18_13_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNI5B15_1_LC_18_13_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 sAddress_RNI5B15_1_LC_18_13_6 (
            .in0(_gnd_net_),
            .in1(N__44897),
            .in2(_gnd_net_),
            .in3(N__44832),
            .lcout(N_139),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_2_LC_18_13_7.C_ON=1'b0;
    defparam sAddress_2_LC_18_13_7.SEQ_MODE=4'b1010;
    defparam sAddress_2_LC_18_13_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 sAddress_2_LC_18_13_7 (
            .in0(_gnd_net_),
            .in1(N__50077),
            .in2(_gnd_net_),
            .in3(N__43869),
            .lcout(sAddressZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47715),
            .ce(N__43779),
            .sr(N__53045));
    defparam sDAC_mem_14_0_LC_18_14_0.C_ON=1'b0;
    defparam sDAC_mem_14_0_LC_18_14_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_0_LC_18_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_0_LC_18_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51268),
            .lcout(sDAC_mem_14Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47720),
            .ce(N__43935),
            .sr(N__53035));
    defparam sDAC_mem_14_1_LC_18_14_1.C_ON=1'b0;
    defparam sDAC_mem_14_1_LC_18_14_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_1_LC_18_14_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_1_LC_18_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50762),
            .lcout(sDAC_mem_14Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47720),
            .ce(N__43935),
            .sr(N__53035));
    defparam sDAC_mem_14_2_LC_18_14_2.C_ON=1'b0;
    defparam sDAC_mem_14_2_LC_18_14_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_2_LC_18_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_2_LC_18_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50090),
            .lcout(sDAC_mem_14Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47720),
            .ce(N__43935),
            .sr(N__53035));
    defparam sDAC_mem_14_3_LC_18_14_3.C_ON=1'b0;
    defparam sDAC_mem_14_3_LC_18_14_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_3_LC_18_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_3_LC_18_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49842),
            .lcout(sDAC_mem_14Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47720),
            .ce(N__43935),
            .sr(N__53035));
    defparam sDAC_mem_14_4_LC_18_14_4.C_ON=1'b0;
    defparam sDAC_mem_14_4_LC_18_14_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_4_LC_18_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_4_LC_18_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49308),
            .lcout(sDAC_mem_14Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47720),
            .ce(N__43935),
            .sr(N__53035));
    defparam sDAC_mem_14_5_LC_18_14_5.C_ON=1'b0;
    defparam sDAC_mem_14_5_LC_18_14_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_5_LC_18_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_5_LC_18_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47132),
            .lcout(sDAC_mem_14Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47720),
            .ce(N__43935),
            .sr(N__53035));
    defparam sDAC_mem_14_6_LC_18_14_6.C_ON=1'b0;
    defparam sDAC_mem_14_6_LC_18_14_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_6_LC_18_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_6_LC_18_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48340),
            .lcout(sDAC_mem_14Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47720),
            .ce(N__43935),
            .sr(N__53035));
    defparam sDAC_mem_14_7_LC_18_14_7.C_ON=1'b0;
    defparam sDAC_mem_14_7_LC_18_14_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_14_7_LC_18_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_14_7_LC_18_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48786),
            .lcout(sDAC_mem_14Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47720),
            .ce(N__43935),
            .sr(N__53035));
    defparam sDAC_data_RNO_19_7_LC_18_15_0.C_ON=1'b0;
    defparam sDAC_data_RNO_19_7_LC_18_15_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_7_LC_18_15_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_7_LC_18_15_0 (
            .in0(N__51973),
            .in1(N__45060),
            .in2(_gnd_net_),
            .in3(N__43929),
            .lcout(sDAC_data_RNO_19Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_7_LC_18_15_1.C_ON=1'b0;
    defparam sDAC_data_RNO_18_7_LC_18_15_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_7_LC_18_15_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_7_LC_18_15_1 (
            .in0(N__51983),
            .in1(N__48885),
            .in2(_gnd_net_),
            .in3(N__43887),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_7_LC_18_15_2.C_ON=1'b0;
    defparam sDAC_data_RNO_9_7_LC_18_15_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_7_LC_18_15_2.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_9_7_LC_18_15_2 (
            .in0(N__45890),
            .in1(N__45492),
            .in2(N__43923),
            .in3(N__43920),
            .lcout(sDAC_data_2_24_ns_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_8_LC_18_15_3.C_ON=1'b0;
    defparam sDAC_data_RNO_18_8_LC_18_15_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_8_LC_18_15_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_8_LC_18_15_3 (
            .in0(N__51984),
            .in1(N__45225),
            .in2(_gnd_net_),
            .in3(N__44148),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_8_LC_18_15_4.C_ON=1'b0;
    defparam sDAC_data_RNO_9_8_LC_18_15_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_8_LC_18_15_4.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_9_8_LC_18_15_4 (
            .in0(N__45891),
            .in1(N__45493),
            .in2(N__43899),
            .in3(N__43875),
            .lcout(sDAC_data_2_24_ns_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_12_4_LC_18_15_5.C_ON=1'b0;
    defparam sDAC_mem_12_4_LC_18_15_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_4_LC_18_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_4_LC_18_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49166),
            .lcout(sDAC_mem_12Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47730),
            .ce(N__47376),
            .sr(N__53026));
    defparam sDAC_data_RNO_19_8_LC_18_15_6.C_ON=1'b0;
    defparam sDAC_data_RNO_19_8_LC_18_15_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_8_LC_18_15_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_8_LC_18_15_6 (
            .in0(N__51974),
            .in1(N__45048),
            .in2(_gnd_net_),
            .in3(N__43881),
            .lcout(sDAC_data_RNO_19Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_12_5_LC_18_15_7.C_ON=1'b0;
    defparam sDAC_mem_12_5_LC_18_15_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_5_LC_18_15_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_5_LC_18_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47147),
            .lcout(sDAC_mem_12Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47730),
            .ce(N__47376),
            .sr(N__53026));
    defparam sEEADC_freq_1_LC_18_16_6.C_ON=1'b0;
    defparam sEEADC_freq_1_LC_18_16_6.SEQ_MODE=4'b1000;
    defparam sEEADC_freq_1_LC_18_16_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEADC_freq_1_LC_18_16_6 (
            .in0(N__50673),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEADC_freqZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47740),
            .ce(N__44126),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_29_3_LC_18_17_6.C_ON=1'b0;
    defparam sDAC_data_RNO_29_3_LC_18_17_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_29_3_LC_18_17_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 sDAC_data_RNO_29_3_LC_18_17_6 (
            .in0(N__44094),
            .in1(N__51890),
            .in2(_gnd_net_),
            .in3(N__44082),
            .lcout(sDAC_data_RNO_29Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_16_3_LC_18_19_0.C_ON=1'b0;
    defparam sDAC_mem_16_3_LC_18_19_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_3_LC_18_19_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_3_LC_18_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49845),
            .lcout(sDAC_mem_16Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47775),
            .ce(N__46631),
            .sr(N__52997));
    defparam sDAC_mem_20_7_LC_19_6_0.C_ON=1'b0;
    defparam sDAC_mem_20_7_LC_19_6_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_20_7_LC_19_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_20_7_LC_19_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48744),
            .lcout(sDAC_mem_20Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47731),
            .ce(N__44031),
            .sr(N__53135));
    defparam sDAC_mem_41_0_LC_19_7_0.C_ON=1'b0;
    defparam sDAC_mem_41_0_LC_19_7_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_0_LC_19_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_0_LC_19_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51239),
            .lcout(sDAC_mem_41Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47721),
            .ce(N__46263),
            .sr(N__53129));
    defparam sDAC_mem_41_1_LC_19_7_1.C_ON=1'b0;
    defparam sDAC_mem_41_1_LC_19_7_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_1_LC_19_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_1_LC_19_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50580),
            .lcout(sDAC_mem_41Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47721),
            .ce(N__46263),
            .sr(N__53129));
    defparam sDAC_mem_41_2_LC_19_7_2.C_ON=1'b0;
    defparam sDAC_mem_41_2_LC_19_7_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_2_LC_19_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_2_LC_19_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50230),
            .lcout(sDAC_mem_41Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47721),
            .ce(N__46263),
            .sr(N__53129));
    defparam sDAC_mem_41_3_LC_19_7_3.C_ON=1'b0;
    defparam sDAC_mem_41_3_LC_19_7_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_3_LC_19_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_3_LC_19_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49737),
            .lcout(sDAC_mem_41Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47721),
            .ce(N__46263),
            .sr(N__53129));
    defparam sDAC_mem_41_4_LC_19_7_4.C_ON=1'b0;
    defparam sDAC_mem_41_4_LC_19_7_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_4_LC_19_7_4.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_41_4_LC_19_7_4 (
            .in0(_gnd_net_),
            .in1(N__49281),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_41Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47721),
            .ce(N__46263),
            .sr(N__53129));
    defparam sDAC_mem_41_5_LC_19_7_5.C_ON=1'b0;
    defparam sDAC_mem_41_5_LC_19_7_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_5_LC_19_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_5_LC_19_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46984),
            .lcout(sDAC_mem_41Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47721),
            .ce(N__46263),
            .sr(N__53129));
    defparam sDAC_mem_41_6_LC_19_7_6.C_ON=1'b0;
    defparam sDAC_mem_41_6_LC_19_7_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_6_LC_19_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_6_LC_19_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48229),
            .lcout(sDAC_mem_41Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47721),
            .ce(N__46263),
            .sr(N__53129));
    defparam sDAC_mem_41_7_LC_19_7_7.C_ON=1'b0;
    defparam sDAC_mem_41_7_LC_19_7_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_41_7_LC_19_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_41_7_LC_19_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48745),
            .lcout(sDAC_mem_41Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47721),
            .ce(N__46263),
            .sr(N__53129));
    defparam sDAC_mem_42_0_LC_19_8_0.C_ON=1'b0;
    defparam sDAC_mem_42_0_LC_19_8_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_0_LC_19_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_42_0_LC_19_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51168),
            .lcout(sDAC_mem_42Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47716),
            .ce(N__44976),
            .sr(N__53115));
    defparam sDAC_mem_42_1_LC_19_8_1.C_ON=1'b0;
    defparam sDAC_mem_42_1_LC_19_8_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_1_LC_19_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_42_1_LC_19_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50581),
            .lcout(sDAC_mem_42Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47716),
            .ce(N__44976),
            .sr(N__53115));
    defparam sDAC_mem_42_2_LC_19_8_2.C_ON=1'b0;
    defparam sDAC_mem_42_2_LC_19_8_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_2_LC_19_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_42_2_LC_19_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50291),
            .lcout(sDAC_mem_42Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47716),
            .ce(N__44976),
            .sr(N__53115));
    defparam sDAC_mem_42_3_LC_19_8_3.C_ON=1'b0;
    defparam sDAC_mem_42_3_LC_19_8_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_3_LC_19_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_42_3_LC_19_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49825),
            .lcout(sDAC_mem_42Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47716),
            .ce(N__44976),
            .sr(N__53115));
    defparam sDAC_mem_42_4_LC_19_8_4.C_ON=1'b0;
    defparam sDAC_mem_42_4_LC_19_8_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_4_LC_19_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_42_4_LC_19_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49335),
            .lcout(sDAC_mem_42Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47716),
            .ce(N__44976),
            .sr(N__53115));
    defparam sDAC_mem_42_5_LC_19_8_5.C_ON=1'b0;
    defparam sDAC_mem_42_5_LC_19_8_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_5_LC_19_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_42_5_LC_19_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47137),
            .lcout(sDAC_mem_42Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47716),
            .ce(N__44976),
            .sr(N__53115));
    defparam sDAC_mem_42_6_LC_19_8_6.C_ON=1'b0;
    defparam sDAC_mem_42_6_LC_19_8_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_6_LC_19_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_42_6_LC_19_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48278),
            .lcout(sDAC_mem_42Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47716),
            .ce(N__44976),
            .sr(N__53115));
    defparam sDAC_mem_42_7_LC_19_8_7.C_ON=1'b0;
    defparam sDAC_mem_42_7_LC_19_8_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_42_7_LC_19_8_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_42_7_LC_19_8_7 (
            .in0(N__48833),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_42Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47716),
            .ce(N__44976),
            .sr(N__53115));
    defparam sDAC_mem_10_0_LC_19_9_0.C_ON=1'b0;
    defparam sDAC_mem_10_0_LC_19_9_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_0_LC_19_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_0_LC_19_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51240),
            .lcout(sDAC_mem_10Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47710),
            .ce(N__44993),
            .sr(N__53103));
    defparam sDAC_mem_10_1_LC_19_9_1.C_ON=1'b0;
    defparam sDAC_mem_10_1_LC_19_9_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_1_LC_19_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_1_LC_19_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50582),
            .lcout(sDAC_mem_10Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47710),
            .ce(N__44993),
            .sr(N__53103));
    defparam sDAC_mem_10_2_LC_19_9_2.C_ON=1'b0;
    defparam sDAC_mem_10_2_LC_19_9_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_2_LC_19_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_2_LC_19_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50286),
            .lcout(sDAC_mem_10Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47710),
            .ce(N__44993),
            .sr(N__53103));
    defparam sDAC_mem_10_3_LC_19_9_3.C_ON=1'b0;
    defparam sDAC_mem_10_3_LC_19_9_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_3_LC_19_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_3_LC_19_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49811),
            .lcout(sDAC_mem_10Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47710),
            .ce(N__44993),
            .sr(N__53103));
    defparam sDAC_mem_10_4_LC_19_9_4.C_ON=1'b0;
    defparam sDAC_mem_10_4_LC_19_9_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_4_LC_19_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_4_LC_19_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49336),
            .lcout(sDAC_mem_10Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47710),
            .ce(N__44993),
            .sr(N__53103));
    defparam sDAC_mem_10_5_LC_19_9_5.C_ON=1'b0;
    defparam sDAC_mem_10_5_LC_19_9_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_5_LC_19_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_5_LC_19_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47138),
            .lcout(sDAC_mem_10Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47710),
            .ce(N__44993),
            .sr(N__53103));
    defparam sDAC_mem_10_6_LC_19_9_6.C_ON=1'b0;
    defparam sDAC_mem_10_6_LC_19_9_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_10_6_LC_19_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_10_6_LC_19_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48279),
            .lcout(sDAC_mem_10Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47710),
            .ce(N__44993),
            .sr(N__53103));
    defparam sAddress_RNI9IH12_10_5_LC_19_10_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_10_5_LC_19_10_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_10_5_LC_19_10_0.LUT_INIT=16'b0000000000000010;
    LogicCell40 sAddress_RNI9IH12_10_5_LC_19_10_0 (
            .in0(N__46294),
            .in1(N__46413),
            .in2(N__44470),
            .in3(N__46563),
            .lcout(sDAC_mem_10_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_6_5_LC_19_10_1.C_ON=1'b0;
    defparam sAddress_RNI9IH12_6_5_LC_19_10_1.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_6_5_LC_19_10_1.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNI9IH12_6_5_LC_19_10_1 (
            .in0(N__46566),
            .in1(N__46123),
            .in2(N__44554),
            .in3(N__46292),
            .lcout(sDAC_mem_15_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_5_5_LC_19_10_2.C_ON=1'b0;
    defparam sAddress_RNI9IH12_5_5_LC_19_10_2.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_5_5_LC_19_10_2.LUT_INIT=16'b0000001000000000;
    LogicCell40 sAddress_RNI9IH12_5_5_LC_19_10_2 (
            .in0(N__46295),
            .in1(N__46414),
            .in2(N__44471),
            .in3(N__46564),
            .lcout(sDAC_mem_42_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI5B15_0_1_LC_19_10_3.C_ON=1'b0;
    defparam sAddress_RNI5B15_0_1_LC_19_10_3.SEQ_MODE=4'b0000;
    defparam sAddress_RNI5B15_0_1_LC_19_10_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 sAddress_RNI5B15_0_1_LC_19_10_3 (
            .in0(_gnd_net_),
            .in1(N__44931),
            .in2(_gnd_net_),
            .in3(N__44855),
            .lcout(N_286),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNIP2UK1_4_LC_19_10_4.C_ON=1'b0;
    defparam sAddress_RNIP2UK1_4_LC_19_10_4.SEQ_MODE=4'b0000;
    defparam sAddress_RNIP2UK1_4_LC_19_10_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 sAddress_RNIP2UK1_4_LC_19_10_4 (
            .in0(N__44778),
            .in1(N__44722),
            .in2(_gnd_net_),
            .in3(N__44636),
            .lcout(N_278),
            .ltout(N_278_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_2_5_LC_19_10_5.C_ON=1'b0;
    defparam sAddress_RNI9IH12_2_5_LC_19_10_5.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_2_5_LC_19_10_5.LUT_INIT=16'b0000000001000000;
    LogicCell40 sAddress_RNI9IH12_2_5_LC_19_10_5 (
            .in0(N__46565),
            .in1(N__44539),
            .in2(N__44481),
            .in3(N__44459),
            .lcout(sDAC_mem_16_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_9_5_LC_19_10_6.C_ON=1'b0;
    defparam sAddress_RNI9IH12_9_5_LC_19_10_6.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_9_5_LC_19_10_6.LUT_INIT=16'b0000000000000010;
    LogicCell40 sAddress_RNI9IH12_9_5_LC_19_10_6 (
            .in0(N__46296),
            .in1(N__46412),
            .in2(N__46133),
            .in3(N__46568),
            .lcout(sDAC_mem_9_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_7_5_LC_19_10_7.C_ON=1'b0;
    defparam sAddress_RNI9IH12_7_5_LC_19_10_7.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_7_5_LC_19_10_7.LUT_INIT=16'b0001000000000000;
    LogicCell40 sAddress_RNI9IH12_7_5_LC_19_10_7 (
            .in0(N__46567),
            .in1(N__46124),
            .in2(N__46247),
            .in3(N__46293),
            .lcout(sDAC_mem_13_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_15_0_LC_19_11_0.C_ON=1'b0;
    defparam sDAC_mem_15_0_LC_19_11_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_0_LC_19_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_0_LC_19_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51241),
            .lcout(sDAC_mem_15Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47702),
            .ce(N__45024),
            .sr(N__53077));
    defparam sDAC_mem_15_1_LC_19_11_1.C_ON=1'b0;
    defparam sDAC_mem_15_1_LC_19_11_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_1_LC_19_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_1_LC_19_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50583),
            .lcout(sDAC_mem_15Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47702),
            .ce(N__45024),
            .sr(N__53077));
    defparam sDAC_mem_15_2_LC_19_11_2.C_ON=1'b0;
    defparam sDAC_mem_15_2_LC_19_11_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_2_LC_19_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_2_LC_19_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50287),
            .lcout(sDAC_mem_15Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47702),
            .ce(N__45024),
            .sr(N__53077));
    defparam sDAC_mem_15_3_LC_19_11_3.C_ON=1'b0;
    defparam sDAC_mem_15_3_LC_19_11_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_3_LC_19_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_3_LC_19_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49819),
            .lcout(sDAC_mem_15Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47702),
            .ce(N__45024),
            .sr(N__53077));
    defparam sDAC_mem_15_4_LC_19_11_4.C_ON=1'b0;
    defparam sDAC_mem_15_4_LC_19_11_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_4_LC_19_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_4_LC_19_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49359),
            .lcout(sDAC_mem_15Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47702),
            .ce(N__45024),
            .sr(N__53077));
    defparam sDAC_mem_15_5_LC_19_11_5.C_ON=1'b0;
    defparam sDAC_mem_15_5_LC_19_11_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_5_LC_19_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_5_LC_19_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47150),
            .lcout(sDAC_mem_15Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47702),
            .ce(N__45024),
            .sr(N__53077));
    defparam sDAC_mem_15_6_LC_19_11_6.C_ON=1'b0;
    defparam sDAC_mem_15_6_LC_19_11_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_6_LC_19_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_6_LC_19_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48330),
            .lcout(sDAC_mem_15Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47702),
            .ce(N__45024),
            .sr(N__53077));
    defparam sDAC_mem_15_7_LC_19_11_7.C_ON=1'b0;
    defparam sDAC_mem_15_7_LC_19_11_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_15_7_LC_19_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_15_7_LC_19_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48812),
            .lcout(sDAC_mem_15Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47702),
            .ce(N__45024),
            .sr(N__53077));
    defparam sDAC_mem_11_0_LC_19_12_0.C_ON=1'b0;
    defparam sDAC_mem_11_0_LC_19_12_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_0_LC_19_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_0_LC_19_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51242),
            .lcout(sDAC_mem_11Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47705),
            .ce(N__45129),
            .sr(N__53066));
    defparam sDAC_mem_11_1_LC_19_12_1.C_ON=1'b0;
    defparam sDAC_mem_11_1_LC_19_12_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_1_LC_19_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_1_LC_19_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50584),
            .lcout(sDAC_mem_11Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47705),
            .ce(N__45129),
            .sr(N__53066));
    defparam sDAC_mem_11_2_LC_19_12_2.C_ON=1'b0;
    defparam sDAC_mem_11_2_LC_19_12_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_2_LC_19_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_2_LC_19_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50307),
            .lcout(sDAC_mem_11Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47705),
            .ce(N__45129),
            .sr(N__53066));
    defparam sDAC_mem_11_3_LC_19_12_3.C_ON=1'b0;
    defparam sDAC_mem_11_3_LC_19_12_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_3_LC_19_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_3_LC_19_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49841),
            .lcout(sDAC_mem_11Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47705),
            .ce(N__45129),
            .sr(N__53066));
    defparam sDAC_mem_11_4_LC_19_12_4.C_ON=1'b0;
    defparam sDAC_mem_11_4_LC_19_12_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_4_LC_19_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_4_LC_19_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49322),
            .lcout(sDAC_mem_11Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47705),
            .ce(N__45129),
            .sr(N__53066));
    defparam sDAC_mem_11_5_LC_19_12_5.C_ON=1'b0;
    defparam sDAC_mem_11_5_LC_19_12_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_5_LC_19_12_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_5_LC_19_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47151),
            .lcout(sDAC_mem_11Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47705),
            .ce(N__45129),
            .sr(N__53066));
    defparam sDAC_mem_11_6_LC_19_12_6.C_ON=1'b0;
    defparam sDAC_mem_11_6_LC_19_12_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_6_LC_19_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_11_6_LC_19_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48325),
            .lcout(sDAC_mem_11Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47705),
            .ce(N__45129),
            .sr(N__53066));
    defparam sDAC_mem_11_7_LC_19_12_7.C_ON=1'b0;
    defparam sDAC_mem_11_7_LC_19_12_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_11_7_LC_19_12_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_11_7_LC_19_12_7 (
            .in0(N__48779),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_11Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47705),
            .ce(N__45129),
            .sr(N__53066));
    defparam sDAC_data_RNO_19_3_LC_19_13_0.C_ON=1'b0;
    defparam sDAC_data_RNO_19_3_LC_19_13_0.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_3_LC_19_13_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_3_LC_19_13_0 (
            .in0(N__52146),
            .in1(N__45123),
            .in2(_gnd_net_),
            .in3(N__45114),
            .lcout(sDAC_data_RNO_19Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_3_LC_19_13_1.C_ON=1'b0;
    defparam sDAC_data_RNO_18_3_LC_19_13_1.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_3_LC_19_13_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_3_LC_19_13_1 (
            .in0(N__52148),
            .in1(N__50778),
            .in2(_gnd_net_),
            .in3(N__45294),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_3_LC_19_13_2.C_ON=1'b0;
    defparam sDAC_data_RNO_9_3_LC_19_13_2.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_3_LC_19_13_2.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_9_3_LC_19_13_2 (
            .in0(N__45910),
            .in1(N__45494),
            .in2(N__45108),
            .in3(N__45105),
            .lcout(sDAC_data_2_24_ns_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_4_LC_19_13_3.C_ON=1'b0;
    defparam sDAC_data_RNO_18_4_LC_19_13_3.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_4_LC_19_13_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_4_LC_19_13_3 (
            .in0(N__52149),
            .in1(N__50316),
            .in2(_gnd_net_),
            .in3(N__45267),
            .lcout(),
            .ltout(sDAC_data_RNO_18Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_9_4_LC_19_13_4.C_ON=1'b0;
    defparam sDAC_data_RNO_9_4_LC_19_13_4.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_9_4_LC_19_13_4.LUT_INIT=16'b0001001110011011;
    LogicCell40 sDAC_data_RNO_9_4_LC_19_13_4 (
            .in0(N__45911),
            .in1(N__45495),
            .in2(N__45303),
            .in3(N__45273),
            .lcout(sDAC_data_2_24_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_12_0_LC_19_13_5.C_ON=1'b0;
    defparam sDAC_mem_12_0_LC_19_13_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_0_LC_19_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_0_LC_19_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51270),
            .lcout(sDAC_mem_12Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47711),
            .ce(N__47375),
            .sr(N__53056));
    defparam sDAC_data_RNO_19_4_LC_19_13_6.C_ON=1'b0;
    defparam sDAC_data_RNO_19_4_LC_19_13_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_4_LC_19_13_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_4_LC_19_13_6 (
            .in0(N__52147),
            .in1(N__45288),
            .in2(_gnd_net_),
            .in3(N__45279),
            .lcout(sDAC_data_RNO_19Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_12_1_LC_19_13_7.C_ON=1'b0;
    defparam sDAC_mem_12_1_LC_19_13_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_1_LC_19_13_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_1_LC_19_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50585),
            .lcout(sDAC_mem_12Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47711),
            .ce(N__47375),
            .sr(N__53056));
    defparam sDAC_mem_27_0_LC_19_14_0.C_ON=1'b0;
    defparam sDAC_mem_27_0_LC_19_14_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_27_0_LC_19_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_27_0_LC_19_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51081),
            .lcout(sDAC_mem_27Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47717),
            .ce(N__45246),
            .sr(N__53046));
    defparam sDAC_mem_13_6_LC_19_15_4.C_ON=1'b0;
    defparam sDAC_mem_13_6_LC_19_15_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_6_LC_19_15_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_6_LC_19_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48232),
            .lcout(sDAC_mem_13Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47722),
            .ce(N__48867),
            .sr(N__53036));
    defparam sDAC_mem_13_5_LC_19_15_6.C_ON=1'b0;
    defparam sDAC_mem_13_5_LC_19_15_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_5_LC_19_15_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_5_LC_19_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47148),
            .lcout(sDAC_mem_13Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47722),
            .ce(N__48867),
            .sr(N__53036));
    defparam sDAC_mem_16_1_LC_19_18_0.C_ON=1'b0;
    defparam sDAC_mem_16_1_LC_19_18_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_16_1_LC_19_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_16_1_LC_19_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50674),
            .lcout(sDAC_mem_16Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47753),
            .ce(N__46630),
            .sr(N__53015));
    defparam sEEDAC_7_LC_20_5_0.C_ON=1'b0;
    defparam sEEDAC_7_LC_20_5_0.SEQ_MODE=4'b1000;
    defparam sEEDAC_7_LC_20_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_7_LC_20_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48729),
            .lcout(sEEDACZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47732),
            .ce(N__47238),
            .sr(_gnd_net_));
    defparam sAddress_RNI9IH12_1_5_LC_20_7_0.C_ON=1'b0;
    defparam sAddress_RNI9IH12_1_5_LC_20_7_0.SEQ_MODE=4'b0000;
    defparam sAddress_RNI9IH12_1_5_LC_20_7_0.LUT_INIT=16'b0000001000000000;
    LogicCell40 sAddress_RNI9IH12_1_5_LC_20_7_0 (
            .in0(N__46559),
            .in1(N__46134),
            .in2(N__46445),
            .in3(N__46319),
            .lcout(sDAC_mem_41_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam reset_rpi_ibuf_RNIRGF52_0_LC_20_8_0.C_ON=1'b0;
    defparam reset_rpi_ibuf_RNIRGF52_0_LC_20_8_0.SEQ_MODE=4'b0000;
    defparam reset_rpi_ibuf_RNIRGF52_0_LC_20_8_0.LUT_INIT=16'b0010001000000000;
    LogicCell40 reset_rpi_ibuf_RNIRGF52_0_LC_20_8_0 (
            .in0(N__46248),
            .in1(N__46128),
            .in2(_gnd_net_),
            .in3(N__46043),
            .lcout(sEEDAC_1_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sEEDAC_0_LC_20_8_1.C_ON=1'b0;
    defparam sEEDAC_0_LC_20_8_1.SEQ_MODE=4'b1000;
    defparam sEEDAC_0_LC_20_8_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEDAC_0_LC_20_8_1 (
            .in0(N__51181),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEDACZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47712),
            .ce(N__47234),
            .sr(_gnd_net_));
    defparam sEEDAC_1_LC_20_8_2.C_ON=1'b0;
    defparam sEEDAC_1_LC_20_8_2.SEQ_MODE=4'b1000;
    defparam sEEDAC_1_LC_20_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_1_LC_20_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50725),
            .lcout(sEEDACZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47712),
            .ce(N__47234),
            .sr(_gnd_net_));
    defparam sEEDAC_2_LC_20_8_3.C_ON=1'b0;
    defparam sEEDAC_2_LC_20_8_3.SEQ_MODE=4'b1000;
    defparam sEEDAC_2_LC_20_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_2_LC_20_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50292),
            .lcout(sEEDACZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47712),
            .ce(N__47234),
            .sr(_gnd_net_));
    defparam sEEDAC_3_LC_20_8_4.C_ON=1'b0;
    defparam sEEDAC_3_LC_20_8_4.SEQ_MODE=4'b1000;
    defparam sEEDAC_3_LC_20_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_3_LC_20_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49826),
            .lcout(sEEDACZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47712),
            .ce(N__47234),
            .sr(_gnd_net_));
    defparam sEEDAC_4_LC_20_8_5.C_ON=1'b0;
    defparam sEEDAC_4_LC_20_8_5.SEQ_MODE=4'b1000;
    defparam sEEDAC_4_LC_20_8_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 sEEDAC_4_LC_20_8_5 (
            .in0(N__49343),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sEEDACZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47712),
            .ce(N__47234),
            .sr(_gnd_net_));
    defparam sEEDAC_5_LC_20_8_6.C_ON=1'b0;
    defparam sEEDAC_5_LC_20_8_6.SEQ_MODE=4'b1000;
    defparam sEEDAC_5_LC_20_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_5_LC_20_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47139),
            .lcout(sEEDACZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47712),
            .ce(N__47234),
            .sr(_gnd_net_));
    defparam sEEDAC_6_LC_20_8_7.C_ON=1'b0;
    defparam sEEDAC_6_LC_20_8_7.SEQ_MODE=4'b1000;
    defparam sEEDAC_6_LC_20_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sEEDAC_6_LC_20_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48280),
            .lcout(sEEDACZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47712),
            .ce(N__47234),
            .sr(_gnd_net_));
    defparam sDAC_mem_9_0_LC_20_9_0.C_ON=1'b0;
    defparam sDAC_mem_9_0_LC_20_9_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_0_LC_20_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_9_0_LC_20_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50981),
            .lcout(sDAC_mem_9Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47706),
            .ce(N__47325),
            .sr(N__53116));
    defparam sDAC_mem_9_1_LC_20_9_1.C_ON=1'b0;
    defparam sDAC_mem_9_1_LC_20_9_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_1_LC_20_9_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_9_1_LC_20_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50753),
            .lcout(sDAC_mem_9Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47706),
            .ce(N__47325),
            .sr(N__53116));
    defparam sDAC_mem_9_2_LC_20_9_2.C_ON=1'b0;
    defparam sDAC_mem_9_2_LC_20_9_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_2_LC_20_9_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_9_2_LC_20_9_2 (
            .in0(N__50308),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_9Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47706),
            .ce(N__47325),
            .sr(N__53116));
    defparam sDAC_mem_9_3_LC_20_9_3.C_ON=1'b0;
    defparam sDAC_mem_9_3_LC_20_9_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_3_LC_20_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_9_3_LC_20_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49843),
            .lcout(sDAC_mem_9Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47706),
            .ce(N__47325),
            .sr(N__53116));
    defparam sDAC_mem_9_4_LC_20_9_4.C_ON=1'b0;
    defparam sDAC_mem_9_4_LC_20_9_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_4_LC_20_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_9_4_LC_20_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49344),
            .lcout(sDAC_mem_9Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47706),
            .ce(N__47325),
            .sr(N__53116));
    defparam sDAC_mem_9_5_LC_20_9_5.C_ON=1'b0;
    defparam sDAC_mem_9_5_LC_20_9_5.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_5_LC_20_9_5.LUT_INIT=16'b1100110011001100;
    LogicCell40 sDAC_mem_9_5_LC_20_9_5 (
            .in0(_gnd_net_),
            .in1(N__47140),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_9Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47706),
            .ce(N__47325),
            .sr(N__53116));
    defparam sDAC_mem_9_6_LC_20_9_6.C_ON=1'b0;
    defparam sDAC_mem_9_6_LC_20_9_6.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_6_LC_20_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_9_6_LC_20_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48281),
            .lcout(sDAC_mem_9Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47706),
            .ce(N__47325),
            .sr(N__53116));
    defparam sDAC_mem_9_7_LC_20_9_7.C_ON=1'b0;
    defparam sDAC_mem_9_7_LC_20_9_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_9_7_LC_20_9_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_9_7_LC_20_9_7 (
            .in0(N__48718),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_9Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47706),
            .ce(N__47325),
            .sr(N__53116));
    defparam sCounterDAC_6_LC_20_10_0.C_ON=1'b0;
    defparam sCounterDAC_6_LC_20_10_0.SEQ_MODE=4'b1010;
    defparam sCounterDAC_6_LC_20_10_0.LUT_INIT=16'b0000011001100110;
    LogicCell40 sCounterDAC_6_LC_20_10_0 (
            .in0(N__52176),
            .in1(N__52444),
            .in2(N__52253),
            .in3(N__53449),
            .lcout(sCounterDACZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53274),
            .ce(),
            .sr(N__53104));
    defparam sCounterDAC_RNI7A77_1_LC_20_10_5.C_ON=1'b0;
    defparam sCounterDAC_RNI7A77_1_LC_20_10_5.SEQ_MODE=4'b0000;
    defparam sCounterDAC_RNI7A77_1_LC_20_10_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 sCounterDAC_RNI7A77_1_LC_20_10_5 (
            .in0(N__52547),
            .in1(N__53357),
            .in2(N__53414),
            .in3(N__52524),
            .lcout(N_14_3),
            .ltout(N_14_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_spi_start_RNO_0_LC_20_10_6.C_ON=1'b0;
    defparam sDAC_spi_start_RNO_0_LC_20_10_6.SEQ_MODE=4'b0000;
    defparam sDAC_spi_start_RNO_0_LC_20_10_6.LUT_INIT=16'b1111000011110010;
    LogicCell40 sDAC_spi_start_RNO_0_LC_20_10_6 (
            .in0(N__47286),
            .in1(N__52548),
            .in2(N__47313),
            .in3(N__52232),
            .lcout(),
            .ltout(N_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_spi_start_LC_20_10_7.C_ON=1'b0;
    defparam sDAC_spi_start_LC_20_10_7.SEQ_MODE=4'b1010;
    defparam sDAC_spi_start_LC_20_10_7.LUT_INIT=16'b1110101000101010;
    LogicCell40 sDAC_spi_start_LC_20_10_7 (
            .in0(N__47300),
            .in1(N__47280),
            .in2(N__47310),
            .in3(N__53337),
            .lcout(sDAC_spi_startZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53274),
            .ce(),
            .sr(N__53104));
    defparam sCounterDAC_RNIPQJ3_3_LC_20_11_0.C_ON=1'b0;
    defparam sCounterDAC_RNIPQJ3_3_LC_20_11_0.SEQ_MODE=4'b0000;
    defparam sCounterDAC_RNIPQJ3_3_LC_20_11_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 sCounterDAC_RNIPQJ3_3_LC_20_11_0 (
            .in0(N__53335),
            .in1(N__52199),
            .in2(_gnd_net_),
            .in3(N__52233),
            .lcout(N_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_spi_start_RNO_2_LC_20_11_1.C_ON=1'b0;
    defparam sDAC_spi_start_RNO_2_LC_20_11_1.SEQ_MODE=4'b0000;
    defparam sDAC_spi_start_RNO_2_LC_20_11_1.LUT_INIT=16'b0000000000010001;
    LogicCell40 sDAC_spi_start_RNO_2_LC_20_11_1 (
            .in0(N__52200),
            .in1(N__52520),
            .in2(_gnd_net_),
            .in3(N__53336),
            .lcout(un1_scounterdac8_i_a2_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_spi_start_RNO_1_LC_20_11_3.C_ON=1'b0;
    defparam sDAC_spi_start_RNO_1_LC_20_11_3.SEQ_MODE=4'b0000;
    defparam sDAC_spi_start_RNO_1_LC_20_11_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 sDAC_spi_start_RNO_1_LC_20_11_3 (
            .in0(N__53410),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53451),
            .lcout(un1_scounterdac8_i_a2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_18_10_LC_20_11_5.C_ON=1'b0;
    defparam sDAC_data_RNO_18_10_LC_20_11_5.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_18_10_LC_20_11_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_18_10_LC_20_11_5 (
            .in0(N__52077),
            .in1(N__48873),
            .in2(_gnd_net_),
            .in3(N__48351),
            .lcout(sDAC_data_RNO_18Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_data_RNO_19_10_LC_20_11_6.C_ON=1'b0;
    defparam sDAC_data_RNO_19_10_LC_20_11_6.SEQ_MODE=4'b0000;
    defparam sDAC_data_RNO_19_10_LC_20_11_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 sDAC_data_RNO_19_10_LC_20_11_6 (
            .in0(N__52076),
            .in1(N__51306),
            .in2(_gnd_net_),
            .in3(N__51300),
            .lcout(sDAC_data_RNO_19Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sDAC_mem_13_0_LC_20_12_0.C_ON=1'b0;
    defparam sDAC_mem_13_0_LC_20_12_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_0_LC_20_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_0_LC_20_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50982),
            .lcout(sDAC_mem_13Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47703),
            .ce(N__48866),
            .sr(N__53078));
    defparam sDAC_mem_13_1_LC_20_12_1.C_ON=1'b0;
    defparam sDAC_mem_13_1_LC_20_12_1.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_1_LC_20_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_1_LC_20_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50576),
            .lcout(sDAC_mem_13Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47703),
            .ce(N__48866),
            .sr(N__53078));
    defparam sDAC_mem_13_2_LC_20_12_2.C_ON=1'b0;
    defparam sDAC_mem_13_2_LC_20_12_2.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_2_LC_20_12_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_13_2_LC_20_12_2 (
            .in0(N__50309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_13Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47703),
            .ce(N__48866),
            .sr(N__53078));
    defparam sDAC_mem_13_3_LC_20_12_3.C_ON=1'b0;
    defparam sDAC_mem_13_3_LC_20_12_3.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_3_LC_20_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_3_LC_20_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49844),
            .lcout(sDAC_mem_13Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47703),
            .ce(N__48866),
            .sr(N__53078));
    defparam sDAC_mem_13_4_LC_20_12_4.C_ON=1'b0;
    defparam sDAC_mem_13_4_LC_20_12_4.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_4_LC_20_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_4_LC_20_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49355),
            .lcout(sDAC_mem_13Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47703),
            .ce(N__48866),
            .sr(N__53078));
    defparam sDAC_mem_13_7_LC_20_12_7.C_ON=1'b0;
    defparam sDAC_mem_13_7_LC_20_12_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_13_7_LC_20_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_13_7_LC_20_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48719),
            .lcout(sDAC_mem_13Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47703),
            .ce(N__48866),
            .sr(N__53078));
    defparam sDAC_mem_12_7_LC_20_13_0.C_ON=1'b0;
    defparam sDAC_mem_12_7_LC_20_13_0.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_7_LC_20_13_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 sDAC_mem_12_7_LC_20_13_0 (
            .in0(N__48728),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(sDAC_mem_12Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47707),
            .ce(N__47377),
            .sr(N__53067));
    defparam sDAC_mem_12_6_LC_20_16_7.C_ON=1'b0;
    defparam sDAC_mem_12_6_LC_20_16_7.SEQ_MODE=4'b1010;
    defparam sDAC_mem_12_6_LC_20_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 sDAC_mem_12_6_LC_20_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48341),
            .lcout(sDAC_mem_12Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47723),
            .ce(N__47391),
            .sr(N__53037));
    defparam sCounterDAC_8_LC_22_8_2.C_ON=1'b0;
    defparam sCounterDAC_8_LC_22_8_2.SEQ_MODE=4'b1010;
    defparam sCounterDAC_8_LC_22_8_2.LUT_INIT=16'b0001010100101010;
    LogicCell40 sCounterDAC_8_LC_22_8_2 (
            .in0(N__53298),
            .in1(N__53450),
            .in2(N__52260),
            .in3(N__53322),
            .lcout(sCounterDACZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53275),
            .ce(),
            .sr(N__53140));
    defparam un2_scounterdac_cry_1_c_LC_22_10_0.C_ON=1'b1;
    defparam un2_scounterdac_cry_1_c_LC_22_10_0.SEQ_MODE=4'b0000;
    defparam un2_scounterdac_cry_1_c_LC_22_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_scounterdac_cry_1_c_LC_22_10_0 (
            .in0(_gnd_net_),
            .in1(N__52512),
            .in2(N__53395),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_22_10_0_),
            .carryout(un2_scounterdac_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_2_LC_22_10_1.C_ON=1'b1;
    defparam sCounterDAC_2_LC_22_10_1.SEQ_MODE=4'b1010;
    defparam sCounterDAC_2_LC_22_10_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 sCounterDAC_2_LC_22_10_1 (
            .in0(_gnd_net_),
            .in1(N__52476),
            .in2(_gnd_net_),
            .in3(N__52236),
            .lcout(sCounterDACZ0Z_2),
            .ltout(),
            .carryin(un2_scounterdac_cry_1),
            .carryout(un2_scounterdac_cry_2),
            .clk(N__53277),
            .ce(),
            .sr(N__53130));
    defparam sCounterDAC_3_LC_22_10_2.C_ON=1'b1;
    defparam sCounterDAC_3_LC_22_10_2.SEQ_MODE=4'b1010;
    defparam sCounterDAC_3_LC_22_10_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 sCounterDAC_3_LC_22_10_2 (
            .in0(_gnd_net_),
            .in1(N__52225),
            .in2(_gnd_net_),
            .in3(N__52206),
            .lcout(sCounterDACZ0Z_3),
            .ltout(),
            .carryin(un2_scounterdac_cry_2),
            .carryout(un2_scounterdac_cry_3),
            .clk(N__53277),
            .ce(),
            .sr(N__53130));
    defparam sCounterDAC_4_LC_22_10_3.C_ON=1'b1;
    defparam sCounterDAC_4_LC_22_10_3.SEQ_MODE=4'b1010;
    defparam sCounterDAC_4_LC_22_10_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 sCounterDAC_4_LC_22_10_3 (
            .in0(_gnd_net_),
            .in1(N__52541),
            .in2(_gnd_net_),
            .in3(N__52203),
            .lcout(sCounterDACZ0Z_4),
            .ltout(),
            .carryin(un2_scounterdac_cry_3),
            .carryout(un2_scounterdac_cry_4),
            .clk(N__53277),
            .ce(),
            .sr(N__53130));
    defparam sCounterDAC_5_LC_22_10_4.C_ON=1'b1;
    defparam sCounterDAC_5_LC_22_10_4.SEQ_MODE=4'b1010;
    defparam sCounterDAC_5_LC_22_10_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 sCounterDAC_5_LC_22_10_4 (
            .in0(_gnd_net_),
            .in1(N__52193),
            .in2(_gnd_net_),
            .in3(N__52179),
            .lcout(sCounterDACZ0Z_5),
            .ltout(),
            .carryin(un2_scounterdac_cry_4),
            .carryout(un2_scounterdac_cry_5),
            .clk(N__53277),
            .ce(),
            .sr(N__53130));
    defparam un2_scounterdac_cry_5_THRU_LUT4_0_LC_22_10_5.C_ON=1'b1;
    defparam un2_scounterdac_cry_5_THRU_LUT4_0_LC_22_10_5.SEQ_MODE=4'b0000;
    defparam un2_scounterdac_cry_5_THRU_LUT4_0_LC_22_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_scounterdac_cry_5_THRU_LUT4_0_LC_22_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52449),
            .in3(N__52167),
            .lcout(un2_scounterdac_cry_5_THRU_CO),
            .ltout(),
            .carryin(un2_scounterdac_cry_5),
            .carryout(un2_scounterdac_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_7_LC_22_10_6.C_ON=1'b1;
    defparam sCounterDAC_7_LC_22_10_6.SEQ_MODE=4'b1010;
    defparam sCounterDAC_7_LC_22_10_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 sCounterDAC_7_LC_22_10_6 (
            .in0(_gnd_net_),
            .in1(N__52488),
            .in2(_gnd_net_),
            .in3(N__52164),
            .lcout(sCounterDACZ0Z_7),
            .ltout(),
            .carryin(un2_scounterdac_cry_6),
            .carryout(un2_scounterdac_cry_7),
            .clk(N__53277),
            .ce(),
            .sr(N__53130));
    defparam un2_scounterdac_cry_7_THRU_LUT4_0_LC_22_10_7.C_ON=1'b1;
    defparam un2_scounterdac_cry_7_THRU_LUT4_0_LC_22_10_7.SEQ_MODE=4'b0000;
    defparam un2_scounterdac_cry_7_THRU_LUT4_0_LC_22_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_scounterdac_cry_7_THRU_LUT4_0_LC_22_10_7 (
            .in0(_gnd_net_),
            .in1(N__53331),
            .in2(_gnd_net_),
            .in3(N__53289),
            .lcout(un2_scounterdac_cry_7_THRU_CO),
            .ltout(),
            .carryin(un2_scounterdac_cry_7),
            .carryout(un2_scounterdac_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_9_LC_22_11_0.C_ON=1'b0;
    defparam sCounterDAC_9_LC_22_11_0.SEQ_MODE=4'b1010;
    defparam sCounterDAC_9_LC_22_11_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 sCounterDAC_9_LC_22_11_0 (
            .in0(_gnd_net_),
            .in1(N__52463),
            .in2(_gnd_net_),
            .in3(N__53286),
            .lcout(sCounterDACZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53279),
            .ce(),
            .sr(N__53117));
    defparam sCounterDAC_0_LC_22_11_1.C_ON=1'b0;
    defparam sCounterDAC_0_LC_22_11_1.SEQ_MODE=4'b1010;
    defparam sCounterDAC_0_LC_22_11_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 sCounterDAC_0_LC_22_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53405),
            .lcout(sCounterDACZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53279),
            .ce(),
            .sr(N__53117));
    defparam sCounterDAC_1_LC_22_11_7.C_ON=1'b0;
    defparam sCounterDAC_1_LC_22_11_7.SEQ_MODE=4'b1010;
    defparam sCounterDAC_1_LC_22_11_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 sCounterDAC_1_LC_22_11_7 (
            .in0(_gnd_net_),
            .in1(N__53406),
            .in2(_gnd_net_),
            .in3(N__52519),
            .lcout(sCounterDACZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__53279),
            .ce(),
            .sr(N__53117));
    defparam \spi_slave_inst.spi_mosi_flash_LC_23_1_2 .C_ON=1'b0;
    defparam \spi_slave_inst.spi_mosi_flash_LC_23_1_2 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.spi_mosi_flash_LC_23_1_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \spi_slave_inst.spi_mosi_flash_LC_23_1_2  (
            .in0(N__52304),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52596),
            .lcout(spi_mosi_flash_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_RNIB1D2_1_LC_23_10_2.C_ON=1'b0;
    defparam sCounterDAC_RNIB1D2_1_LC_23_10_2.SEQ_MODE=4'b0000;
    defparam sCounterDAC_RNIB1D2_1_LC_23_10_2.LUT_INIT=16'b0000000000110011;
    LogicCell40 sCounterDAC_RNIB1D2_1_LC_23_10_2 (
            .in0(_gnd_net_),
            .in1(N__52540),
            .in2(_gnd_net_),
            .in3(N__52511),
            .lcout(op_eq_scounterdac10_0_a2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_RNI4HQ4_9_LC_23_10_4.C_ON=1'b0;
    defparam sCounterDAC_RNI4HQ4_9_LC_23_10_4.SEQ_MODE=4'b0000;
    defparam sCounterDAC_RNI4HQ4_9_LC_23_10_4.LUT_INIT=16'b0000000000000100;
    LogicCell40 sCounterDAC_RNI4HQ4_9_LC_23_10_4 (
            .in0(N__52487),
            .in1(N__52475),
            .in2(N__52464),
            .in3(N__52445),
            .lcout(N_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.spi_cs_flash_LC_24_1_1 .C_ON=1'b0;
    defparam \spi_slave_inst.spi_cs_flash_LC_24_1_1 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.spi_cs_flash_LC_24_1_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \spi_slave_inst.spi_cs_flash_LC_24_1_1  (
            .in0(N__52296),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52414),
            .lcout(spi_cs_flash_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \spi_slave_inst.spi_sclk_flash_LC_24_1_5 .C_ON=1'b0;
    defparam \spi_slave_inst.spi_sclk_flash_LC_24_1_5 .SEQ_MODE=4'b0000;
    defparam \spi_slave_inst.spi_sclk_flash_LC_24_1_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \spi_slave_inst.spi_sclk_flash_LC_24_1_5  (
            .in0(N__52347),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52297),
            .lcout(spi_sclk_flash_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sCounterDAC_RNIBR1C_0_LC_24_10_3.C_ON=1'b0;
    defparam sCounterDAC_RNIBR1C_0_LC_24_10_3.SEQ_MODE=4'b0000;
    defparam sCounterDAC_RNIBR1C_0_LC_24_10_3.LUT_INIT=16'b0000100000000000;
    LogicCell40 sCounterDAC_RNIBR1C_0_LC_24_10_3 (
            .in0(N__53457),
            .in1(N__53436),
            .in2(N__53415),
            .in3(N__53364),
            .lcout(op_eq_scounterdac10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // MATTY_MAIN_VHDL
